-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Sep 14 2025 10:30:51

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DA : out std_logic_vector(2 downto 0);
    A : in std_logic_vector(20 downto 0);
    TBIn : out std_logic;
    RAMSPACEn : in std_logic;
    DBRn : in std_logic;
    RAMENn : out std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    PRnW : out std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    BLSn : out std_logic;
    TCIn : out std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__13161\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13006\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12684\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12549\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11967\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11714\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10629\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10177\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7257\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \N_112_0\ : std_logic;
signal \U712_REG_SM_REG_TACK_7_0\ : std_logic;
signal \N_19_0_cascade_\ : std_logic;
signal \U712_REG_SM_STATE_COUNT_3\ : std_logic;
signal \N_19_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_CHIP_RAM_m113_0\ : std_logic;
signal \U712_CHIP_RAM.N_87_0\ : std_logic;
signal \U712_CHIP_RAM.N_87_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_97_0_cascade_\ : std_logic;
signal \U712_REG_SM_STATE_COUNT_7\ : std_logic;
signal \U712_REG_SM_STATE_COUNT_0\ : std_logic;
signal \U712_CHIP_RAM.N_79_0\ : std_logic;
signal \U712_REG_SM_STATE_COUNT_5\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.N_103_0\ : std_logic;
signal \U712_REG_SM_STATE_COUNT_8\ : std_logic;
signal \U712_CHIP_RAM.N_103_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.m106_nsZ0Z_1\ : std_logic;
signal i62_mux : std_logic;
signal \U712_REG_SM_WRITE_CYCLE\ : std_logic;
signal \PRnW_c\ : std_logic;
signal \U712_CHIP_RAM.N_332\ : std_logic;
signal \INVU712_CYCLE_TERM.TACK_ENC_net\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_2\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \U712_CYCLE_TERM.TACK_RST_0_i\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_REG_SM_REG_CYCLE_START\ : std_logic;
signal \U712_REG_SM_START_RST\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_3\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U712_CHIP_RAM.m223_ns_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_4\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.m231_0\ : std_logic;
signal \U712_CHIP_RAM.N_236\ : std_logic;
signal \U712_REG_SM_STATE_COUNT_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_83_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_83_0\ : std_logic;
signal \U712_CHIP_RAM.N_94_0_cascade_\ : std_logic;
signal \U712_REG_SM_STATE_COUNT_1\ : std_logic;
signal \U712_REG_SM_STATE_COUNT_2\ : std_logic;
signal \DBR_SYNC_i_1\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ1Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_7_0\ : std_logic;
signal \N_86_0\ : std_logic;
signal \U712_REG_SM_C3_SYNC_1\ : std_logic;
signal \BLSn_c\ : std_logic;
signal \U712_REG_SM.N_86_0_0\ : std_logic;
signal \U712_CYCLE_TERM.N_36_0_cascade_\ : std_logic;
signal \TACK_OUT\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STARTZ0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \INVU712_CYCLE_TERM.TACK_OUTC_net\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_146_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_154_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.m38_1\ : std_logic;
signal \U712_CHIP_RAM.N_34_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_359\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_28_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_47_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_215\ : std_logic;
signal \bfn_10_14_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.N_56_0_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.N_330\ : std_logic;
signal \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\ : std_logic;
signal \U712_REG_SM_UDSn_6_0\ : std_logic;
signal \UDSn_c\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \A_c_9\ : std_logic;
signal \U712_CHIP_RAM.m186_0_cascade_\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U712_CHIP_RAM.m192_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.m192_1\ : std_logic;
signal \U712_CHIP_RAM.d_N_6_5\ : std_logic;
signal \U712_CHIP_RAM.d_N_6_1\ : std_logic;
signal \U712_CHIP_RAM.N_353_mux\ : std_logic;
signal \U712_CHIP_RAM.N_168_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.m64_ns_1\ : std_logic;
signal \U712_CHIP_RAM.i67_mux_cascade_\ : std_logic;
signal \U712_CHIP_RAM.m66_ns_1\ : std_logic;
signal \U712_CHIP_RAM.N_146_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_151_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_2\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lt7\ : std_logic;
signal \U712_CHIP_RAM.N_28_0\ : std_logic;
signal \U712_CHIP_RAM.N_219\ : std_logic;
signal \U712_CHIP_RAM.m41_1\ : std_logic;
signal \U712_CHIP_RAM.N_31_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.m217_ns_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_218\ : std_logic;
signal \U712_CHIP_RAM.m212_ns_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_30_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_213\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.N_333_mux_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_51_0\ : std_logic;
signal \U712_CHIP_RAM.N_51_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_54_0\ : std_logic;
signal \U712_CHIP_RAM.m53_ns_1\ : std_logic;
signal \U712_CHIP_RAM.N_333_mux\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \U712_CHIP_RAM.m189_1\ : std_logic;
signal \U712_CHIP_RAM.m188_1\ : std_logic;
signal \U712_CHIP_RAM.d_N_6_2\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U712_CHIP_RAM.m188_0\ : std_logic;
signal \U712_CHIP_RAM.d_N_6\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U712_CHIP_RAM.m189_0\ : std_logic;
signal \A_c_14\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \U712_CHIP_RAM.m186_1\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.N_198_cascade_\ : std_logic;
signal \CLK40_PLL\ : std_logic;
signal \CLK40_PLL_iso_i\ : std_logic;
signal \U712_CHIP_RAM.m187_1\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.N_3_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.m187_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_163_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_67_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.N_48_0\ : std_logic;
signal \U712_CHIP_RAM.N_363\ : std_logic;
signal \U712_CHIP_RAM.N_158_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_58_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.d_N_6_0\ : std_logic;
signal \U712_CHIP_RAM.N_43_0\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\ : std_logic;
signal \A_c_6\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_START_RNIJD6OZ0Z3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_204_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_364\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.N_26_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_30_0\ : std_logic;
signal \U712_CHIP_RAM.N_62_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_RNI9THUZ0Z5\ : std_logic;
signal \U712_CHIP_RAM.CLK_EN_RNOZ0Z_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CLK_EN_RNOZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_174_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER43\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.N_62_0\ : std_logic;
signal \U712_CHIP_RAM.N_52_0\ : std_logic;
signal \U712_CHIP_RAM.N_208_cascade_\ : std_logic;
signal \N_99_0\ : std_logic;
signal \LDSn_c\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \RASn_c\ : std_logic;
signal \U712_CHIP_RAM.d_N_7\ : std_logic;
signal \U712_CHIP_RAM.m185_0\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U712_CHIP_RAM.m191_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.d_N_6_4\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.m184_m2_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.m184_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.m184_1\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U712_CHIP_RAM.N_3_0\ : std_logic;
signal \U712_CHIP_RAM.m186_m2_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.m190_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.m190_1\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.d_N_6_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.d_N_7_0\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.N_204\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_31_0\ : std_logic;
signal \U712_CHIP_RAM.DBENn_8_0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0\ : std_logic;
signal \LATCH_CLK_c\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.N_99_0_0\ : std_logic;
signal \U712_REG_SM_C1_SYNC_1\ : std_logic;
signal \U712_REG_SM_LDSn_6_0\ : std_logic;
signal \U712_CHIP_RAM.m185_1\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \A_c_19\ : std_logic;
signal \U712_CHIP_RAM.m194_0\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.m191_1\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.N_198_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \CUMBEn_c\ : std_logic;
signal \LMBEn_c\ : std_logic;
signal \CLMBEn_c\ : std_logic;
signal \CUUBEn_c\ : std_logic;
signal \U712_CHIP_RAM.N_346\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \U712_CHIP_RAM.N_346_cascade_\ : std_logic;
signal \CLLBEn_c\ : std_logic;
signal \LLBEn_c\ : std_logic;
signal \A_c_0\ : std_logic;
signal \UUBEn_c\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \A_c_1\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \U712_CHIP_RAM.N_325_mux\ : std_logic;
signal \UMBEn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \WEn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.N_345\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \DMA_LATCH_EN_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_0\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLEm\ : std_logic;
signal \N_338_mux\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_WRITE_CYCLEZ0\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \N_328_mux\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \DA_wire\ : std_logic_vector(2 downto 0);
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \PRnW_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \BLSn_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    TBIn <= \TBIn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    ASn <= \ASn_wire\;
    DA <= \DA_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    TCIn <= \TCIn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    PRnW <= \PRnW_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    \C3_wire\ <= C3;
    BLSn <= \BLSn_wire\;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL\,
            REFERENCECLK => \N__4511\,
            RESETB => \N__8729\,
            BYPASS => \GNDG0\,
            PLLOUTCOREA => OPEN,
            SDI => \GNDG0\,
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => \GNDG0\,
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => \GNDG0\
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13161\,
            DIN => \N__13160\,
            DOUT => \N__13159\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13161\,
            PADOUT => \N__13160\,
            PADIN => \N__13159\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10274\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13152\,
            DIN => \N__13151\,
            DOUT => \N__13150\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13152\,
            PADOUT => \N__13151\,
            PADIN => \N__13150\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13143\,
            DIN => \N__13142\,
            DOUT => \N__13141\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13143\,
            PADOUT => \N__13142\,
            PADIN => \N__13141\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12026\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13134\,
            DIN => \N__13133\,
            DOUT => \N__13132\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13134\,
            PADOUT => \N__13133\,
            PADIN => \N__13132\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10661\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13125\,
            DIN => \N__13124\,
            DOUT => \N__13123\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13125\,
            PADOUT => \N__13124\,
            PADIN => \N__13123\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13116\,
            DIN => \N__13115\,
            DOUT => \N__13114\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13116\,
            PADOUT => \N__13115\,
            PADIN => \N__13114\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13107\,
            DIN => \N__13106\,
            DOUT => \N__13105\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13107\,
            PADOUT => \N__13106\,
            PADIN => \N__13105\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13098\,
            DIN => \N__13097\,
            DOUT => \N__13096\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13098\,
            PADOUT => \N__13097\,
            PADIN => \N__13096\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13089\,
            DIN => \N__13088\,
            DOUT => \N__13087\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13089\,
            PADOUT => \N__13088\,
            PADIN => \N__13087\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13080\,
            DIN => \N__13079\,
            DOUT => \N__13078\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13080\,
            PADOUT => \N__13079\,
            PADIN => \N__13078\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13071\,
            DIN => \N__13070\,
            DOUT => \N__13069\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13071\,
            PADOUT => \N__13070\,
            PADIN => \N__13069\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13062\,
            DIN => \N__13061\,
            DOUT => \N__13060\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13062\,
            PADOUT => \N__13061\,
            PADIN => \N__13060\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9692\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13053\,
            DIN => \N__13052\,
            DOUT => \N__13051\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13053\,
            PADOUT => \N__13052\,
            PADIN => \N__13051\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10121\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13044\,
            DIN => \N__13043\,
            DOUT => \N__13042\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13044\,
            PADOUT => \N__13043\,
            PADIN => \N__13042\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13035\,
            DIN => \N__13034\,
            DOUT => \N__13033\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13035\,
            PADOUT => \N__13034\,
            PADIN => \N__13033\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5161\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13026\,
            DIN => \N__13025\,
            DOUT => \N__13024\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13026\,
            PADOUT => \N__13025\,
            PADIN => \N__13024\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13017\,
            DIN => \N__13016\,
            DOUT => \N__13015\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13017\,
            PADOUT => \N__13016\,
            PADIN => \N__13015\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13008\,
            DIN => \N__13007\,
            DOUT => \N__13006\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13008\,
            PADOUT => \N__13007\,
            PADIN => \N__13006\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4676\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12999\,
            DIN => \N__12998\,
            DOUT => \N__12997\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12999\,
            PADOUT => \N__12998\,
            PADIN => \N__12997\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12990\,
            DIN => \N__12989\,
            DOUT => \N__12988\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12990\,
            PADOUT => \N__12989\,
            PADIN => \N__12988\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12981\,
            DIN => \N__12980\,
            DOUT => \N__12979\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12981\,
            PADOUT => \N__12980\,
            PADIN => \N__12979\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6905\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12972\,
            DIN => \N__12971\,
            DOUT => \N__12970\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12972\,
            PADOUT => \N__12971\,
            PADIN => \N__12970\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12963\,
            DIN => \N__12962\,
            DOUT => \N__12961\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12963\,
            PADOUT => \N__12962\,
            PADIN => \N__12961\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11960\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12954\,
            DIN => \N__12953\,
            DOUT => \N__12952\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12954\,
            PADOUT => \N__12953\,
            PADIN => \N__12952\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12945\,
            DIN => \N__12944\,
            DOUT => \N__12943\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12945\,
            PADOUT => \N__12944\,
            PADIN => \N__12943\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10193\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12936\,
            DIN => \N__12935\,
            DOUT => \N__12934\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12936\,
            PADOUT => \N__12935\,
            PADIN => \N__12934\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4878\,
            DIN0 => OPEN,
            DOUT0 => \N__5562\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12927\,
            DIN => \N__12926\,
            DOUT => \N__12925\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12927\,
            PADOUT => \N__12926\,
            PADIN => \N__12925\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12918\,
            DIN => \N__12917\,
            DOUT => \N__12916\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12918\,
            PADOUT => \N__12917\,
            PADIN => \N__12916\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12909\,
            DIN => \N__12908\,
            DOUT => \N__12907\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12909\,
            PADOUT => \N__12908\,
            PADIN => \N__12907\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12900\,
            DIN => \N__12899\,
            DOUT => \N__12898\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12900\,
            PADOUT => \N__12899\,
            PADIN => \N__12898\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12891\,
            DIN => \N__12890\,
            DOUT => \N__12889\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12891\,
            PADOUT => \N__12890\,
            PADIN => \N__12889\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12882\,
            DIN => \N__12881\,
            DOUT => \N__12880\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12882\,
            PADOUT => \N__12881\,
            PADIN => \N__12880\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12269\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12873\,
            DIN => \N__12872\,
            DOUT => \N__12871\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12873\,
            PADOUT => \N__12872\,
            PADIN => \N__12871\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12864\,
            DIN => \N__12863\,
            DOUT => \N__12862\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12864\,
            PADOUT => \N__12863\,
            PADIN => \N__12862\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12855\,
            DIN => \N__12854\,
            DOUT => \N__12853\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12855\,
            PADOUT => \N__12854\,
            PADIN => \N__12853\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12846\,
            DIN => \N__12845\,
            DOUT => \N__12844\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12846\,
            PADOUT => \N__12845\,
            PADIN => \N__12844\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12837\,
            DIN => \N__12836\,
            DOUT => \N__12835\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12837\,
            PADOUT => \N__12836\,
            PADIN => \N__12835\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12828\,
            DIN => \N__12827\,
            DOUT => \N__12826\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12828\,
            PADOUT => \N__12827\,
            PADIN => \N__12826\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7910\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12819\,
            DIN => \N__12818\,
            DOUT => \N__12817\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12819\,
            PADOUT => \N__12818\,
            PADIN => \N__12817\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12810\,
            DIN => \N__12809\,
            DOUT => \N__12808\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12810\,
            PADOUT => \N__12809\,
            PADIN => \N__12808\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12801\,
            DIN => \N__12800\,
            DOUT => \N__12799\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12801\,
            PADOUT => \N__12800\,
            PADIN => \N__12799\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9485\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12792\,
            DIN => \N__12791\,
            DOUT => \N__12790\,
            PACKAGEPIN => \DA_wire\(0)
        );

    \DA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12792\,
            PADOUT => \N__12791\,
            PADIN => \N__12790\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6020\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12783\,
            DIN => \N__12782\,
            DOUT => \N__12781\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12783\,
            PADOUT => \N__12782\,
            PADIN => \N__12781\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12774\,
            DIN => \N__12773\,
            DOUT => \N__12772\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12774\,
            PADOUT => \N__12773\,
            PADIN => \N__12772\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6722\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12765\,
            DIN => \N__12764\,
            DOUT => \N__12763\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12765\,
            PADOUT => \N__12764\,
            PADIN => \N__12763\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6770\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12756\,
            DIN => \N__12755\,
            DOUT => \N__12754\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12756\,
            PADOUT => \N__12755\,
            PADIN => \N__12754\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5614\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12747\,
            DIN => \N__12746\,
            DOUT => \N__12745\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12747\,
            PADOUT => \N__12746\,
            PADIN => \N__12745\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12738\,
            DIN => \N__12737\,
            DOUT => \N__12736\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12738\,
            PADOUT => \N__12737\,
            PADIN => \N__12736\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9524\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12729\,
            DIN => \N__12728\,
            DOUT => \N__12727\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12729\,
            PADOUT => \N__12728\,
            PADIN => \N__12727\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4883\,
            DIN0 => OPEN,
            DOUT0 => \N__5563\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12720\,
            DIN => \N__12719\,
            DOUT => \N__12718\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12720\,
            PADOUT => \N__12719\,
            PADIN => \N__12718\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9821\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12711\,
            DIN => \N__12710\,
            DOUT => \N__12709\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12711\,
            PADOUT => \N__12710\,
            PADIN => \N__12709\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7235\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12702\,
            DIN => \N__12701\,
            DOUT => \N__12700\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12702\,
            PADOUT => \N__12701\,
            PADIN => \N__12700\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9578\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12693\,
            DIN => \N__12692\,
            DOUT => \N__12691\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12693\,
            PADOUT => \N__12692\,
            PADIN => \N__12691\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12684\,
            DIN => \N__12683\,
            DOUT => \N__12682\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12684\,
            PADOUT => \N__12683\,
            PADIN => \N__12682\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12675\,
            DIN => \N__12674\,
            DOUT => \N__12673\,
            PACKAGEPIN => \DA_wire\(2)
        );

    \DA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12675\,
            PADOUT => \N__12674\,
            PADIN => \N__12673\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7205\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12666\,
            DIN => \N__12665\,
            DOUT => \N__12664\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12666\,
            PADOUT => \N__12665\,
            PADIN => \N__12664\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12657\,
            DIN => \N__12656\,
            DOUT => \N__12655\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12657\,
            PADOUT => \N__12656\,
            PADIN => \N__12655\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12648\,
            DIN => \N__12647\,
            DOUT => \N__12646\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12648\,
            PADOUT => \N__12647\,
            PADIN => \N__12646\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6884\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12639\,
            DIN => \N__12638\,
            DOUT => \N__12637\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12639\,
            PADOUT => \N__12638\,
            PADIN => \N__12637\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9554\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12630\,
            DIN => \N__12629\,
            DOUT => \N__12628\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12630\,
            PADOUT => \N__12629\,
            PADIN => \N__12628\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12621\,
            DIN => \N__12620\,
            DOUT => \N__12619\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12621\,
            PADOUT => \N__12620\,
            PADIN => \N__12619\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9503\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12612\,
            DIN => \N__12611\,
            DOUT => \N__12610\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12612\,
            PADOUT => \N__12611\,
            PADIN => \N__12610\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4882\,
            DIN0 => OPEN,
            DOUT0 => \N__5564\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12603\,
            DIN => \N__12602\,
            DOUT => \N__12601\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12603\,
            PADOUT => \N__12602\,
            PADIN => \N__12601\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6929\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12594\,
            DIN => \N__12593\,
            DOUT => \N__12592\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12594\,
            PADOUT => \N__12593\,
            PADIN => \N__12592\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12585\,
            DIN => \N__12584\,
            DOUT => \N__12583\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12585\,
            PADOUT => \N__12584\,
            PADIN => \N__12583\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12576\,
            DIN => \N__12575\,
            DOUT => \N__12574\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12576\,
            PADOUT => \N__12575\,
            PADIN => \N__12574\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6041\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12567\,
            DIN => \N__12566\,
            DOUT => \N__12565\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12567\,
            PADOUT => \N__12566\,
            PADIN => \N__12565\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12558\,
            DIN => \N__12557\,
            DOUT => \N__12556\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12558\,
            PADOUT => \N__12557\,
            PADIN => \N__12556\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12549\,
            DIN => \N__12548\,
            DOUT => \N__12547\,
            PACKAGEPIN => \DA_wire\(1)
        );

    \DA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12549\,
            PADOUT => \N__12548\,
            PADIN => \N__12547\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8471\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12540\,
            DIN => \N__12539\,
            DOUT => \N__12538\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12540\,
            PADOUT => \N__12539\,
            PADIN => \N__12538\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12531\,
            DIN => \N__12530\,
            DOUT => \N__12529\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12531\,
            PADOUT => \N__12530\,
            PADIN => \N__12529\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12522\,
            DIN => \N__12521\,
            DOUT => \N__12520\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12522\,
            PADOUT => \N__12521\,
            PADIN => \N__12520\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9329\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12513\,
            DIN => \N__12512\,
            DOUT => \N__12511\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12513\,
            PADOUT => \N__12512\,
            PADIN => \N__12511\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6098\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12504\,
            DIN => \N__12503\,
            DOUT => \N__12502\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12504\,
            PADOUT => \N__12503\,
            PADIN => \N__12502\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9923\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12495\,
            DIN => \N__12494\,
            DOUT => \N__12493\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12495\,
            PADOUT => \N__12494\,
            PADIN => \N__12493\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7613\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12486\,
            DIN => \N__12485\,
            DOUT => \N__12484\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12486\,
            PADOUT => \N__12485\,
            PADIN => \N__12484\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12477\,
            DIN => \N__12476\,
            DOUT => \N__12475\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12477\,
            PADOUT => \N__12476\,
            PADIN => \N__12475\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12468\,
            DIN => \N__12467\,
            DOUT => \N__12466\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12468\,
            PADOUT => \N__12467\,
            PADIN => \N__12466\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8243\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12459\,
            DIN => \N__12458\,
            DOUT => \N__12457\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12459\,
            PADOUT => \N__12458\,
            PADIN => \N__12457\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12450\,
            DIN => \N__12449\,
            DOUT => \N__12448\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12450\,
            PADOUT => \N__12449\,
            PADIN => \N__12448\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12441\,
            DIN => \N__12440\,
            DOUT => \N__12439\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12441\,
            PADOUT => \N__12440\,
            PADIN => \N__12439\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8507\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12432\,
            DIN => \N__12431\,
            DOUT => \N__12430\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12432\,
            PADOUT => \N__12431\,
            PADIN => \N__12430\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8177\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12423\,
            DIN => \N__12422\,
            DOUT => \N__12421\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12423\,
            PADOUT => \N__12422\,
            PADIN => \N__12421\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6831\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PRnW_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12414\,
            DIN => \N__12413\,
            DOUT => \N__12412\,
            PACKAGEPIN => \PRnW_wire\
        );

    \PRnW_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12414\,
            PADOUT => \N__12413\,
            PADIN => \N__12412\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4931\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12405\,
            DIN => \N__12404\,
            DOUT => \N__12403\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12405\,
            PADOUT => \N__12404\,
            PADIN => \N__12403\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12396\,
            DIN => \N__12395\,
            DOUT => \N__12394\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12396\,
            PADOUT => \N__12395\,
            PADIN => \N__12394\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6833\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12387\,
            DIN => \N__12386\,
            DOUT => \N__12385\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12387\,
            PADOUT => \N__12386\,
            PADIN => \N__12385\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4526\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12378\,
            DIN => \N__12377\,
            DOUT => \N__12376\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12378\,
            PADOUT => \N__12377\,
            PADIN => \N__12376\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6746\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12369\,
            DIN => \N__12368\,
            DOUT => \N__12367\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12369\,
            PADOUT => \N__12368\,
            PADIN => \N__12367\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12360\,
            DIN => \N__12359\,
            DOUT => \N__12358\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12360\,
            PADOUT => \N__12359\,
            PADIN => \N__12358\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12351\,
            DIN => \N__12350\,
            DOUT => \N__12349\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12351\,
            PADOUT => \N__12350\,
            PADIN => \N__12349\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BLSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12342\,
            DIN => \N__12341\,
            DOUT => \N__12340\,
            PACKAGEPIN => \BLSn_wire\
        );

    \BLSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12342\,
            PADOUT => \N__12341\,
            PADIN => \N__12340\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5618\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12333\,
            DIN => \N__12332\,
            DOUT => \N__12331\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12333\,
            PADOUT => \N__12332\,
            PADIN => \N__12331\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12324\,
            DIN => \N__12323\,
            DOUT => \N__12322\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12324\,
            PADOUT => \N__12323\,
            PADIN => \N__12322\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6832\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12315\,
            DIN => \N__12314\,
            DOUT => \N__12313\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12315\,
            PADOUT => \N__12314\,
            PADIN => \N__12313\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10871\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12306\,
            DIN => \N__12305\,
            DOUT => \N__12304\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12306\,
            PADOUT => \N__12305\,
            PADIN => \N__12304\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10214\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12297\,
            DIN => \N__12296\,
            DOUT => \N__12295\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12297\,
            PADOUT => \N__12296\,
            PADIN => \N__12295\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9263\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12288\,
            DIN => \N__12287\,
            DOUT => \N__12286\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12288\,
            PADOUT => \N__12287\,
            PADIN => \N__12286\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2982\ : IoInMux
    port map (
            O => \N__12269\,
            I => \N__12266\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__12266\,
            I => \N__12263\
        );

    \I__2980\ : Span4Mux_s3_v
    port map (
            O => \N__12263\,
            I => \N__12260\
        );

    \I__2979\ : Span4Mux_v
    port map (
            O => \N__12260\,
            I => \N__12257\
        );

    \I__2978\ : Sp12to4
    port map (
            O => \N__12257\,
            I => \N__12254\
        );

    \I__2977\ : Span12Mux_h
    port map (
            O => \N__12254\,
            I => \N__12251\
        );

    \I__2976\ : Odrv12
    port map (
            O => \N__12251\,
            I => \DMA_LATCH_EN_c\
        );

    \I__2975\ : CascadeMux
    port map (
            O => \N__12248\,
            I => \N__12244\
        );

    \I__2974\ : InMux
    port map (
            O => \N__12247\,
            I => \N__12237\
        );

    \I__2973\ : InMux
    port map (
            O => \N__12244\,
            I => \N__12234\
        );

    \I__2972\ : CascadeMux
    port map (
            O => \N__12243\,
            I => \N__12231\
        );

    \I__2971\ : CascadeMux
    port map (
            O => \N__12242\,
            I => \N__12221\
        );

    \I__2970\ : CascadeMux
    port map (
            O => \N__12241\,
            I => \N__12218\
        );

    \I__2969\ : CascadeMux
    port map (
            O => \N__12240\,
            I => \N__12215\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__12237\,
            I => \N__12209\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__12234\,
            I => \N__12209\
        );

    \I__2966\ : InMux
    port map (
            O => \N__12231\,
            I => \N__12206\
        );

    \I__2965\ : InMux
    port map (
            O => \N__12230\,
            I => \N__12203\
        );

    \I__2964\ : CascadeMux
    port map (
            O => \N__12229\,
            I => \N__12200\
        );

    \I__2963\ : CascadeMux
    port map (
            O => \N__12228\,
            I => \N__12196\
        );

    \I__2962\ : CascadeMux
    port map (
            O => \N__12227\,
            I => \N__12193\
        );

    \I__2961\ : CascadeMux
    port map (
            O => \N__12226\,
            I => \N__12190\
        );

    \I__2960\ : CascadeMux
    port map (
            O => \N__12225\,
            I => \N__12187\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__12224\,
            I => \N__12178\
        );

    \I__2958\ : InMux
    port map (
            O => \N__12221\,
            I => \N__12171\
        );

    \I__2957\ : InMux
    port map (
            O => \N__12218\,
            I => \N__12171\
        );

    \I__2956\ : InMux
    port map (
            O => \N__12215\,
            I => \N__12171\
        );

    \I__2955\ : InMux
    port map (
            O => \N__12214\,
            I => \N__12168\
        );

    \I__2954\ : Span4Mux_h
    port map (
            O => \N__12209\,
            I => \N__12165\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__12206\,
            I => \N__12160\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__12203\,
            I => \N__12157\
        );

    \I__2951\ : InMux
    port map (
            O => \N__12200\,
            I => \N__12154\
        );

    \I__2950\ : InMux
    port map (
            O => \N__12199\,
            I => \N__12141\
        );

    \I__2949\ : InMux
    port map (
            O => \N__12196\,
            I => \N__12141\
        );

    \I__2948\ : InMux
    port map (
            O => \N__12193\,
            I => \N__12141\
        );

    \I__2947\ : InMux
    port map (
            O => \N__12190\,
            I => \N__12134\
        );

    \I__2946\ : InMux
    port map (
            O => \N__12187\,
            I => \N__12134\
        );

    \I__2945\ : InMux
    port map (
            O => \N__12186\,
            I => \N__12134\
        );

    \I__2944\ : InMux
    port map (
            O => \N__12185\,
            I => \N__12127\
        );

    \I__2943\ : InMux
    port map (
            O => \N__12184\,
            I => \N__12127\
        );

    \I__2942\ : InMux
    port map (
            O => \N__12183\,
            I => \N__12127\
        );

    \I__2941\ : CascadeMux
    port map (
            O => \N__12182\,
            I => \N__12124\
        );

    \I__2940\ : CascadeMux
    port map (
            O => \N__12181\,
            I => \N__12115\
        );

    \I__2939\ : InMux
    port map (
            O => \N__12178\,
            I => \N__12112\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__12171\,
            I => \N__12107\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__12168\,
            I => \N__12107\
        );

    \I__2936\ : Span4Mux_v
    port map (
            O => \N__12165\,
            I => \N__12104\
        );

    \I__2935\ : InMux
    port map (
            O => \N__12164\,
            I => \N__12099\
        );

    \I__2934\ : InMux
    port map (
            O => \N__12163\,
            I => \N__12099\
        );

    \I__2933\ : Span4Mux_h
    port map (
            O => \N__12160\,
            I => \N__12092\
        );

    \I__2932\ : Span4Mux_v
    port map (
            O => \N__12157\,
            I => \N__12092\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__12154\,
            I => \N__12092\
        );

    \I__2930\ : InMux
    port map (
            O => \N__12153\,
            I => \N__12085\
        );

    \I__2929\ : InMux
    port map (
            O => \N__12152\,
            I => \N__12085\
        );

    \I__2928\ : InMux
    port map (
            O => \N__12151\,
            I => \N__12085\
        );

    \I__2927\ : InMux
    port map (
            O => \N__12150\,
            I => \N__12080\
        );

    \I__2926\ : InMux
    port map (
            O => \N__12149\,
            I => \N__12080\
        );

    \I__2925\ : InMux
    port map (
            O => \N__12148\,
            I => \N__12077\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__12141\,
            I => \N__12070\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__12134\,
            I => \N__12070\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__12127\,
            I => \N__12070\
        );

    \I__2921\ : InMux
    port map (
            O => \N__12124\,
            I => \N__12063\
        );

    \I__2920\ : InMux
    port map (
            O => \N__12123\,
            I => \N__12063\
        );

    \I__2919\ : InMux
    port map (
            O => \N__12122\,
            I => \N__12063\
        );

    \I__2918\ : InMux
    port map (
            O => \N__12121\,
            I => \N__12056\
        );

    \I__2917\ : InMux
    port map (
            O => \N__12120\,
            I => \N__12056\
        );

    \I__2916\ : InMux
    port map (
            O => \N__12119\,
            I => \N__12056\
        );

    \I__2915\ : InMux
    port map (
            O => \N__12118\,
            I => \N__12051\
        );

    \I__2914\ : InMux
    port map (
            O => \N__12115\,
            I => \N__12051\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__12112\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2912\ : Odrv4
    port map (
            O => \N__12107\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2911\ : Odrv4
    port map (
            O => \N__12104\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__12099\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2909\ : Odrv4
    port map (
            O => \N__12092\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__12085\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__12080\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__12077\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2905\ : Odrv12
    port map (
            O => \N__12070\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__12063\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__12056\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__12051\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2901\ : IoInMux
    port map (
            O => \N__12026\,
            I => \N__12023\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__12023\,
            I => \N__12020\
        );

    \I__2899\ : Span12Mux_s9_v
    port map (
            O => \N__12020\,
            I => \N__12017\
        );

    \I__2898\ : Odrv12
    port map (
            O => \N__12017\,
            I => \CASn_c\
        );

    \I__2897\ : InMux
    port map (
            O => \N__12014\,
            I => \N__12010\
        );

    \I__2896\ : InMux
    port map (
            O => \N__12013\,
            I => \N__12007\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__12010\,
            I => \N__12003\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__12007\,
            I => \N__12000\
        );

    \I__2893\ : CascadeMux
    port map (
            O => \N__12006\,
            I => \N__11997\
        );

    \I__2892\ : Span4Mux_h
    port map (
            O => \N__12003\,
            I => \N__11991\
        );

    \I__2891\ : Span4Mux_h
    port map (
            O => \N__12000\,
            I => \N__11991\
        );

    \I__2890\ : InMux
    port map (
            O => \N__11997\,
            I => \N__11988\
        );

    \I__2889\ : InMux
    port map (
            O => \N__11996\,
            I => \N__11985\
        );

    \I__2888\ : Span4Mux_v
    port map (
            O => \N__11991\,
            I => \N__11979\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__11988\,
            I => \N__11979\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__11985\,
            I => \N__11976\
        );

    \I__2885\ : InMux
    port map (
            O => \N__11984\,
            I => \N__11973\
        );

    \I__2884\ : Span4Mux_h
    port map (
            O => \N__11979\,
            I => \N__11970\
        );

    \I__2883\ : Span4Mux_h
    port map (
            O => \N__11976\,
            I => \N__11967\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__11973\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2881\ : Odrv4
    port map (
            O => \N__11970\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2880\ : Odrv4
    port map (
            O => \N__11967\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2879\ : IoInMux
    port map (
            O => \N__11960\,
            I => \N__11957\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__11957\,
            I => \N__11954\
        );

    \I__2877\ : Span4Mux_s1_v
    port map (
            O => \N__11954\,
            I => \N__11951\
        );

    \I__2876\ : Span4Mux_v
    port map (
            O => \N__11951\,
            I => \N__11948\
        );

    \I__2875\ : Span4Mux_v
    port map (
            O => \N__11948\,
            I => \N__11945\
        );

    \I__2874\ : Odrv4
    port map (
            O => \N__11945\,
            I => \CRCSn_c\
        );

    \I__2873\ : InMux
    port map (
            O => \N__11942\,
            I => \N__11939\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__11939\,
            I => \N__11933\
        );

    \I__2871\ : InMux
    port map (
            O => \N__11938\,
            I => \N__11930\
        );

    \I__2870\ : InMux
    port map (
            O => \N__11937\,
            I => \N__11927\
        );

    \I__2869\ : InMux
    port map (
            O => \N__11936\,
            I => \N__11924\
        );

    \I__2868\ : Span4Mux_v
    port map (
            O => \N__11933\,
            I => \N__11921\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__11930\,
            I => \N__11918\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__11927\,
            I => \N__11913\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__11924\,
            I => \N__11913\
        );

    \I__2864\ : Span4Mux_h
    port map (
            O => \N__11921\,
            I => \N__11908\
        );

    \I__2863\ : Span4Mux_v
    port map (
            O => \N__11918\,
            I => \N__11908\
        );

    \I__2862\ : Span12Mux_v
    port map (
            O => \N__11913\,
            I => \N__11905\
        );

    \I__2861\ : Sp12to4
    port map (
            O => \N__11908\,
            I => \N__11902\
        );

    \I__2860\ : Span12Mux_h
    port map (
            O => \N__11905\,
            I => \N__11899\
        );

    \I__2859\ : Odrv12
    port map (
            O => \N__11902\,
            I => \DRA_c_8\
        );

    \I__2858\ : Odrv12
    port map (
            O => \N__11899\,
            I => \DRA_c_8\
        );

    \I__2857\ : InMux
    port map (
            O => \N__11894\,
            I => \N__11890\
        );

    \I__2856\ : InMux
    port map (
            O => \N__11893\,
            I => \N__11887\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__11890\,
            I => \N__11880\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__11887\,
            I => \N__11880\
        );

    \I__2853\ : InMux
    port map (
            O => \N__11886\,
            I => \N__11877\
        );

    \I__2852\ : InMux
    port map (
            O => \N__11885\,
            I => \N__11874\
        );

    \I__2851\ : Span4Mux_h
    port map (
            O => \N__11880\,
            I => \N__11867\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__11877\,
            I => \N__11867\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__11874\,
            I => \N__11867\
        );

    \I__2848\ : Span4Mux_v
    port map (
            O => \N__11867\,
            I => \N__11864\
        );

    \I__2847\ : Sp12to4
    port map (
            O => \N__11864\,
            I => \N__11861\
        );

    \I__2846\ : Span12Mux_h
    port map (
            O => \N__11861\,
            I => \N__11858\
        );

    \I__2845\ : Odrv12
    port map (
            O => \N__11858\,
            I => \DRA_c_7\
        );

    \I__2844\ : InMux
    port map (
            O => \N__11855\,
            I => \N__11852\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__11852\,
            I => \N__11849\
        );

    \I__2842\ : Odrv4
    port map (
            O => \N__11849\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2841\ : InMux
    port map (
            O => \N__11846\,
            I => \N__11842\
        );

    \I__2840\ : InMux
    port map (
            O => \N__11845\,
            I => \N__11838\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__11842\,
            I => \N__11835\
        );

    \I__2838\ : InMux
    port map (
            O => \N__11841\,
            I => \N__11832\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__11838\,
            I => \N__11829\
        );

    \I__2836\ : Span4Mux_v
    port map (
            O => \N__11835\,
            I => \N__11825\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__11832\,
            I => \N__11822\
        );

    \I__2834\ : Span4Mux_h
    port map (
            O => \N__11829\,
            I => \N__11819\
        );

    \I__2833\ : InMux
    port map (
            O => \N__11828\,
            I => \N__11816\
        );

    \I__2832\ : Span4Mux_h
    port map (
            O => \N__11825\,
            I => \N__11811\
        );

    \I__2831\ : Span4Mux_v
    port map (
            O => \N__11822\,
            I => \N__11811\
        );

    \I__2830\ : Sp12to4
    port map (
            O => \N__11819\,
            I => \N__11806\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__11816\,
            I => \N__11806\
        );

    \I__2828\ : Span4Mux_v
    port map (
            O => \N__11811\,
            I => \N__11803\
        );

    \I__2827\ : Span12Mux_v
    port map (
            O => \N__11806\,
            I => \N__11798\
        );

    \I__2826\ : Sp12to4
    port map (
            O => \N__11803\,
            I => \N__11798\
        );

    \I__2825\ : Span12Mux_h
    port map (
            O => \N__11798\,
            I => \N__11795\
        );

    \I__2824\ : Span12Mux_v
    port map (
            O => \N__11795\,
            I => \N__11792\
        );

    \I__2823\ : Odrv12
    port map (
            O => \N__11792\,
            I => \DRA_c_9\
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__11789\,
            I => \N__11786\
        );

    \I__2821\ : InMux
    port map (
            O => \N__11786\,
            I => \N__11783\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__11783\,
            I => \N__11772\
        );

    \I__2819\ : CascadeMux
    port map (
            O => \N__11782\,
            I => \N__11769\
        );

    \I__2818\ : InMux
    port map (
            O => \N__11781\,
            I => \N__11766\
        );

    \I__2817\ : InMux
    port map (
            O => \N__11780\,
            I => \N__11761\
        );

    \I__2816\ : InMux
    port map (
            O => \N__11779\,
            I => \N__11761\
        );

    \I__2815\ : InMux
    port map (
            O => \N__11778\,
            I => \N__11756\
        );

    \I__2814\ : InMux
    port map (
            O => \N__11777\,
            I => \N__11756\
        );

    \I__2813\ : InMux
    port map (
            O => \N__11776\,
            I => \N__11753\
        );

    \I__2812\ : InMux
    port map (
            O => \N__11775\,
            I => \N__11743\
        );

    \I__2811\ : Span4Mux_v
    port map (
            O => \N__11772\,
            I => \N__11740\
        );

    \I__2810\ : InMux
    port map (
            O => \N__11769\,
            I => \N__11737\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__11766\,
            I => \N__11728\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__11761\,
            I => \N__11728\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__11756\,
            I => \N__11728\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__11753\,
            I => \N__11728\
        );

    \I__2805\ : InMux
    port map (
            O => \N__11752\,
            I => \N__11723\
        );

    \I__2804\ : InMux
    port map (
            O => \N__11751\,
            I => \N__11723\
        );

    \I__2803\ : InMux
    port map (
            O => \N__11750\,
            I => \N__11720\
        );

    \I__2802\ : InMux
    port map (
            O => \N__11749\,
            I => \N__11717\
        );

    \I__2801\ : InMux
    port map (
            O => \N__11748\,
            I => \N__11714\
        );

    \I__2800\ : InMux
    port map (
            O => \N__11747\,
            I => \N__11711\
        );

    \I__2799\ : InMux
    port map (
            O => \N__11746\,
            I => \N__11707\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__11743\,
            I => \N__11702\
        );

    \I__2797\ : Span4Mux_v
    port map (
            O => \N__11740\,
            I => \N__11695\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__11737\,
            I => \N__11695\
        );

    \I__2795\ : Span4Mux_v
    port map (
            O => \N__11728\,
            I => \N__11682\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__11723\,
            I => \N__11682\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__11720\,
            I => \N__11682\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__11717\,
            I => \N__11682\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__11714\,
            I => \N__11682\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__11711\,
            I => \N__11682\
        );

    \I__2789\ : CascadeMux
    port map (
            O => \N__11710\,
            I => \N__11679\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__11707\,
            I => \N__11676\
        );

    \I__2787\ : InMux
    port map (
            O => \N__11706\,
            I => \N__11671\
        );

    \I__2786\ : InMux
    port map (
            O => \N__11705\,
            I => \N__11671\
        );

    \I__2785\ : Span4Mux_v
    port map (
            O => \N__11702\,
            I => \N__11668\
        );

    \I__2784\ : InMux
    port map (
            O => \N__11701\,
            I => \N__11665\
        );

    \I__2783\ : InMux
    port map (
            O => \N__11700\,
            I => \N__11662\
        );

    \I__2782\ : Span4Mux_h
    port map (
            O => \N__11695\,
            I => \N__11657\
        );

    \I__2781\ : Span4Mux_v
    port map (
            O => \N__11682\,
            I => \N__11657\
        );

    \I__2780\ : InMux
    port map (
            O => \N__11679\,
            I => \N__11654\
        );

    \I__2779\ : Sp12to4
    port map (
            O => \N__11676\,
            I => \N__11651\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__11671\,
            I => \N__11642\
        );

    \I__2777\ : Sp12to4
    port map (
            O => \N__11668\,
            I => \N__11642\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__11665\,
            I => \N__11642\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__11662\,
            I => \N__11642\
        );

    \I__2774\ : Sp12to4
    port map (
            O => \N__11657\,
            I => \N__11637\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__11654\,
            I => \N__11637\
        );

    \I__2772\ : Span12Mux_v
    port map (
            O => \N__11651\,
            I => \N__11634\
        );

    \I__2771\ : Span12Mux_h
    port map (
            O => \N__11642\,
            I => \N__11631\
        );

    \I__2770\ : Span12Mux_h
    port map (
            O => \N__11637\,
            I => \N__11628\
        );

    \I__2769\ : Span12Mux_h
    port map (
            O => \N__11634\,
            I => \N__11623\
        );

    \I__2768\ : Span12Mux_v
    port map (
            O => \N__11631\,
            I => \N__11623\
        );

    \I__2767\ : Span12Mux_v
    port map (
            O => \N__11628\,
            I => \N__11620\
        );

    \I__2766\ : Odrv12
    port map (
            O => \N__11623\,
            I => \AGNUS_REV_c\
        );

    \I__2765\ : Odrv12
    port map (
            O => \N__11620\,
            I => \AGNUS_REV_c\
        );

    \I__2764\ : InMux
    port map (
            O => \N__11615\,
            I => \N__11612\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__11612\,
            I => \N__11609\
        );

    \I__2762\ : Span4Mux_v
    port map (
            O => \N__11609\,
            I => \N__11606\
        );

    \I__2761\ : Odrv4
    port map (
            O => \N__11606\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2760\ : ClkMux
    port map (
            O => \N__11603\,
            I => \N__11579\
        );

    \I__2759\ : ClkMux
    port map (
            O => \N__11602\,
            I => \N__11579\
        );

    \I__2758\ : ClkMux
    port map (
            O => \N__11601\,
            I => \N__11579\
        );

    \I__2757\ : ClkMux
    port map (
            O => \N__11600\,
            I => \N__11579\
        );

    \I__2756\ : ClkMux
    port map (
            O => \N__11599\,
            I => \N__11579\
        );

    \I__2755\ : ClkMux
    port map (
            O => \N__11598\,
            I => \N__11579\
        );

    \I__2754\ : ClkMux
    port map (
            O => \N__11597\,
            I => \N__11579\
        );

    \I__2753\ : ClkMux
    port map (
            O => \N__11596\,
            I => \N__11579\
        );

    \I__2752\ : GlobalMux
    port map (
            O => \N__11579\,
            I => \N__11576\
        );

    \I__2751\ : gio2CtrlBuf
    port map (
            O => \N__11576\,
            I => \C3_c_g\
        );

    \I__2750\ : CEMux
    port map (
            O => \N__11573\,
            I => \N__11528\
        );

    \I__2749\ : CEMux
    port map (
            O => \N__11572\,
            I => \N__11528\
        );

    \I__2748\ : CEMux
    port map (
            O => \N__11571\,
            I => \N__11528\
        );

    \I__2747\ : CEMux
    port map (
            O => \N__11570\,
            I => \N__11528\
        );

    \I__2746\ : CEMux
    port map (
            O => \N__11569\,
            I => \N__11528\
        );

    \I__2745\ : CEMux
    port map (
            O => \N__11568\,
            I => \N__11528\
        );

    \I__2744\ : CEMux
    port map (
            O => \N__11567\,
            I => \N__11528\
        );

    \I__2743\ : CEMux
    port map (
            O => \N__11566\,
            I => \N__11528\
        );

    \I__2742\ : CEMux
    port map (
            O => \N__11565\,
            I => \N__11528\
        );

    \I__2741\ : CEMux
    port map (
            O => \N__11564\,
            I => \N__11528\
        );

    \I__2740\ : CEMux
    port map (
            O => \N__11563\,
            I => \N__11528\
        );

    \I__2739\ : CEMux
    port map (
            O => \N__11562\,
            I => \N__11528\
        );

    \I__2738\ : CEMux
    port map (
            O => \N__11561\,
            I => \N__11528\
        );

    \I__2737\ : CEMux
    port map (
            O => \N__11560\,
            I => \N__11528\
        );

    \I__2736\ : CEMux
    port map (
            O => \N__11559\,
            I => \N__11528\
        );

    \I__2735\ : GlobalMux
    port map (
            O => \N__11528\,
            I => \N__11525\
        );

    \I__2734\ : gio2CtrlBuf
    port map (
            O => \N__11525\,
            I => \DBRn_c_i_0_g\
        );

    \I__2733\ : InMux
    port map (
            O => \N__11522\,
            I => \N__11518\
        );

    \I__2732\ : InMux
    port map (
            O => \N__11521\,
            I => \N__11515\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__11518\,
            I => \N__11512\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__11515\,
            I => \N__11509\
        );

    \I__2729\ : Span4Mux_v
    port map (
            O => \N__11512\,
            I => \N__11504\
        );

    \I__2728\ : Span4Mux_v
    port map (
            O => \N__11509\,
            I => \N__11504\
        );

    \I__2727\ : Sp12to4
    port map (
            O => \N__11504\,
            I => \N__11501\
        );

    \I__2726\ : Odrv12
    port map (
            O => \N__11501\,
            I => \RAS0n_c\
        );

    \I__2725\ : InMux
    port map (
            O => \N__11498\,
            I => \N__11495\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__11495\,
            I => \N__11492\
        );

    \I__2723\ : Span12Mux_h
    port map (
            O => \N__11492\,
            I => \N__11489\
        );

    \I__2722\ : Odrv12
    port map (
            O => \N__11489\,
            I => \RAS1n_c\
        );

    \I__2721\ : InMux
    port map (
            O => \N__11486\,
            I => \N__11483\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__11483\,
            I => \N__11480\
        );

    \I__2719\ : Span12Mux_h
    port map (
            O => \N__11480\,
            I => \N__11477\
        );

    \I__2718\ : Odrv12
    port map (
            O => \N__11477\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2717\ : InMux
    port map (
            O => \N__11474\,
            I => \N__11471\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__11471\,
            I => \N__11432\
        );

    \I__2715\ : ClkMux
    port map (
            O => \N__11470\,
            I => \N__11330\
        );

    \I__2714\ : ClkMux
    port map (
            O => \N__11469\,
            I => \N__11330\
        );

    \I__2713\ : ClkMux
    port map (
            O => \N__11468\,
            I => \N__11330\
        );

    \I__2712\ : ClkMux
    port map (
            O => \N__11467\,
            I => \N__11330\
        );

    \I__2711\ : ClkMux
    port map (
            O => \N__11466\,
            I => \N__11330\
        );

    \I__2710\ : ClkMux
    port map (
            O => \N__11465\,
            I => \N__11330\
        );

    \I__2709\ : ClkMux
    port map (
            O => \N__11464\,
            I => \N__11330\
        );

    \I__2708\ : ClkMux
    port map (
            O => \N__11463\,
            I => \N__11330\
        );

    \I__2707\ : ClkMux
    port map (
            O => \N__11462\,
            I => \N__11330\
        );

    \I__2706\ : ClkMux
    port map (
            O => \N__11461\,
            I => \N__11330\
        );

    \I__2705\ : ClkMux
    port map (
            O => \N__11460\,
            I => \N__11330\
        );

    \I__2704\ : ClkMux
    port map (
            O => \N__11459\,
            I => \N__11330\
        );

    \I__2703\ : ClkMux
    port map (
            O => \N__11458\,
            I => \N__11330\
        );

    \I__2702\ : ClkMux
    port map (
            O => \N__11457\,
            I => \N__11330\
        );

    \I__2701\ : ClkMux
    port map (
            O => \N__11456\,
            I => \N__11330\
        );

    \I__2700\ : ClkMux
    port map (
            O => \N__11455\,
            I => \N__11330\
        );

    \I__2699\ : ClkMux
    port map (
            O => \N__11454\,
            I => \N__11330\
        );

    \I__2698\ : ClkMux
    port map (
            O => \N__11453\,
            I => \N__11330\
        );

    \I__2697\ : ClkMux
    port map (
            O => \N__11452\,
            I => \N__11330\
        );

    \I__2696\ : ClkMux
    port map (
            O => \N__11451\,
            I => \N__11330\
        );

    \I__2695\ : ClkMux
    port map (
            O => \N__11450\,
            I => \N__11330\
        );

    \I__2694\ : ClkMux
    port map (
            O => \N__11449\,
            I => \N__11330\
        );

    \I__2693\ : ClkMux
    port map (
            O => \N__11448\,
            I => \N__11330\
        );

    \I__2692\ : ClkMux
    port map (
            O => \N__11447\,
            I => \N__11330\
        );

    \I__2691\ : ClkMux
    port map (
            O => \N__11446\,
            I => \N__11330\
        );

    \I__2690\ : ClkMux
    port map (
            O => \N__11445\,
            I => \N__11330\
        );

    \I__2689\ : ClkMux
    port map (
            O => \N__11444\,
            I => \N__11330\
        );

    \I__2688\ : ClkMux
    port map (
            O => \N__11443\,
            I => \N__11330\
        );

    \I__2687\ : ClkMux
    port map (
            O => \N__11442\,
            I => \N__11330\
        );

    \I__2686\ : ClkMux
    port map (
            O => \N__11441\,
            I => \N__11330\
        );

    \I__2685\ : ClkMux
    port map (
            O => \N__11440\,
            I => \N__11330\
        );

    \I__2684\ : ClkMux
    port map (
            O => \N__11439\,
            I => \N__11330\
        );

    \I__2683\ : ClkMux
    port map (
            O => \N__11438\,
            I => \N__11330\
        );

    \I__2682\ : ClkMux
    port map (
            O => \N__11437\,
            I => \N__11330\
        );

    \I__2681\ : ClkMux
    port map (
            O => \N__11436\,
            I => \N__11330\
        );

    \I__2680\ : ClkMux
    port map (
            O => \N__11435\,
            I => \N__11330\
        );

    \I__2679\ : Glb2LocalMux
    port map (
            O => \N__11432\,
            I => \N__11330\
        );

    \I__2678\ : ClkMux
    port map (
            O => \N__11431\,
            I => \N__11330\
        );

    \I__2677\ : ClkMux
    port map (
            O => \N__11430\,
            I => \N__11330\
        );

    \I__2676\ : ClkMux
    port map (
            O => \N__11429\,
            I => \N__11330\
        );

    \I__2675\ : ClkMux
    port map (
            O => \N__11428\,
            I => \N__11330\
        );

    \I__2674\ : ClkMux
    port map (
            O => \N__11427\,
            I => \N__11330\
        );

    \I__2673\ : ClkMux
    port map (
            O => \N__11426\,
            I => \N__11330\
        );

    \I__2672\ : ClkMux
    port map (
            O => \N__11425\,
            I => \N__11330\
        );

    \I__2671\ : ClkMux
    port map (
            O => \N__11424\,
            I => \N__11330\
        );

    \I__2670\ : ClkMux
    port map (
            O => \N__11423\,
            I => \N__11330\
        );

    \I__2669\ : GlobalMux
    port map (
            O => \N__11330\,
            I => \CLK80_PLL\
        );

    \I__2668\ : InMux
    port map (
            O => \N__11327\,
            I => \N__11320\
        );

    \I__2667\ : InMux
    port map (
            O => \N__11326\,
            I => \N__11317\
        );

    \I__2666\ : InMux
    port map (
            O => \N__11325\,
            I => \N__11314\
        );

    \I__2665\ : InMux
    port map (
            O => \N__11324\,
            I => \N__11311\
        );

    \I__2664\ : InMux
    port map (
            O => \N__11323\,
            I => \N__11308\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__11320\,
            I => \N__11303\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__11317\,
            I => \N__11272\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__11314\,
            I => \N__11269\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__11311\,
            I => \N__11251\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__11308\,
            I => \N__11247\
        );

    \I__2658\ : SRMux
    port map (
            O => \N__11307\,
            I => \N__11135\
        );

    \I__2657\ : SRMux
    port map (
            O => \N__11306\,
            I => \N__11135\
        );

    \I__2656\ : Glb2LocalMux
    port map (
            O => \N__11303\,
            I => \N__11135\
        );

    \I__2655\ : SRMux
    port map (
            O => \N__11302\,
            I => \N__11135\
        );

    \I__2654\ : SRMux
    port map (
            O => \N__11301\,
            I => \N__11135\
        );

    \I__2653\ : SRMux
    port map (
            O => \N__11300\,
            I => \N__11135\
        );

    \I__2652\ : SRMux
    port map (
            O => \N__11299\,
            I => \N__11135\
        );

    \I__2651\ : SRMux
    port map (
            O => \N__11298\,
            I => \N__11135\
        );

    \I__2650\ : SRMux
    port map (
            O => \N__11297\,
            I => \N__11135\
        );

    \I__2649\ : SRMux
    port map (
            O => \N__11296\,
            I => \N__11135\
        );

    \I__2648\ : SRMux
    port map (
            O => \N__11295\,
            I => \N__11135\
        );

    \I__2647\ : SRMux
    port map (
            O => \N__11294\,
            I => \N__11135\
        );

    \I__2646\ : SRMux
    port map (
            O => \N__11293\,
            I => \N__11135\
        );

    \I__2645\ : SRMux
    port map (
            O => \N__11292\,
            I => \N__11135\
        );

    \I__2644\ : SRMux
    port map (
            O => \N__11291\,
            I => \N__11135\
        );

    \I__2643\ : SRMux
    port map (
            O => \N__11290\,
            I => \N__11135\
        );

    \I__2642\ : SRMux
    port map (
            O => \N__11289\,
            I => \N__11135\
        );

    \I__2641\ : SRMux
    port map (
            O => \N__11288\,
            I => \N__11135\
        );

    \I__2640\ : SRMux
    port map (
            O => \N__11287\,
            I => \N__11135\
        );

    \I__2639\ : SRMux
    port map (
            O => \N__11286\,
            I => \N__11135\
        );

    \I__2638\ : SRMux
    port map (
            O => \N__11285\,
            I => \N__11135\
        );

    \I__2637\ : SRMux
    port map (
            O => \N__11284\,
            I => \N__11135\
        );

    \I__2636\ : SRMux
    port map (
            O => \N__11283\,
            I => \N__11135\
        );

    \I__2635\ : SRMux
    port map (
            O => \N__11282\,
            I => \N__11135\
        );

    \I__2634\ : SRMux
    port map (
            O => \N__11281\,
            I => \N__11135\
        );

    \I__2633\ : SRMux
    port map (
            O => \N__11280\,
            I => \N__11135\
        );

    \I__2632\ : SRMux
    port map (
            O => \N__11279\,
            I => \N__11135\
        );

    \I__2631\ : SRMux
    port map (
            O => \N__11278\,
            I => \N__11135\
        );

    \I__2630\ : SRMux
    port map (
            O => \N__11277\,
            I => \N__11135\
        );

    \I__2629\ : SRMux
    port map (
            O => \N__11276\,
            I => \N__11135\
        );

    \I__2628\ : SRMux
    port map (
            O => \N__11275\,
            I => \N__11135\
        );

    \I__2627\ : Glb2LocalMux
    port map (
            O => \N__11272\,
            I => \N__11135\
        );

    \I__2626\ : Glb2LocalMux
    port map (
            O => \N__11269\,
            I => \N__11135\
        );

    \I__2625\ : SRMux
    port map (
            O => \N__11268\,
            I => \N__11135\
        );

    \I__2624\ : SRMux
    port map (
            O => \N__11267\,
            I => \N__11135\
        );

    \I__2623\ : SRMux
    port map (
            O => \N__11266\,
            I => \N__11135\
        );

    \I__2622\ : SRMux
    port map (
            O => \N__11265\,
            I => \N__11135\
        );

    \I__2621\ : SRMux
    port map (
            O => \N__11264\,
            I => \N__11135\
        );

    \I__2620\ : SRMux
    port map (
            O => \N__11263\,
            I => \N__11135\
        );

    \I__2619\ : SRMux
    port map (
            O => \N__11262\,
            I => \N__11135\
        );

    \I__2618\ : SRMux
    port map (
            O => \N__11261\,
            I => \N__11135\
        );

    \I__2617\ : SRMux
    port map (
            O => \N__11260\,
            I => \N__11135\
        );

    \I__2616\ : SRMux
    port map (
            O => \N__11259\,
            I => \N__11135\
        );

    \I__2615\ : SRMux
    port map (
            O => \N__11258\,
            I => \N__11135\
        );

    \I__2614\ : SRMux
    port map (
            O => \N__11257\,
            I => \N__11135\
        );

    \I__2613\ : SRMux
    port map (
            O => \N__11256\,
            I => \N__11135\
        );

    \I__2612\ : SRMux
    port map (
            O => \N__11255\,
            I => \N__11135\
        );

    \I__2611\ : SRMux
    port map (
            O => \N__11254\,
            I => \N__11135\
        );

    \I__2610\ : Glb2LocalMux
    port map (
            O => \N__11251\,
            I => \N__11135\
        );

    \I__2609\ : SRMux
    port map (
            O => \N__11250\,
            I => \N__11135\
        );

    \I__2608\ : Glb2LocalMux
    port map (
            O => \N__11247\,
            I => \N__11135\
        );

    \I__2607\ : SRMux
    port map (
            O => \N__11246\,
            I => \N__11135\
        );

    \I__2606\ : SRMux
    port map (
            O => \N__11245\,
            I => \N__11135\
        );

    \I__2605\ : SRMux
    port map (
            O => \N__11244\,
            I => \N__11135\
        );

    \I__2604\ : GlobalMux
    port map (
            O => \N__11135\,
            I => \N__11132\
        );

    \I__2603\ : gio2CtrlBuf
    port map (
            O => \N__11132\,
            I => \RESETn_c_i_g\
        );

    \I__2602\ : InMux
    port map (
            O => \N__11129\,
            I => \N__11126\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__11126\,
            I => \N__11123\
        );

    \I__2600\ : Sp12to4
    port map (
            O => \N__11123\,
            I => \N__11119\
        );

    \I__2599\ : InMux
    port map (
            O => \N__11122\,
            I => \N__11116\
        );

    \I__2598\ : Span12Mux_v
    port map (
            O => \N__11119\,
            I => \N__11113\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__11116\,
            I => \N__11110\
        );

    \I__2596\ : Span12Mux_h
    port map (
            O => \N__11113\,
            I => \N__11105\
        );

    \I__2595\ : Span12Mux_v
    port map (
            O => \N__11110\,
            I => \N__11102\
        );

    \I__2594\ : InMux
    port map (
            O => \N__11109\,
            I => \N__11099\
        );

    \I__2593\ : InMux
    port map (
            O => \N__11108\,
            I => \N__11096\
        );

    \I__2592\ : Odrv12
    port map (
            O => \N__11105\,
            I => \REG_CYCLEm\
        );

    \I__2591\ : Odrv12
    port map (
            O => \N__11102\,
            I => \REG_CYCLEm\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__11099\,
            I => \REG_CYCLEm\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__11096\,
            I => \REG_CYCLEm\
        );

    \I__2588\ : InMux
    port map (
            O => \N__11087\,
            I => \N__11084\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__11084\,
            I => \N__11081\
        );

    \I__2586\ : Span4Mux_v
    port map (
            O => \N__11081\,
            I => \N__11077\
        );

    \I__2585\ : CascadeMux
    port map (
            O => \N__11080\,
            I => \N__11073\
        );

    \I__2584\ : Span4Mux_h
    port map (
            O => \N__11077\,
            I => \N__11067\
        );

    \I__2583\ : InMux
    port map (
            O => \N__11076\,
            I => \N__11057\
        );

    \I__2582\ : InMux
    port map (
            O => \N__11073\,
            I => \N__11052\
        );

    \I__2581\ : InMux
    port map (
            O => \N__11072\,
            I => \N__11052\
        );

    \I__2580\ : InMux
    port map (
            O => \N__11071\,
            I => \N__11047\
        );

    \I__2579\ : InMux
    port map (
            O => \N__11070\,
            I => \N__11047\
        );

    \I__2578\ : Span4Mux_h
    port map (
            O => \N__11067\,
            I => \N__11040\
        );

    \I__2577\ : InMux
    port map (
            O => \N__11066\,
            I => \N__11031\
        );

    \I__2576\ : InMux
    port map (
            O => \N__11065\,
            I => \N__11031\
        );

    \I__2575\ : InMux
    port map (
            O => \N__11064\,
            I => \N__11031\
        );

    \I__2574\ : InMux
    port map (
            O => \N__11063\,
            I => \N__11031\
        );

    \I__2573\ : CascadeMux
    port map (
            O => \N__11062\,
            I => \N__11026\
        );

    \I__2572\ : CascadeMux
    port map (
            O => \N__11061\,
            I => \N__11023\
        );

    \I__2571\ : InMux
    port map (
            O => \N__11060\,
            I => \N__11019\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__11057\,
            I => \N__11016\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__11052\,
            I => \N__11013\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__11047\,
            I => \N__11010\
        );

    \I__2567\ : InMux
    port map (
            O => \N__11046\,
            I => \N__11005\
        );

    \I__2566\ : InMux
    port map (
            O => \N__11045\,
            I => \N__11005\
        );

    \I__2565\ : CascadeMux
    port map (
            O => \N__11044\,
            I => \N__11001\
        );

    \I__2564\ : InMux
    port map (
            O => \N__11043\,
            I => \N__10995\
        );

    \I__2563\ : Span4Mux_v
    port map (
            O => \N__11040\,
            I => \N__10987\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__11031\,
            I => \N__10987\
        );

    \I__2561\ : InMux
    port map (
            O => \N__11030\,
            I => \N__10984\
        );

    \I__2560\ : InMux
    port map (
            O => \N__11029\,
            I => \N__10981\
        );

    \I__2559\ : InMux
    port map (
            O => \N__11026\,
            I => \N__10976\
        );

    \I__2558\ : InMux
    port map (
            O => \N__11023\,
            I => \N__10976\
        );

    \I__2557\ : InMux
    port map (
            O => \N__11022\,
            I => \N__10973\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__11019\,
            I => \N__10970\
        );

    \I__2555\ : Span4Mux_v
    port map (
            O => \N__11016\,
            I => \N__10961\
        );

    \I__2554\ : Span4Mux_h
    port map (
            O => \N__11013\,
            I => \N__10961\
        );

    \I__2553\ : Span4Mux_v
    port map (
            O => \N__11010\,
            I => \N__10961\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__11005\,
            I => \N__10961\
        );

    \I__2551\ : InMux
    port map (
            O => \N__11004\,
            I => \N__10958\
        );

    \I__2550\ : InMux
    port map (
            O => \N__11001\,
            I => \N__10955\
        );

    \I__2549\ : InMux
    port map (
            O => \N__11000\,
            I => \N__10948\
        );

    \I__2548\ : InMux
    port map (
            O => \N__10999\,
            I => \N__10948\
        );

    \I__2547\ : InMux
    port map (
            O => \N__10998\,
            I => \N__10948\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__10995\,
            I => \N__10945\
        );

    \I__2545\ : InMux
    port map (
            O => \N__10994\,
            I => \N__10940\
        );

    \I__2544\ : InMux
    port map (
            O => \N__10993\,
            I => \N__10940\
        );

    \I__2543\ : InMux
    port map (
            O => \N__10992\,
            I => \N__10934\
        );

    \I__2542\ : Span4Mux_h
    port map (
            O => \N__10987\,
            I => \N__10929\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__10984\,
            I => \N__10929\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__10981\,
            I => \N__10916\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__10976\,
            I => \N__10916\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__10973\,
            I => \N__10916\
        );

    \I__2537\ : Span4Mux_h
    port map (
            O => \N__10970\,
            I => \N__10916\
        );

    \I__2536\ : Span4Mux_h
    port map (
            O => \N__10961\,
            I => \N__10916\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__10958\,
            I => \N__10916\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__10955\,
            I => \N__10908\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__10948\,
            I => \N__10908\
        );

    \I__2532\ : Span4Mux_v
    port map (
            O => \N__10945\,
            I => \N__10908\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__10940\,
            I => \N__10905\
        );

    \I__2530\ : InMux
    port map (
            O => \N__10939\,
            I => \N__10898\
        );

    \I__2529\ : InMux
    port map (
            O => \N__10938\,
            I => \N__10898\
        );

    \I__2528\ : InMux
    port map (
            O => \N__10937\,
            I => \N__10898\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__10934\,
            I => \N__10895\
        );

    \I__2526\ : Span4Mux_v
    port map (
            O => \N__10929\,
            I => \N__10890\
        );

    \I__2525\ : Span4Mux_v
    port map (
            O => \N__10916\,
            I => \N__10890\
        );

    \I__2524\ : InMux
    port map (
            O => \N__10915\,
            I => \N__10887\
        );

    \I__2523\ : Span4Mux_h
    port map (
            O => \N__10908\,
            I => \N__10880\
        );

    \I__2522\ : Span4Mux_v
    port map (
            O => \N__10905\,
            I => \N__10880\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__10898\,
            I => \N__10880\
        );

    \I__2520\ : Odrv4
    port map (
            O => \N__10895\,
            I => \U712_CHIP_RAM.CPU_CYCLEm\
        );

    \I__2519\ : Odrv4
    port map (
            O => \N__10890\,
            I => \U712_CHIP_RAM.CPU_CYCLEm\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__10887\,
            I => \U712_CHIP_RAM.CPU_CYCLEm\
        );

    \I__2517\ : Odrv4
    port map (
            O => \N__10880\,
            I => \U712_CHIP_RAM.CPU_CYCLEm\
        );

    \I__2516\ : IoInMux
    port map (
            O => \N__10871\,
            I => \N__10868\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__10868\,
            I => \N__10865\
        );

    \I__2514\ : Span4Mux_s3_v
    port map (
            O => \N__10865\,
            I => \N__10862\
        );

    \I__2513\ : Span4Mux_v
    port map (
            O => \N__10862\,
            I => \N__10859\
        );

    \I__2512\ : Odrv4
    port map (
            O => \N__10859\,
            I => \N_338_mux\
        );

    \I__2511\ : InMux
    port map (
            O => \N__10856\,
            I => \N__10853\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__10853\,
            I => \N__10849\
        );

    \I__2509\ : InMux
    port map (
            O => \N__10852\,
            I => \N__10846\
        );

    \I__2508\ : Span4Mux_h
    port map (
            O => \N__10849\,
            I => \N__10840\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__10846\,
            I => \N__10840\
        );

    \I__2506\ : InMux
    port map (
            O => \N__10845\,
            I => \N__10837\
        );

    \I__2505\ : Span4Mux_v
    port map (
            O => \N__10840\,
            I => \N__10831\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__10837\,
            I => \N__10831\
        );

    \I__2503\ : CascadeMux
    port map (
            O => \N__10836\,
            I => \N__10827\
        );

    \I__2502\ : Sp12to4
    port map (
            O => \N__10831\,
            I => \N__10824\
        );

    \I__2501\ : InMux
    port map (
            O => \N__10830\,
            I => \N__10819\
        );

    \I__2500\ : InMux
    port map (
            O => \N__10827\,
            I => \N__10819\
        );

    \I__2499\ : Span12Mux_v
    port map (
            O => \N__10824\,
            I => \N__10816\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__10819\,
            I => \N__10813\
        );

    \I__2497\ : Span12Mux_h
    port map (
            O => \N__10816\,
            I => \N__10810\
        );

    \I__2496\ : Span12Mux_v
    port map (
            O => \N__10813\,
            I => \N__10807\
        );

    \I__2495\ : Odrv12
    port map (
            O => \N__10810\,
            I => \CASLn_c\
        );

    \I__2494\ : Odrv12
    port map (
            O => \N__10807\,
            I => \CASLn_c\
        );

    \I__2493\ : InMux
    port map (
            O => \N__10802\,
            I => \N__10798\
        );

    \I__2492\ : InMux
    port map (
            O => \N__10801\,
            I => \N__10795\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__10798\,
            I => \N__10789\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__10795\,
            I => \N__10786\
        );

    \I__2489\ : InMux
    port map (
            O => \N__10794\,
            I => \N__10781\
        );

    \I__2488\ : InMux
    port map (
            O => \N__10793\,
            I => \N__10781\
        );

    \I__2487\ : InMux
    port map (
            O => \N__10792\,
            I => \N__10778\
        );

    \I__2486\ : Span4Mux_v
    port map (
            O => \N__10789\,
            I => \N__10775\
        );

    \I__2485\ : Span4Mux_v
    port map (
            O => \N__10786\,
            I => \N__10772\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__10781\,
            I => \N__10769\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__10778\,
            I => \N__10766\
        );

    \I__2482\ : Sp12to4
    port map (
            O => \N__10775\,
            I => \N__10763\
        );

    \I__2481\ : Span4Mux_h
    port map (
            O => \N__10772\,
            I => \N__10758\
        );

    \I__2480\ : Span4Mux_v
    port map (
            O => \N__10769\,
            I => \N__10758\
        );

    \I__2479\ : Span4Mux_v
    port map (
            O => \N__10766\,
            I => \N__10755\
        );

    \I__2478\ : Span12Mux_h
    port map (
            O => \N__10763\,
            I => \N__10748\
        );

    \I__2477\ : Sp12to4
    port map (
            O => \N__10758\,
            I => \N__10748\
        );

    \I__2476\ : Sp12to4
    port map (
            O => \N__10755\,
            I => \N__10748\
        );

    \I__2475\ : Span12Mux_h
    port map (
            O => \N__10748\,
            I => \N__10745\
        );

    \I__2474\ : Odrv12
    port map (
            O => \N__10745\,
            I => \RnW_c\
        );

    \I__2473\ : CascadeMux
    port map (
            O => \N__10742\,
            I => \N__10739\
        );

    \I__2472\ : InMux
    port map (
            O => \N__10739\,
            I => \N__10736\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__10736\,
            I => \N__10732\
        );

    \I__2470\ : InMux
    port map (
            O => \N__10735\,
            I => \N__10729\
        );

    \I__2469\ : Sp12to4
    port map (
            O => \N__10732\,
            I => \N__10724\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__10729\,
            I => \N__10724\
        );

    \I__2467\ : Span12Mux_h
    port map (
            O => \N__10724\,
            I => \N__10720\
        );

    \I__2466\ : InMux
    port map (
            O => \N__10723\,
            I => \N__10717\
        );

    \I__2465\ : Odrv12
    port map (
            O => \N__10720\,
            I => \U712_CHIP_RAM.DMA_WRITE_CYCLEZ0\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__10717\,
            I => \U712_CHIP_RAM.DMA_WRITE_CYCLEZ0\
        );

    \I__2463\ : InMux
    port map (
            O => \N__10712\,
            I => \N__10709\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__10709\,
            I => \N__10704\
        );

    \I__2461\ : InMux
    port map (
            O => \N__10708\,
            I => \N__10701\
        );

    \I__2460\ : InMux
    port map (
            O => \N__10707\,
            I => \N__10698\
        );

    \I__2459\ : Span4Mux_v
    port map (
            O => \N__10704\,
            I => \N__10693\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__10701\,
            I => \N__10693\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__10698\,
            I => \N__10690\
        );

    \I__2456\ : Span4Mux_v
    port map (
            O => \N__10693\,
            I => \N__10685\
        );

    \I__2455\ : Span4Mux_h
    port map (
            O => \N__10690\,
            I => \N__10685\
        );

    \I__2454\ : Span4Mux_h
    port map (
            O => \N__10685\,
            I => \N__10680\
        );

    \I__2453\ : InMux
    port map (
            O => \N__10684\,
            I => \N__10675\
        );

    \I__2452\ : InMux
    port map (
            O => \N__10683\,
            I => \N__10675\
        );

    \I__2451\ : Span4Mux_h
    port map (
            O => \N__10680\,
            I => \N__10670\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__10675\,
            I => \N__10670\
        );

    \I__2449\ : Span4Mux_h
    port map (
            O => \N__10670\,
            I => \N__10667\
        );

    \I__2448\ : Span4Mux_v
    port map (
            O => \N__10667\,
            I => \N__10664\
        );

    \I__2447\ : Odrv4
    port map (
            O => \N__10664\,
            I => \CASUn_c\
        );

    \I__2446\ : IoInMux
    port map (
            O => \N__10661\,
            I => \N__10658\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__10658\,
            I => \N__10655\
        );

    \I__2444\ : IoSpan4Mux
    port map (
            O => \N__10655\,
            I => \N__10652\
        );

    \I__2443\ : Span4Mux_s3_h
    port map (
            O => \N__10652\,
            I => \N__10649\
        );

    \I__2442\ : Odrv4
    port map (
            O => \N__10649\,
            I => \N_328_mux\
        );

    \I__2441\ : InMux
    port map (
            O => \N__10646\,
            I => \N__10643\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__10643\,
            I => \N__10639\
        );

    \I__2439\ : InMux
    port map (
            O => \N__10642\,
            I => \N__10636\
        );

    \I__2438\ : Span4Mux_h
    port map (
            O => \N__10639\,
            I => \N__10631\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__10636\,
            I => \N__10631\
        );

    \I__2436\ : Span4Mux_v
    port map (
            O => \N__10631\,
            I => \N__10626\
        );

    \I__2435\ : InMux
    port map (
            O => \N__10630\,
            I => \N__10623\
        );

    \I__2434\ : InMux
    port map (
            O => \N__10629\,
            I => \N__10620\
        );

    \I__2433\ : Span4Mux_v
    port map (
            O => \N__10626\,
            I => \N__10617\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__10623\,
            I => \N__10612\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__10620\,
            I => \N__10612\
        );

    \I__2430\ : Sp12to4
    port map (
            O => \N__10617\,
            I => \N__10607\
        );

    \I__2429\ : Span12Mux_v
    port map (
            O => \N__10612\,
            I => \N__10607\
        );

    \I__2428\ : Span12Mux_h
    port map (
            O => \N__10607\,
            I => \N__10604\
        );

    \I__2427\ : Odrv12
    port map (
            O => \N__10604\,
            I => \DRA_c_6\
        );

    \I__2426\ : InMux
    port map (
            O => \N__10601\,
            I => \N__10598\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__10598\,
            I => \N__10595\
        );

    \I__2424\ : Span4Mux_h
    port map (
            O => \N__10595\,
            I => \N__10592\
        );

    \I__2423\ : Odrv4
    port map (
            O => \N__10592\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__2422\ : InMux
    port map (
            O => \N__10589\,
            I => \N__10586\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__10586\,
            I => \N__10583\
        );

    \I__2420\ : Odrv4
    port map (
            O => \N__10583\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__2419\ : InMux
    port map (
            O => \N__10580\,
            I => \N__10576\
        );

    \I__2418\ : InMux
    port map (
            O => \N__10579\,
            I => \N__10573\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__10576\,
            I => \N__10566\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__10573\,
            I => \N__10566\
        );

    \I__2415\ : InMux
    port map (
            O => \N__10572\,
            I => \N__10563\
        );

    \I__2414\ : InMux
    port map (
            O => \N__10571\,
            I => \N__10560\
        );

    \I__2413\ : Span4Mux_v
    port map (
            O => \N__10566\,
            I => \N__10557\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__10563\,
            I => \N__10552\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__10560\,
            I => \N__10552\
        );

    \I__2410\ : Span4Mux_v
    port map (
            O => \N__10557\,
            I => \N__10549\
        );

    \I__2409\ : Span12Mux_v
    port map (
            O => \N__10552\,
            I => \N__10544\
        );

    \I__2408\ : Sp12to4
    port map (
            O => \N__10549\,
            I => \N__10544\
        );

    \I__2407\ : Span12Mux_h
    port map (
            O => \N__10544\,
            I => \N__10541\
        );

    \I__2406\ : Odrv12
    port map (
            O => \N__10541\,
            I => \DRA_c_3\
        );

    \I__2405\ : InMux
    port map (
            O => \N__10538\,
            I => \N__10535\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__10535\,
            I => \N__10532\
        );

    \I__2403\ : Odrv4
    port map (
            O => \N__10532\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__2402\ : InMux
    port map (
            O => \N__10529\,
            I => \N__10524\
        );

    \I__2401\ : InMux
    port map (
            O => \N__10528\,
            I => \N__10521\
        );

    \I__2400\ : InMux
    port map (
            O => \N__10527\,
            I => \N__10518\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__10524\,
            I => \N__10510\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__10521\,
            I => \N__10510\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__10518\,
            I => \N__10510\
        );

    \I__2396\ : InMux
    port map (
            O => \N__10517\,
            I => \N__10507\
        );

    \I__2395\ : Span4Mux_v
    port map (
            O => \N__10510\,
            I => \N__10504\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__10507\,
            I => \N__10501\
        );

    \I__2393\ : Sp12to4
    port map (
            O => \N__10504\,
            I => \N__10498\
        );

    \I__2392\ : Span4Mux_h
    port map (
            O => \N__10501\,
            I => \N__10495\
        );

    \I__2391\ : Span12Mux_h
    port map (
            O => \N__10498\,
            I => \N__10492\
        );

    \I__2390\ : Sp12to4
    port map (
            O => \N__10495\,
            I => \N__10489\
        );

    \I__2389\ : Span12Mux_v
    port map (
            O => \N__10492\,
            I => \N__10486\
        );

    \I__2388\ : Span12Mux_v
    port map (
            O => \N__10489\,
            I => \N__10483\
        );

    \I__2387\ : Odrv12
    port map (
            O => \N__10486\,
            I => \DRA_c_2\
        );

    \I__2386\ : Odrv12
    port map (
            O => \N__10483\,
            I => \DRA_c_2\
        );

    \I__2385\ : InMux
    port map (
            O => \N__10478\,
            I => \N__10475\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__10475\,
            I => \N__10472\
        );

    \I__2383\ : Span4Mux_h
    port map (
            O => \N__10472\,
            I => \N__10469\
        );

    \I__2382\ : Span4Mux_h
    port map (
            O => \N__10469\,
            I => \N__10466\
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__10466\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__2380\ : InMux
    port map (
            O => \N__10463\,
            I => \N__10460\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__10460\,
            I => \N__10457\
        );

    \I__2378\ : Span4Mux_h
    port map (
            O => \N__10457\,
            I => \N__10454\
        );

    \I__2377\ : Odrv4
    port map (
            O => \N__10454\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2376\ : InMux
    port map (
            O => \N__10451\,
            I => \N__10447\
        );

    \I__2375\ : InMux
    port map (
            O => \N__10450\,
            I => \N__10444\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__10447\,
            I => \N__10441\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__10444\,
            I => \N__10438\
        );

    \I__2372\ : Sp12to4
    port map (
            O => \N__10441\,
            I => \N__10435\
        );

    \I__2371\ : Span12Mux_h
    port map (
            O => \N__10438\,
            I => \N__10432\
        );

    \I__2370\ : Span12Mux_v
    port map (
            O => \N__10435\,
            I => \N__10429\
        );

    \I__2369\ : Span12Mux_v
    port map (
            O => \N__10432\,
            I => \N__10426\
        );

    \I__2368\ : Span12Mux_h
    port map (
            O => \N__10429\,
            I => \N__10423\
        );

    \I__2367\ : Odrv12
    port map (
            O => \N__10426\,
            I => \DRA_c_0\
        );

    \I__2366\ : Odrv12
    port map (
            O => \N__10423\,
            I => \DRA_c_0\
        );

    \I__2365\ : InMux
    port map (
            O => \N__10418\,
            I => \N__10414\
        );

    \I__2364\ : InMux
    port map (
            O => \N__10417\,
            I => \N__10410\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__10414\,
            I => \N__10406\
        );

    \I__2362\ : InMux
    port map (
            O => \N__10413\,
            I => \N__10403\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__10410\,
            I => \N__10400\
        );

    \I__2360\ : InMux
    port map (
            O => \N__10409\,
            I => \N__10397\
        );

    \I__2359\ : Span4Mux_v
    port map (
            O => \N__10406\,
            I => \N__10390\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__10403\,
            I => \N__10390\
        );

    \I__2357\ : Span4Mux_v
    port map (
            O => \N__10400\,
            I => \N__10390\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__10397\,
            I => \N__10387\
        );

    \I__2355\ : Sp12to4
    port map (
            O => \N__10390\,
            I => \N__10384\
        );

    \I__2354\ : Span4Mux_h
    port map (
            O => \N__10387\,
            I => \N__10381\
        );

    \I__2353\ : Span12Mux_h
    port map (
            O => \N__10384\,
            I => \N__10378\
        );

    \I__2352\ : Sp12to4
    port map (
            O => \N__10381\,
            I => \N__10375\
        );

    \I__2351\ : Span12Mux_v
    port map (
            O => \N__10378\,
            I => \N__10372\
        );

    \I__2350\ : Span12Mux_v
    port map (
            O => \N__10375\,
            I => \N__10369\
        );

    \I__2349\ : Odrv12
    port map (
            O => \N__10372\,
            I => \DRA_c_1\
        );

    \I__2348\ : Odrv12
    port map (
            O => \N__10369\,
            I => \DRA_c_1\
        );

    \I__2347\ : InMux
    port map (
            O => \N__10364\,
            I => \N__10361\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__10361\,
            I => \N__10358\
        );

    \I__2345\ : Span4Mux_h
    port map (
            O => \N__10358\,
            I => \N__10355\
        );

    \I__2344\ : Odrv4
    port map (
            O => \N__10355\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__2343\ : CascadeMux
    port map (
            O => \N__10352\,
            I => \N__10347\
        );

    \I__2342\ : InMux
    port map (
            O => \N__10351\,
            I => \N__10344\
        );

    \I__2341\ : InMux
    port map (
            O => \N__10350\,
            I => \N__10341\
        );

    \I__2340\ : InMux
    port map (
            O => \N__10347\,
            I => \N__10338\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__10344\,
            I => \N__10332\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__10341\,
            I => \N__10332\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__10338\,
            I => \N__10327\
        );

    \I__2336\ : InMux
    port map (
            O => \N__10337\,
            I => \N__10324\
        );

    \I__2335\ : Span4Mux_v
    port map (
            O => \N__10332\,
            I => \N__10321\
        );

    \I__2334\ : InMux
    port map (
            O => \N__10331\,
            I => \N__10318\
        );

    \I__2333\ : InMux
    port map (
            O => \N__10330\,
            I => \N__10315\
        );

    \I__2332\ : Span4Mux_v
    port map (
            O => \N__10327\,
            I => \N__10312\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__10324\,
            I => \N__10309\
        );

    \I__2330\ : Odrv4
    port map (
            O => \N__10321\,
            I => \U712_CHIP_RAM.DMA_CYCLEm\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__10318\,
            I => \U712_CHIP_RAM.DMA_CYCLEm\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__10315\,
            I => \U712_CHIP_RAM.DMA_CYCLEm\
        );

    \I__2327\ : Odrv4
    port map (
            O => \N__10312\,
            I => \U712_CHIP_RAM.DMA_CYCLEm\
        );

    \I__2326\ : Odrv4
    port map (
            O => \N__10309\,
            I => \U712_CHIP_RAM.DMA_CYCLEm\
        );

    \I__2325\ : InMux
    port map (
            O => \N__10298\,
            I => \N__10292\
        );

    \I__2324\ : InMux
    port map (
            O => \N__10297\,
            I => \N__10292\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__10292\,
            I => \U712_CHIP_RAM.N_345\
        );

    \I__2322\ : InMux
    port map (
            O => \N__10289\,
            I => \N__10286\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__10286\,
            I => \N__10283\
        );

    \I__2320\ : Odrv4
    port map (
            O => \N__10283\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__2319\ : InMux
    port map (
            O => \N__10280\,
            I => \N__10277\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__10277\,
            I => \U712_CHIP_RAM.N_346\
        );

    \I__2317\ : IoInMux
    port map (
            O => \N__10274\,
            I => \N__10271\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__10271\,
            I => \N__10268\
        );

    \I__2315\ : IoSpan4Mux
    port map (
            O => \N__10268\,
            I => \N__10265\
        );

    \I__2314\ : Sp12to4
    port map (
            O => \N__10265\,
            I => \N__10259\
        );

    \I__2313\ : CascadeMux
    port map (
            O => \N__10264\,
            I => \N__10256\
        );

    \I__2312\ : CascadeMux
    port map (
            O => \N__10263\,
            I => \N__10253\
        );

    \I__2311\ : CascadeMux
    port map (
            O => \N__10262\,
            I => \N__10249\
        );

    \I__2310\ : Span12Mux_s7_v
    port map (
            O => \N__10259\,
            I => \N__10246\
        );

    \I__2309\ : InMux
    port map (
            O => \N__10256\,
            I => \N__10243\
        );

    \I__2308\ : InMux
    port map (
            O => \N__10253\,
            I => \N__10236\
        );

    \I__2307\ : InMux
    port map (
            O => \N__10252\,
            I => \N__10236\
        );

    \I__2306\ : InMux
    port map (
            O => \N__10249\,
            I => \N__10236\
        );

    \I__2305\ : Span12Mux_h
    port map (
            O => \N__10246\,
            I => \N__10232\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__10243\,
            I => \N__10227\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__10236\,
            I => \N__10227\
        );

    \I__2302\ : InMux
    port map (
            O => \N__10235\,
            I => \N__10224\
        );

    \I__2301\ : Odrv12
    port map (
            O => \N__10232\,
            I => \DBENn_c\
        );

    \I__2300\ : Odrv4
    port map (
            O => \N__10227\,
            I => \DBENn_c\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__10224\,
            I => \DBENn_c\
        );

    \I__2298\ : CascadeMux
    port map (
            O => \N__10217\,
            I => \U712_CHIP_RAM.N_346_cascade_\
        );

    \I__2297\ : IoInMux
    port map (
            O => \N__10214\,
            I => \N__10211\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__10211\,
            I => \N__10208\
        );

    \I__2295\ : IoSpan4Mux
    port map (
            O => \N__10208\,
            I => \N__10205\
        );

    \I__2294\ : Sp12to4
    port map (
            O => \N__10205\,
            I => \N__10202\
        );

    \I__2293\ : Span12Mux_s7_v
    port map (
            O => \N__10202\,
            I => \N__10199\
        );

    \I__2292\ : Span12Mux_v
    port map (
            O => \N__10199\,
            I => \N__10196\
        );

    \I__2291\ : Odrv12
    port map (
            O => \N__10196\,
            I => \CLLBEn_c\
        );

    \I__2290\ : IoInMux
    port map (
            O => \N__10193\,
            I => \N__10190\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__10190\,
            I => \N__10187\
        );

    \I__2288\ : IoSpan4Mux
    port map (
            O => \N__10187\,
            I => \N__10183\
        );

    \I__2287\ : InMux
    port map (
            O => \N__10186\,
            I => \N__10180\
        );

    \I__2286\ : Sp12to4
    port map (
            O => \N__10183\,
            I => \N__10177\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__10180\,
            I => \N__10174\
        );

    \I__2284\ : Odrv12
    port map (
            O => \N__10177\,
            I => \LLBEn_c\
        );

    \I__2283\ : Odrv4
    port map (
            O => \N__10174\,
            I => \LLBEn_c\
        );

    \I__2282\ : CascadeMux
    port map (
            O => \N__10169\,
            I => \N__10164\
        );

    \I__2281\ : InMux
    port map (
            O => \N__10168\,
            I => \N__10161\
        );

    \I__2280\ : InMux
    port map (
            O => \N__10167\,
            I => \N__10156\
        );

    \I__2279\ : InMux
    port map (
            O => \N__10164\,
            I => \N__10156\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__10161\,
            I => \N__10152\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__10156\,
            I => \N__10149\
        );

    \I__2276\ : InMux
    port map (
            O => \N__10155\,
            I => \N__10146\
        );

    \I__2275\ : Span4Mux_v
    port map (
            O => \N__10152\,
            I => \N__10143\
        );

    \I__2274\ : Span4Mux_v
    port map (
            O => \N__10149\,
            I => \N__10140\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__10146\,
            I => \N__10137\
        );

    \I__2272\ : Sp12to4
    port map (
            O => \N__10143\,
            I => \N__10134\
        );

    \I__2271\ : Span4Mux_h
    port map (
            O => \N__10140\,
            I => \N__10129\
        );

    \I__2270\ : Span4Mux_v
    port map (
            O => \N__10137\,
            I => \N__10129\
        );

    \I__2269\ : Span12Mux_h
    port map (
            O => \N__10134\,
            I => \N__10124\
        );

    \I__2268\ : Sp12to4
    port map (
            O => \N__10129\,
            I => \N__10124\
        );

    \I__2267\ : Odrv12
    port map (
            O => \N__10124\,
            I => \A_c_0\
        );

    \I__2266\ : IoInMux
    port map (
            O => \N__10121\,
            I => \N__10118\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__10118\,
            I => \N__10115\
        );

    \I__2264\ : Span4Mux_s2_v
    port map (
            O => \N__10115\,
            I => \N__10111\
        );

    \I__2263\ : InMux
    port map (
            O => \N__10114\,
            I => \N__10108\
        );

    \I__2262\ : Span4Mux_v
    port map (
            O => \N__10111\,
            I => \N__10105\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__10108\,
            I => \N__10102\
        );

    \I__2260\ : Odrv4
    port map (
            O => \N__10105\,
            I => \UUBEn_c\
        );

    \I__2259\ : Odrv12
    port map (
            O => \N__10102\,
            I => \UUBEn_c\
        );

    \I__2258\ : CascadeMux
    port map (
            O => \N__10097\,
            I => \N__10091\
        );

    \I__2257\ : InMux
    port map (
            O => \N__10096\,
            I => \N__10083\
        );

    \I__2256\ : InMux
    port map (
            O => \N__10095\,
            I => \N__10083\
        );

    \I__2255\ : InMux
    port map (
            O => \N__10094\,
            I => \N__10083\
        );

    \I__2254\ : InMux
    port map (
            O => \N__10091\,
            I => \N__10078\
        );

    \I__2253\ : InMux
    port map (
            O => \N__10090\,
            I => \N__10078\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__10083\,
            I => \N__10074\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__10078\,
            I => \N__10071\
        );

    \I__2250\ : InMux
    port map (
            O => \N__10077\,
            I => \N__10068\
        );

    \I__2249\ : Span4Mux_v
    port map (
            O => \N__10074\,
            I => \N__10065\
        );

    \I__2248\ : Span4Mux_v
    port map (
            O => \N__10071\,
            I => \N__10062\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__10068\,
            I => \N__10059\
        );

    \I__2246\ : Span4Mux_v
    port map (
            O => \N__10065\,
            I => \N__10056\
        );

    \I__2245\ : Span4Mux_h
    port map (
            O => \N__10062\,
            I => \N__10051\
        );

    \I__2244\ : Span4Mux_v
    port map (
            O => \N__10059\,
            I => \N__10051\
        );

    \I__2243\ : Sp12to4
    port map (
            O => \N__10056\,
            I => \N__10048\
        );

    \I__2242\ : Span4Mux_v
    port map (
            O => \N__10051\,
            I => \N__10045\
        );

    \I__2241\ : Span12Mux_h
    port map (
            O => \N__10048\,
            I => \N__10040\
        );

    \I__2240\ : Sp12to4
    port map (
            O => \N__10045\,
            I => \N__10040\
        );

    \I__2239\ : Odrv12
    port map (
            O => \N__10040\,
            I => \SIZ_c_0\
        );

    \I__2238\ : InMux
    port map (
            O => \N__10037\,
            I => \N__10027\
        );

    \I__2237\ : InMux
    port map (
            O => \N__10036\,
            I => \N__10027\
        );

    \I__2236\ : InMux
    port map (
            O => \N__10035\,
            I => \N__10027\
        );

    \I__2235\ : InMux
    port map (
            O => \N__10034\,
            I => \N__10024\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__10027\,
            I => \N__10021\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__10024\,
            I => \N__10018\
        );

    \I__2232\ : Span4Mux_v
    port map (
            O => \N__10021\,
            I => \N__10015\
        );

    \I__2231\ : Span4Mux_v
    port map (
            O => \N__10018\,
            I => \N__10012\
        );

    \I__2230\ : Sp12to4
    port map (
            O => \N__10015\,
            I => \N__10007\
        );

    \I__2229\ : Sp12to4
    port map (
            O => \N__10012\,
            I => \N__10007\
        );

    \I__2228\ : Span12Mux_h
    port map (
            O => \N__10007\,
            I => \N__10004\
        );

    \I__2227\ : Odrv12
    port map (
            O => \N__10004\,
            I => \A_c_1\
        );

    \I__2226\ : CascadeMux
    port map (
            O => \N__10001\,
            I => \N__9996\
        );

    \I__2225\ : CascadeMux
    port map (
            O => \N__10000\,
            I => \N__9993\
        );

    \I__2224\ : CascadeMux
    port map (
            O => \N__9999\,
            I => \N__9990\
        );

    \I__2223\ : InMux
    port map (
            O => \N__9996\,
            I => \N__9984\
        );

    \I__2222\ : InMux
    port map (
            O => \N__9993\,
            I => \N__9979\
        );

    \I__2221\ : InMux
    port map (
            O => \N__9990\,
            I => \N__9979\
        );

    \I__2220\ : InMux
    port map (
            O => \N__9989\,
            I => \N__9974\
        );

    \I__2219\ : InMux
    port map (
            O => \N__9988\,
            I => \N__9974\
        );

    \I__2218\ : InMux
    port map (
            O => \N__9987\,
            I => \N__9971\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__9984\,
            I => \N__9964\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__9979\,
            I => \N__9964\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__9974\,
            I => \N__9964\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__9971\,
            I => \N__9961\
        );

    \I__2213\ : Sp12to4
    port map (
            O => \N__9964\,
            I => \N__9958\
        );

    \I__2212\ : Sp12to4
    port map (
            O => \N__9961\,
            I => \N__9955\
        );

    \I__2211\ : Span12Mux_v
    port map (
            O => \N__9958\,
            I => \N__9952\
        );

    \I__2210\ : Span12Mux_v
    port map (
            O => \N__9955\,
            I => \N__9949\
        );

    \I__2209\ : Span12Mux_h
    port map (
            O => \N__9952\,
            I => \N__9946\
        );

    \I__2208\ : Span12Mux_h
    port map (
            O => \N__9949\,
            I => \N__9943\
        );

    \I__2207\ : Odrv12
    port map (
            O => \N__9946\,
            I => \SIZ_c_1\
        );

    \I__2206\ : Odrv12
    port map (
            O => \N__9943\,
            I => \SIZ_c_1\
        );

    \I__2205\ : InMux
    port map (
            O => \N__9938\,
            I => \N__9933\
        );

    \I__2204\ : InMux
    port map (
            O => \N__9937\,
            I => \N__9928\
        );

    \I__2203\ : InMux
    port map (
            O => \N__9936\,
            I => \N__9928\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__9933\,
            I => \U712_CHIP_RAM.N_325_mux\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__9928\,
            I => \U712_CHIP_RAM.N_325_mux\
        );

    \I__2200\ : IoInMux
    port map (
            O => \N__9923\,
            I => \N__9920\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__9920\,
            I => \N__9917\
        );

    \I__2198\ : IoSpan4Mux
    port map (
            O => \N__9917\,
            I => \N__9914\
        );

    \I__2197\ : Span4Mux_s1_v
    port map (
            O => \N__9914\,
            I => \N__9911\
        );

    \I__2196\ : Span4Mux_h
    port map (
            O => \N__9911\,
            I => \N__9907\
        );

    \I__2195\ : InMux
    port map (
            O => \N__9910\,
            I => \N__9904\
        );

    \I__2194\ : Sp12to4
    port map (
            O => \N__9907\,
            I => \N__9899\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__9904\,
            I => \N__9899\
        );

    \I__2192\ : Odrv12
    port map (
            O => \N__9899\,
            I => \UMBEn_c\
        );

    \I__2191\ : InMux
    port map (
            O => \N__9896\,
            I => \N__9893\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__9893\,
            I => \N__9888\
        );

    \I__2189\ : CascadeMux
    port map (
            O => \N__9892\,
            I => \N__9885\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__9891\,
            I => \N__9881\
        );

    \I__2187\ : Span4Mux_h
    port map (
            O => \N__9888\,
            I => \N__9877\
        );

    \I__2186\ : InMux
    port map (
            O => \N__9885\,
            I => \N__9874\
        );

    \I__2185\ : InMux
    port map (
            O => \N__9884\,
            I => \N__9870\
        );

    \I__2184\ : InMux
    port map (
            O => \N__9881\,
            I => \N__9867\
        );

    \I__2183\ : InMux
    port map (
            O => \N__9880\,
            I => \N__9864\
        );

    \I__2182\ : Span4Mux_v
    port map (
            O => \N__9877\,
            I => \N__9859\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__9874\,
            I => \N__9859\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__9873\,
            I => \N__9856\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__9870\,
            I => \N__9849\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__9867\,
            I => \N__9849\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__9864\,
            I => \N__9846\
        );

    \I__2176\ : Span4Mux_h
    port map (
            O => \N__9859\,
            I => \N__9843\
        );

    \I__2175\ : InMux
    port map (
            O => \N__9856\,
            I => \N__9840\
        );

    \I__2174\ : InMux
    port map (
            O => \N__9855\,
            I => \N__9837\
        );

    \I__2173\ : InMux
    port map (
            O => \N__9854\,
            I => \N__9834\
        );

    \I__2172\ : Odrv4
    port map (
            O => \N__9849\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2171\ : Odrv4
    port map (
            O => \N__9846\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2170\ : Odrv4
    port map (
            O => \N__9843\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__9840\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__9837\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__9834\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2166\ : IoInMux
    port map (
            O => \N__9821\,
            I => \N__9818\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__9818\,
            I => \N__9815\
        );

    \I__2164\ : IoSpan4Mux
    port map (
            O => \N__9815\,
            I => \N__9812\
        );

    \I__2163\ : Sp12to4
    port map (
            O => \N__9812\,
            I => \N__9809\
        );

    \I__2162\ : Span12Mux_s7_v
    port map (
            O => \N__9809\,
            I => \N__9806\
        );

    \I__2161\ : Odrv12
    port map (
            O => \N__9806\,
            I => \WEn_c\
        );

    \I__2160\ : InMux
    port map (
            O => \N__9803\,
            I => \N__9800\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__9800\,
            I => \N__9797\
        );

    \I__2158\ : Odrv4
    port map (
            O => \N__9797\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2157\ : InMux
    port map (
            O => \N__9794\,
            I => \N__9789\
        );

    \I__2156\ : InMux
    port map (
            O => \N__9793\,
            I => \N__9786\
        );

    \I__2155\ : InMux
    port map (
            O => \N__9792\,
            I => \N__9783\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__9789\,
            I => \N__9775\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__9786\,
            I => \N__9775\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__9783\,
            I => \N__9775\
        );

    \I__2151\ : InMux
    port map (
            O => \N__9782\,
            I => \N__9772\
        );

    \I__2150\ : Span4Mux_v
    port map (
            O => \N__9775\,
            I => \N__9767\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__9772\,
            I => \N__9767\
        );

    \I__2148\ : Span4Mux_v
    port map (
            O => \N__9767\,
            I => \N__9764\
        );

    \I__2147\ : Span4Mux_v
    port map (
            O => \N__9764\,
            I => \N__9761\
        );

    \I__2146\ : Sp12to4
    port map (
            O => \N__9761\,
            I => \N__9758\
        );

    \I__2145\ : Span12Mux_h
    port map (
            O => \N__9758\,
            I => \N__9755\
        );

    \I__2144\ : Odrv12
    port map (
            O => \N__9755\,
            I => \DRA_c_4\
        );

    \I__2143\ : InMux
    port map (
            O => \N__9752\,
            I => \N__9749\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__9749\,
            I => \N__9746\
        );

    \I__2141\ : Odrv12
    port map (
            O => \N__9746\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__2140\ : InMux
    port map (
            O => \N__9743\,
            I => \N__9737\
        );

    \I__2139\ : InMux
    port map (
            O => \N__9742\,
            I => \N__9734\
        );

    \I__2138\ : InMux
    port map (
            O => \N__9741\,
            I => \N__9729\
        );

    \I__2137\ : InMux
    port map (
            O => \N__9740\,
            I => \N__9729\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9737\,
            I => \N__9722\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__9734\,
            I => \N__9722\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__9729\,
            I => \N__9722\
        );

    \I__2133\ : Span4Mux_v
    port map (
            O => \N__9722\,
            I => \N__9719\
        );

    \I__2132\ : Sp12to4
    port map (
            O => \N__9719\,
            I => \N__9716\
        );

    \I__2131\ : Span12Mux_h
    port map (
            O => \N__9716\,
            I => \N__9713\
        );

    \I__2130\ : Span12Mux_v
    port map (
            O => \N__9713\,
            I => \N__9710\
        );

    \I__2129\ : Odrv12
    port map (
            O => \N__9710\,
            I => \DRA_c_5\
        );

    \I__2128\ : InMux
    port map (
            O => \N__9707\,
            I => \N__9704\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__9704\,
            I => \N__9701\
        );

    \I__2126\ : Odrv4
    port map (
            O => \N__9701\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__2125\ : InMux
    port map (
            O => \N__9698\,
            I => \N__9695\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__9695\,
            I => \U712_CHIP_RAM.m191_1\
        );

    \I__2123\ : IoInMux
    port map (
            O => \N__9692\,
            I => \N__9689\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__9689\,
            I => \N__9686\
        );

    \I__2121\ : IoSpan4Mux
    port map (
            O => \N__9686\,
            I => \N__9683\
        );

    \I__2120\ : IoSpan4Mux
    port map (
            O => \N__9683\,
            I => \N__9680\
        );

    \I__2119\ : Span4Mux_s3_h
    port map (
            O => \N__9680\,
            I => \N__9677\
        );

    \I__2118\ : Sp12to4
    port map (
            O => \N__9677\,
            I => \N__9674\
        );

    \I__2117\ : Odrv12
    port map (
            O => \N__9674\,
            I => \CMA_c_7\
        );

    \I__2116\ : CEMux
    port map (
            O => \N__9671\,
            I => \N__9668\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__9668\,
            I => \N__9663\
        );

    \I__2114\ : CEMux
    port map (
            O => \N__9667\,
            I => \N__9660\
        );

    \I__2113\ : CEMux
    port map (
            O => \N__9666\,
            I => \N__9657\
        );

    \I__2112\ : Span4Mux_v
    port map (
            O => \N__9663\,
            I => \N__9654\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__9660\,
            I => \N__9651\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__9657\,
            I => \N__9648\
        );

    \I__2109\ : Span4Mux_h
    port map (
            O => \N__9654\,
            I => \N__9642\
        );

    \I__2108\ : Span4Mux_h
    port map (
            O => \N__9651\,
            I => \N__9637\
        );

    \I__2107\ : Span4Mux_h
    port map (
            O => \N__9648\,
            I => \N__9637\
        );

    \I__2106\ : CEMux
    port map (
            O => \N__9647\,
            I => \N__9634\
        );

    \I__2105\ : CEMux
    port map (
            O => \N__9646\,
            I => \N__9631\
        );

    \I__2104\ : CEMux
    port map (
            O => \N__9645\,
            I => \N__9628\
        );

    \I__2103\ : Odrv4
    port map (
            O => \N__9642\,
            I => \U712_CHIP_RAM.N_198_0\
        );

    \I__2102\ : Odrv4
    port map (
            O => \N__9637\,
            I => \U712_CHIP_RAM.N_198_0\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__9634\,
            I => \U712_CHIP_RAM.N_198_0\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__9631\,
            I => \U712_CHIP_RAM.N_198_0\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__9628\,
            I => \U712_CHIP_RAM.N_198_0\
        );

    \I__2098\ : InMux
    port map (
            O => \N__9617\,
            I => \N__9614\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__9614\,
            I => \N__9611\
        );

    \I__2096\ : Odrv12
    port map (
            O => \N__9611\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__2095\ : InMux
    port map (
            O => \N__9608\,
            I => \N__9605\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__9605\,
            I => \N__9602\
        );

    \I__2093\ : Odrv4
    port map (
            O => \N__9602\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__2092\ : InMux
    port map (
            O => \N__9599\,
            I => \N__9596\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__9596\,
            I => \N__9593\
        );

    \I__2090\ : Odrv4
    port map (
            O => \N__9593\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__2089\ : InMux
    port map (
            O => \N__9590\,
            I => \N__9587\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__9587\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__2087\ : InMux
    port map (
            O => \N__9584\,
            I => \N__9581\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__9581\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2085\ : IoInMux
    port map (
            O => \N__9578\,
            I => \N__9575\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__9575\,
            I => \N__9572\
        );

    \I__2083\ : Span4Mux_s2_h
    port map (
            O => \N__9572\,
            I => \N__9569\
        );

    \I__2082\ : Span4Mux_v
    port map (
            O => \N__9569\,
            I => \N__9566\
        );

    \I__2081\ : Sp12to4
    port map (
            O => \N__9566\,
            I => \N__9563\
        );

    \I__2080\ : Span12Mux_h
    port map (
            O => \N__9563\,
            I => \N__9560\
        );

    \I__2079\ : Span12Mux_v
    port map (
            O => \N__9560\,
            I => \N__9557\
        );

    \I__2078\ : Odrv12
    port map (
            O => \N__9557\,
            I => \CUMBEn_c\
        );

    \I__2077\ : IoInMux
    port map (
            O => \N__9554\,
            I => \N__9551\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__9551\,
            I => \N__9548\
        );

    \I__2075\ : Span4Mux_s1_v
    port map (
            O => \N__9548\,
            I => \N__9544\
        );

    \I__2074\ : InMux
    port map (
            O => \N__9547\,
            I => \N__9541\
        );

    \I__2073\ : Span4Mux_v
    port map (
            O => \N__9544\,
            I => \N__9538\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__9541\,
            I => \N__9535\
        );

    \I__2071\ : Span4Mux_v
    port map (
            O => \N__9538\,
            I => \N__9532\
        );

    \I__2070\ : Span4Mux_v
    port map (
            O => \N__9535\,
            I => \N__9529\
        );

    \I__2069\ : Odrv4
    port map (
            O => \N__9532\,
            I => \LMBEn_c\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__9529\,
            I => \LMBEn_c\
        );

    \I__2067\ : IoInMux
    port map (
            O => \N__9524\,
            I => \N__9521\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__9521\,
            I => \N__9518\
        );

    \I__2065\ : Span4Mux_s2_h
    port map (
            O => \N__9518\,
            I => \N__9515\
        );

    \I__2064\ : Sp12to4
    port map (
            O => \N__9515\,
            I => \N__9512\
        );

    \I__2063\ : Span12Mux_s10_v
    port map (
            O => \N__9512\,
            I => \N__9509\
        );

    \I__2062\ : Span12Mux_h
    port map (
            O => \N__9509\,
            I => \N__9506\
        );

    \I__2061\ : Odrv12
    port map (
            O => \N__9506\,
            I => \CLMBEn_c\
        );

    \I__2060\ : IoInMux
    port map (
            O => \N__9503\,
            I => \N__9500\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__9500\,
            I => \N__9497\
        );

    \I__2058\ : Span4Mux_s2_h
    port map (
            O => \N__9497\,
            I => \N__9494\
        );

    \I__2057\ : Sp12to4
    port map (
            O => \N__9494\,
            I => \N__9491\
        );

    \I__2056\ : Span12Mux_v
    port map (
            O => \N__9491\,
            I => \N__9488\
        );

    \I__2055\ : Odrv12
    port map (
            O => \N__9488\,
            I => \CUUBEn_c\
        );

    \I__2054\ : IoInMux
    port map (
            O => \N__9485\,
            I => \N__9482\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__9482\,
            I => \N__9479\
        );

    \I__2052\ : Span12Mux_s7_v
    port map (
            O => \N__9479\,
            I => \N__9476\
        );

    \I__2051\ : Span12Mux_h
    port map (
            O => \N__9476\,
            I => \N__9473\
        );

    \I__2050\ : Odrv12
    port map (
            O => \N__9473\,
            I => \ASn_c\
        );

    \I__2049\ : CEMux
    port map (
            O => \N__9470\,
            I => \N__9467\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__9467\,
            I => \N__9464\
        );

    \I__2047\ : Span4Mux_v
    port map (
            O => \N__9464\,
            I => \N__9461\
        );

    \I__2046\ : Odrv4
    port map (
            O => \N__9461\,
            I => \U712_REG_SM.N_99_0_0\
        );

    \I__2045\ : CascadeMux
    port map (
            O => \N__9458\,
            I => \N__9454\
        );

    \I__2044\ : InMux
    port map (
            O => \N__9457\,
            I => \N__9447\
        );

    \I__2043\ : InMux
    port map (
            O => \N__9454\,
            I => \N__9444\
        );

    \I__2042\ : InMux
    port map (
            O => \N__9453\,
            I => \N__9441\
        );

    \I__2041\ : InMux
    port map (
            O => \N__9452\,
            I => \N__9436\
        );

    \I__2040\ : InMux
    port map (
            O => \N__9451\,
            I => \N__9432\
        );

    \I__2039\ : CascadeMux
    port map (
            O => \N__9450\,
            I => \N__9427\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__9447\,
            I => \N__9422\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__9444\,
            I => \N__9419\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__9441\,
            I => \N__9416\
        );

    \I__2035\ : InMux
    port map (
            O => \N__9440\,
            I => \N__9411\
        );

    \I__2034\ : CascadeMux
    port map (
            O => \N__9439\,
            I => \N__9408\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__9436\,
            I => \N__9405\
        );

    \I__2032\ : InMux
    port map (
            O => \N__9435\,
            I => \N__9402\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__9432\,
            I => \N__9399\
        );

    \I__2030\ : InMux
    port map (
            O => \N__9431\,
            I => \N__9396\
        );

    \I__2029\ : InMux
    port map (
            O => \N__9430\,
            I => \N__9389\
        );

    \I__2028\ : InMux
    port map (
            O => \N__9427\,
            I => \N__9389\
        );

    \I__2027\ : InMux
    port map (
            O => \N__9426\,
            I => \N__9389\
        );

    \I__2026\ : InMux
    port map (
            O => \N__9425\,
            I => \N__9386\
        );

    \I__2025\ : Span4Mux_h
    port map (
            O => \N__9422\,
            I => \N__9381\
        );

    \I__2024\ : Span4Mux_v
    port map (
            O => \N__9419\,
            I => \N__9381\
        );

    \I__2023\ : Span4Mux_v
    port map (
            O => \N__9416\,
            I => \N__9378\
        );

    \I__2022\ : InMux
    port map (
            O => \N__9415\,
            I => \N__9373\
        );

    \I__2021\ : InMux
    port map (
            O => \N__9414\,
            I => \N__9373\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__9411\,
            I => \N__9370\
        );

    \I__2019\ : InMux
    port map (
            O => \N__9408\,
            I => \N__9367\
        );

    \I__2018\ : Span4Mux_h
    port map (
            O => \N__9405\,
            I => \N__9362\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__9402\,
            I => \N__9362\
        );

    \I__2016\ : Odrv12
    port map (
            O => \N__9399\,
            I => \U712_REG_SM_C1_SYNC_1\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__9396\,
            I => \U712_REG_SM_C1_SYNC_1\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__9389\,
            I => \U712_REG_SM_C1_SYNC_1\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__9386\,
            I => \U712_REG_SM_C1_SYNC_1\
        );

    \I__2012\ : Odrv4
    port map (
            O => \N__9381\,
            I => \U712_REG_SM_C1_SYNC_1\
        );

    \I__2011\ : Odrv4
    port map (
            O => \N__9378\,
            I => \U712_REG_SM_C1_SYNC_1\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__9373\,
            I => \U712_REG_SM_C1_SYNC_1\
        );

    \I__2009\ : Odrv4
    port map (
            O => \N__9370\,
            I => \U712_REG_SM_C1_SYNC_1\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__9367\,
            I => \U712_REG_SM_C1_SYNC_1\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__9362\,
            I => \U712_REG_SM_C1_SYNC_1\
        );

    \I__2006\ : InMux
    port map (
            O => \N__9341\,
            I => \N__9338\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__9338\,
            I => \U712_REG_SM_LDSn_6_0\
        );

    \I__2004\ : InMux
    port map (
            O => \N__9335\,
            I => \N__9332\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__9332\,
            I => \U712_CHIP_RAM.m185_1\
        );

    \I__2002\ : IoInMux
    port map (
            O => \N__9329\,
            I => \N__9326\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__9326\,
            I => \N__9323\
        );

    \I__2000\ : Span4Mux_s3_h
    port map (
            O => \N__9323\,
            I => \N__9320\
        );

    \I__1999\ : Span4Mux_v
    port map (
            O => \N__9320\,
            I => \N__9317\
        );

    \I__1998\ : Sp12to4
    port map (
            O => \N__9317\,
            I => \N__9314\
        );

    \I__1997\ : Span12Mux_h
    port map (
            O => \N__9314\,
            I => \N__9311\
        );

    \I__1996\ : Odrv12
    port map (
            O => \N__9311\,
            I => \CMA_c_5\
        );

    \I__1995\ : InMux
    port map (
            O => \N__9308\,
            I => \N__9305\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__9305\,
            I => \N__9302\
        );

    \I__1993\ : Span4Mux_h
    port map (
            O => \N__9302\,
            I => \N__9299\
        );

    \I__1992\ : Odrv4
    port map (
            O => \N__9299\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__1991\ : InMux
    port map (
            O => \N__9296\,
            I => \N__9293\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__9293\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__1989\ : InMux
    port map (
            O => \N__9290\,
            I => \N__9287\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__9287\,
            I => \N__9284\
        );

    \I__1987\ : Span4Mux_v
    port map (
            O => \N__9284\,
            I => \N__9281\
        );

    \I__1986\ : Span4Mux_v
    port map (
            O => \N__9281\,
            I => \N__9278\
        );

    \I__1985\ : Sp12to4
    port map (
            O => \N__9278\,
            I => \N__9275\
        );

    \I__1984\ : Span12Mux_h
    port map (
            O => \N__9275\,
            I => \N__9272\
        );

    \I__1983\ : Odrv12
    port map (
            O => \N__9272\,
            I => \A_c_19\
        );

    \I__1982\ : InMux
    port map (
            O => \N__9269\,
            I => \N__9266\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__9266\,
            I => \U712_CHIP_RAM.m194_0\
        );

    \I__1980\ : IoInMux
    port map (
            O => \N__9263\,
            I => \N__9260\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__9260\,
            I => \N__9257\
        );

    \I__1978\ : Span4Mux_s3_h
    port map (
            O => \N__9257\,
            I => \N__9254\
        );

    \I__1977\ : Span4Mux_v
    port map (
            O => \N__9254\,
            I => \N__9251\
        );

    \I__1976\ : Sp12to4
    port map (
            O => \N__9251\,
            I => \N__9248\
        );

    \I__1975\ : Span12Mux_h
    port map (
            O => \N__9248\,
            I => \N__9245\
        );

    \I__1974\ : Odrv12
    port map (
            O => \N__9245\,
            I => \CMA_c_9\
        );

    \I__1973\ : InMux
    port map (
            O => \N__9242\,
            I => \N__9238\
        );

    \I__1972\ : InMux
    port map (
            O => \N__9241\,
            I => \N__9235\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__9238\,
            I => \N__9229\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__9235\,
            I => \N__9225\
        );

    \I__1969\ : InMux
    port map (
            O => \N__9234\,
            I => \N__9222\
        );

    \I__1968\ : InMux
    port map (
            O => \N__9233\,
            I => \N__9217\
        );

    \I__1967\ : InMux
    port map (
            O => \N__9232\,
            I => \N__9214\
        );

    \I__1966\ : Span4Mux_h
    port map (
            O => \N__9229\,
            I => \N__9211\
        );

    \I__1965\ : InMux
    port map (
            O => \N__9228\,
            I => \N__9208\
        );

    \I__1964\ : Span12Mux_v
    port map (
            O => \N__9225\,
            I => \N__9205\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__9222\,
            I => \N__9202\
        );

    \I__1962\ : InMux
    port map (
            O => \N__9221\,
            I => \N__9199\
        );

    \I__1961\ : InMux
    port map (
            O => \N__9220\,
            I => \N__9196\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__9217\,
            I => \N__9187\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__9214\,
            I => \N__9187\
        );

    \I__1958\ : Span4Mux_v
    port map (
            O => \N__9211\,
            I => \N__9187\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__9208\,
            I => \N__9187\
        );

    \I__1956\ : Odrv12
    port map (
            O => \N__9205\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1955\ : Odrv4
    port map (
            O => \N__9202\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__9199\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__9196\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1952\ : Odrv4
    port map (
            O => \N__9187\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1951\ : InMux
    port map (
            O => \N__9176\,
            I => \N__9173\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__9173\,
            I => \N__9170\
        );

    \I__1949\ : Odrv4
    port map (
            O => \N__9170\,
            I => \U712_CHIP_RAM.d_N_7_0\
        );

    \I__1948\ : InMux
    port map (
            O => \N__9167\,
            I => \N__9164\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__9164\,
            I => \N__9161\
        );

    \I__1946\ : Span4Mux_v
    port map (
            O => \N__9161\,
            I => \N__9158\
        );

    \I__1945\ : Sp12to4
    port map (
            O => \N__9158\,
            I => \N__9155\
        );

    \I__1944\ : Span12Mux_v
    port map (
            O => \N__9155\,
            I => \N__9152\
        );

    \I__1943\ : Span12Mux_h
    port map (
            O => \N__9152\,
            I => \N__9149\
        );

    \I__1942\ : Odrv12
    port map (
            O => \N__9149\,
            I => \A_c_18\
        );

    \I__1941\ : InMux
    port map (
            O => \N__9146\,
            I => \N__9142\
        );

    \I__1940\ : InMux
    port map (
            O => \N__9145\,
            I => \N__9139\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__9142\,
            I => \N__9136\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__9139\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\
        );

    \I__1937\ : Odrv4
    port map (
            O => \N__9136\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\
        );

    \I__1936\ : CascadeMux
    port map (
            O => \N__9131\,
            I => \N__9127\
        );

    \I__1935\ : InMux
    port map (
            O => \N__9130\,
            I => \N__9115\
        );

    \I__1934\ : InMux
    port map (
            O => \N__9127\,
            I => \N__9112\
        );

    \I__1933\ : InMux
    port map (
            O => \N__9126\,
            I => \N__9107\
        );

    \I__1932\ : InMux
    port map (
            O => \N__9125\,
            I => \N__9107\
        );

    \I__1931\ : InMux
    port map (
            O => \N__9124\,
            I => \N__9104\
        );

    \I__1930\ : InMux
    port map (
            O => \N__9123\,
            I => \N__9099\
        );

    \I__1929\ : InMux
    port map (
            O => \N__9122\,
            I => \N__9096\
        );

    \I__1928\ : CascadeMux
    port map (
            O => \N__9121\,
            I => \N__9093\
        );

    \I__1927\ : CascadeMux
    port map (
            O => \N__9120\,
            I => \N__9090\
        );

    \I__1926\ : InMux
    port map (
            O => \N__9119\,
            I => \N__9081\
        );

    \I__1925\ : InMux
    port map (
            O => \N__9118\,
            I => \N__9081\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__9115\,
            I => \N__9078\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__9112\,
            I => \N__9071\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__9107\,
            I => \N__9071\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__9104\,
            I => \N__9071\
        );

    \I__1920\ : InMux
    port map (
            O => \N__9103\,
            I => \N__9068\
        );

    \I__1919\ : InMux
    port map (
            O => \N__9102\,
            I => \N__9065\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__9099\,
            I => \N__9062\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__9096\,
            I => \N__9059\
        );

    \I__1916\ : InMux
    port map (
            O => \N__9093\,
            I => \N__9056\
        );

    \I__1915\ : InMux
    port map (
            O => \N__9090\,
            I => \N__9049\
        );

    \I__1914\ : InMux
    port map (
            O => \N__9089\,
            I => \N__9049\
        );

    \I__1913\ : InMux
    port map (
            O => \N__9088\,
            I => \N__9049\
        );

    \I__1912\ : InMux
    port map (
            O => \N__9087\,
            I => \N__9044\
        );

    \I__1911\ : InMux
    port map (
            O => \N__9086\,
            I => \N__9044\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__9081\,
            I => \N__9037\
        );

    \I__1909\ : Span4Mux_h
    port map (
            O => \N__9078\,
            I => \N__9037\
        );

    \I__1908\ : Span4Mux_h
    port map (
            O => \N__9071\,
            I => \N__9037\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__9068\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__9065\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1905\ : Odrv4
    port map (
            O => \N__9062\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1904\ : Odrv4
    port map (
            O => \N__9059\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__9056\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__9049\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__9044\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1900\ : Odrv4
    port map (
            O => \N__9037\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1899\ : InMux
    port map (
            O => \N__9020\,
            I => \N__9017\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__9017\,
            I => \U712_CHIP_RAM.N_204\
        );

    \I__1897\ : InMux
    port map (
            O => \N__9014\,
            I => \N__9011\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__9011\,
            I => \N__9008\
        );

    \I__1895\ : Span4Mux_h
    port map (
            O => \N__9008\,
            I => \N__9005\
        );

    \I__1894\ : Sp12to4
    port map (
            O => \N__9005\,
            I => \N__9002\
        );

    \I__1893\ : Span12Mux_v
    port map (
            O => \N__9002\,
            I => \N__8999\
        );

    \I__1892\ : Span12Mux_h
    port map (
            O => \N__8999\,
            I => \N__8996\
        );

    \I__1891\ : Odrv12
    port map (
            O => \N__8996\,
            I => \A_c_3\
        );

    \I__1890\ : InMux
    port map (
            O => \N__8993\,
            I => \N__8989\
        );

    \I__1889\ : InMux
    port map (
            O => \N__8992\,
            I => \N__8986\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__8989\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__8986\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\
        );

    \I__1886\ : InMux
    port map (
            O => \N__8981\,
            I => \N__8967\
        );

    \I__1885\ : InMux
    port map (
            O => \N__8980\,
            I => \N__8967\
        );

    \I__1884\ : InMux
    port map (
            O => \N__8979\,
            I => \N__8967\
        );

    \I__1883\ : InMux
    port map (
            O => \N__8978\,
            I => \N__8962\
        );

    \I__1882\ : InMux
    port map (
            O => \N__8977\,
            I => \N__8962\
        );

    \I__1881\ : InMux
    port map (
            O => \N__8976\,
            I => \N__8955\
        );

    \I__1880\ : InMux
    port map (
            O => \N__8975\,
            I => \N__8955\
        );

    \I__1879\ : InMux
    port map (
            O => \N__8974\,
            I => \N__8955\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__8967\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__8962\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__8955\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\
        );

    \I__1875\ : InMux
    port map (
            O => \N__8948\,
            I => \N__8945\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__8945\,
            I => \N__8942\
        );

    \I__1873\ : Span12Mux_h
    port map (
            O => \N__8942\,
            I => \N__8939\
        );

    \I__1872\ : Odrv12
    port map (
            O => \N__8939\,
            I => \A_c_8\
        );

    \I__1871\ : InMux
    port map (
            O => \N__8936\,
            I => \N__8932\
        );

    \I__1870\ : InMux
    port map (
            O => \N__8935\,
            I => \N__8929\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__8932\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__8929\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\
        );

    \I__1867\ : InMux
    port map (
            O => \N__8924\,
            I => \N__8916\
        );

    \I__1866\ : InMux
    port map (
            O => \N__8923\,
            I => \N__8910\
        );

    \I__1865\ : InMux
    port map (
            O => \N__8922\,
            I => \N__8907\
        );

    \I__1864\ : InMux
    port map (
            O => \N__8921\,
            I => \N__8900\
        );

    \I__1863\ : InMux
    port map (
            O => \N__8920\,
            I => \N__8900\
        );

    \I__1862\ : InMux
    port map (
            O => \N__8919\,
            I => \N__8900\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__8916\,
            I => \N__8896\
        );

    \I__1860\ : InMux
    port map (
            O => \N__8915\,
            I => \N__8889\
        );

    \I__1859\ : InMux
    port map (
            O => \N__8914\,
            I => \N__8889\
        );

    \I__1858\ : InMux
    port map (
            O => \N__8913\,
            I => \N__8889\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__8910\,
            I => \N__8875\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__8907\,
            I => \N__8875\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__8900\,
            I => \N__8875\
        );

    \I__1854\ : CascadeMux
    port map (
            O => \N__8899\,
            I => \N__8868\
        );

    \I__1853\ : Span4Mux_v
    port map (
            O => \N__8896\,
            I => \N__8861\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__8889\,
            I => \N__8861\
        );

    \I__1851\ : InMux
    port map (
            O => \N__8888\,
            I => \N__8854\
        );

    \I__1850\ : InMux
    port map (
            O => \N__8887\,
            I => \N__8854\
        );

    \I__1849\ : InMux
    port map (
            O => \N__8886\,
            I => \N__8854\
        );

    \I__1848\ : InMux
    port map (
            O => \N__8885\,
            I => \N__8847\
        );

    \I__1847\ : InMux
    port map (
            O => \N__8884\,
            I => \N__8847\
        );

    \I__1846\ : InMux
    port map (
            O => \N__8883\,
            I => \N__8847\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__8882\,
            I => \N__8842\
        );

    \I__1844\ : Span4Mux_v
    port map (
            O => \N__8875\,
            I => \N__8838\
        );

    \I__1843\ : InMux
    port map (
            O => \N__8874\,
            I => \N__8833\
        );

    \I__1842\ : InMux
    port map (
            O => \N__8873\,
            I => \N__8833\
        );

    \I__1841\ : InMux
    port map (
            O => \N__8872\,
            I => \N__8830\
        );

    \I__1840\ : InMux
    port map (
            O => \N__8871\,
            I => \N__8821\
        );

    \I__1839\ : InMux
    port map (
            O => \N__8868\,
            I => \N__8821\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8867\,
            I => \N__8821\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8866\,
            I => \N__8821\
        );

    \I__1836\ : Span4Mux_h
    port map (
            O => \N__8861\,
            I => \N__8816\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__8854\,
            I => \N__8816\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__8847\,
            I => \N__8813\
        );

    \I__1833\ : InMux
    port map (
            O => \N__8846\,
            I => \N__8808\
        );

    \I__1832\ : InMux
    port map (
            O => \N__8845\,
            I => \N__8808\
        );

    \I__1831\ : InMux
    port map (
            O => \N__8842\,
            I => \N__8803\
        );

    \I__1830\ : InMux
    port map (
            O => \N__8841\,
            I => \N__8803\
        );

    \I__1829\ : Odrv4
    port map (
            O => \N__8838\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__8833\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8830\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__8821\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1825\ : Odrv4
    port map (
            O => \N__8816\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1824\ : Odrv4
    port map (
            O => \N__8813\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__8808\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__8803\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1821\ : InMux
    port map (
            O => \N__8786\,
            I => \N__8781\
        );

    \I__1820\ : InMux
    port map (
            O => \N__8785\,
            I => \N__8776\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__8784\,
            I => \N__8773\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__8781\,
            I => \N__8768\
        );

    \I__1817\ : InMux
    port map (
            O => \N__8780\,
            I => \N__8763\
        );

    \I__1816\ : InMux
    port map (
            O => \N__8779\,
            I => \N__8763\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__8776\,
            I => \N__8760\
        );

    \I__1814\ : InMux
    port map (
            O => \N__8773\,
            I => \N__8757\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8772\,
            I => \N__8754\
        );

    \I__1812\ : InMux
    port map (
            O => \N__8771\,
            I => \N__8751\
        );

    \I__1811\ : Odrv4
    port map (
            O => \N__8768\,
            I => \U712_CHIP_RAM.N_31_0\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__8763\,
            I => \U712_CHIP_RAM.N_31_0\
        );

    \I__1809\ : Odrv4
    port map (
            O => \N__8760\,
            I => \U712_CHIP_RAM.N_31_0\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__8757\,
            I => \U712_CHIP_RAM.N_31_0\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__8754\,
            I => \U712_CHIP_RAM.N_31_0\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__8751\,
            I => \U712_CHIP_RAM.N_31_0\
        );

    \I__1805\ : CascadeMux
    port map (
            O => \N__8738\,
            I => \N__8735\
        );

    \I__1804\ : InMux
    port map (
            O => \N__8735\,
            I => \N__8732\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__8732\,
            I => \U712_CHIP_RAM.DBENn_8_0\
        );

    \I__1802\ : IoInMux
    port map (
            O => \N__8729\,
            I => \N__8726\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__8726\,
            I => \N__8723\
        );

    \I__1800\ : IoSpan4Mux
    port map (
            O => \N__8723\,
            I => \N__8720\
        );

    \I__1799\ : Sp12to4
    port map (
            O => \N__8720\,
            I => \N__8716\
        );

    \I__1798\ : InMux
    port map (
            O => \N__8719\,
            I => \N__8713\
        );

    \I__1797\ : Span12Mux_s7_v
    port map (
            O => \N__8716\,
            I => \N__8710\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__8713\,
            I => \N__8707\
        );

    \I__1795\ : Odrv12
    port map (
            O => \N__8710\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1794\ : Odrv4
    port map (
            O => \N__8707\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1793\ : CascadeMux
    port map (
            O => \N__8702\,
            I => \N__8699\
        );

    \I__1792\ : InMux
    port map (
            O => \N__8699\,
            I => \N__8696\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__8696\,
            I => \N__8693\
        );

    \I__1790\ : Span4Mux_h
    port map (
            O => \N__8693\,
            I => \N__8690\
        );

    \I__1789\ : Odrv4
    port map (
            O => \N__8690\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__1788\ : CascadeMux
    port map (
            O => \N__8687\,
            I => \N__8682\
        );

    \I__1787\ : CascadeMux
    port map (
            O => \N__8686\,
            I => \N__8677\
        );

    \I__1786\ : CascadeMux
    port map (
            O => \N__8685\,
            I => \N__8673\
        );

    \I__1785\ : InMux
    port map (
            O => \N__8682\,
            I => \N__8659\
        );

    \I__1784\ : InMux
    port map (
            O => \N__8681\,
            I => \N__8659\
        );

    \I__1783\ : CascadeMux
    port map (
            O => \N__8680\,
            I => \N__8655\
        );

    \I__1782\ : InMux
    port map (
            O => \N__8677\,
            I => \N__8650\
        );

    \I__1781\ : InMux
    port map (
            O => \N__8676\,
            I => \N__8647\
        );

    \I__1780\ : InMux
    port map (
            O => \N__8673\,
            I => \N__8642\
        );

    \I__1779\ : InMux
    port map (
            O => \N__8672\,
            I => \N__8642\
        );

    \I__1778\ : InMux
    port map (
            O => \N__8671\,
            I => \N__8636\
        );

    \I__1777\ : InMux
    port map (
            O => \N__8670\,
            I => \N__8629\
        );

    \I__1776\ : InMux
    port map (
            O => \N__8669\,
            I => \N__8629\
        );

    \I__1775\ : InMux
    port map (
            O => \N__8668\,
            I => \N__8629\
        );

    \I__1774\ : InMux
    port map (
            O => \N__8667\,
            I => \N__8618\
        );

    \I__1773\ : InMux
    port map (
            O => \N__8666\,
            I => \N__8618\
        );

    \I__1772\ : InMux
    port map (
            O => \N__8665\,
            I => \N__8618\
        );

    \I__1771\ : InMux
    port map (
            O => \N__8664\,
            I => \N__8615\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__8659\,
            I => \N__8612\
        );

    \I__1769\ : InMux
    port map (
            O => \N__8658\,
            I => \N__8603\
        );

    \I__1768\ : InMux
    port map (
            O => \N__8655\,
            I => \N__8603\
        );

    \I__1767\ : InMux
    port map (
            O => \N__8654\,
            I => \N__8603\
        );

    \I__1766\ : InMux
    port map (
            O => \N__8653\,
            I => \N__8603\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__8650\,
            I => \N__8596\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8647\,
            I => \N__8596\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__8642\,
            I => \N__8596\
        );

    \I__1762\ : CascadeMux
    port map (
            O => \N__8641\,
            I => \N__8590\
        );

    \I__1761\ : InMux
    port map (
            O => \N__8640\,
            I => \N__8586\
        );

    \I__1760\ : InMux
    port map (
            O => \N__8639\,
            I => \N__8582\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__8636\,
            I => \N__8577\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__8629\,
            I => \N__8577\
        );

    \I__1757\ : InMux
    port map (
            O => \N__8628\,
            I => \N__8570\
        );

    \I__1756\ : InMux
    port map (
            O => \N__8627\,
            I => \N__8570\
        );

    \I__1755\ : InMux
    port map (
            O => \N__8626\,
            I => \N__8570\
        );

    \I__1754\ : InMux
    port map (
            O => \N__8625\,
            I => \N__8567\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__8618\,
            I => \N__8564\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__8615\,
            I => \N__8555\
        );

    \I__1751\ : Span4Mux_v
    port map (
            O => \N__8612\,
            I => \N__8555\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__8603\,
            I => \N__8555\
        );

    \I__1749\ : Span4Mux_v
    port map (
            O => \N__8596\,
            I => \N__8555\
        );

    \I__1748\ : InMux
    port map (
            O => \N__8595\,
            I => \N__8548\
        );

    \I__1747\ : InMux
    port map (
            O => \N__8594\,
            I => \N__8548\
        );

    \I__1746\ : InMux
    port map (
            O => \N__8593\,
            I => \N__8548\
        );

    \I__1745\ : InMux
    port map (
            O => \N__8590\,
            I => \N__8545\
        );

    \I__1744\ : InMux
    port map (
            O => \N__8589\,
            I => \N__8542\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__8586\,
            I => \N__8539\
        );

    \I__1742\ : InMux
    port map (
            O => \N__8585\,
            I => \N__8536\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__8582\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1740\ : Odrv4
    port map (
            O => \N__8577\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__8570\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__8567\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1737\ : Odrv4
    port map (
            O => \N__8564\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1736\ : Odrv4
    port map (
            O => \N__8555\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__8548\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__8545\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__8542\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1732\ : Odrv12
    port map (
            O => \N__8539\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__8536\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1730\ : InMux
    port map (
            O => \N__8513\,
            I => \N__8510\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__8510\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0\
        );

    \I__1728\ : IoInMux
    port map (
            O => \N__8507\,
            I => \N__8504\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__8504\,
            I => \N__8501\
        );

    \I__1726\ : Span12Mux_s1_v
    port map (
            O => \N__8501\,
            I => \N__8498\
        );

    \I__1725\ : Span12Mux_v
    port map (
            O => \N__8498\,
            I => \N__8494\
        );

    \I__1724\ : InMux
    port map (
            O => \N__8497\,
            I => \N__8491\
        );

    \I__1723\ : Odrv12
    port map (
            O => \N__8494\,
            I => \LATCH_CLK_c\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__8491\,
            I => \LATCH_CLK_c\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__8486\,
            I => \U712_CHIP_RAM.m191_0_cascade_\
        );

    \I__1720\ : InMux
    port map (
            O => \N__8483\,
            I => \N__8480\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__8480\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__1718\ : InMux
    port map (
            O => \N__8477\,
            I => \N__8474\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__8474\,
            I => \U712_CHIP_RAM.d_N_6_4\
        );

    \I__1716\ : IoInMux
    port map (
            O => \N__8471\,
            I => \N__8468\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__8468\,
            I => \N__8465\
        );

    \I__1714\ : Span4Mux_s0_v
    port map (
            O => \N__8465\,
            I => \N__8462\
        );

    \I__1713\ : Span4Mux_v
    port map (
            O => \N__8462\,
            I => \N__8458\
        );

    \I__1712\ : InMux
    port map (
            O => \N__8461\,
            I => \N__8455\
        );

    \I__1711\ : Span4Mux_v
    port map (
            O => \N__8458\,
            I => \N__8452\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__8455\,
            I => \N__8449\
        );

    \I__1709\ : Sp12to4
    port map (
            O => \N__8452\,
            I => \N__8446\
        );

    \I__1708\ : Span4Mux_v
    port map (
            O => \N__8449\,
            I => \N__8443\
        );

    \I__1707\ : Span12Mux_h
    port map (
            O => \N__8446\,
            I => \N__8440\
        );

    \I__1706\ : Sp12to4
    port map (
            O => \N__8443\,
            I => \N__8437\
        );

    \I__1705\ : Span12Mux_v
    port map (
            O => \N__8440\,
            I => \N__8432\
        );

    \I__1704\ : Span12Mux_h
    port map (
            O => \N__8437\,
            I => \N__8432\
        );

    \I__1703\ : Odrv12
    port map (
            O => \N__8432\,
            I => \A_c_10\
        );

    \I__1702\ : CascadeMux
    port map (
            O => \N__8429\,
            I => \N__8426\
        );

    \I__1701\ : InMux
    port map (
            O => \N__8426\,
            I => \N__8422\
        );

    \I__1700\ : InMux
    port map (
            O => \N__8425\,
            I => \N__8419\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__8422\,
            I => \N__8416\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__8419\,
            I => \N__8413\
        );

    \I__1697\ : Span4Mux_h
    port map (
            O => \N__8416\,
            I => \N__8410\
        );

    \I__1696\ : Span4Mux_v
    port map (
            O => \N__8413\,
            I => \N__8405\
        );

    \I__1695\ : Span4Mux_v
    port map (
            O => \N__8410\,
            I => \N__8405\
        );

    \I__1694\ : Odrv4
    port map (
            O => \N__8405\,
            I => \U712_CHIP_RAM.m184_m2_0_a2_0\
        );

    \I__1693\ : CascadeMux
    port map (
            O => \N__8402\,
            I => \U712_CHIP_RAM.m184_0_cascade_\
        );

    \I__1692\ : InMux
    port map (
            O => \N__8399\,
            I => \N__8396\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__8396\,
            I => \U712_CHIP_RAM.m184_1\
        );

    \I__1690\ : InMux
    port map (
            O => \N__8393\,
            I => \N__8390\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__8390\,
            I => \N__8387\
        );

    \I__1688\ : Span4Mux_v
    port map (
            O => \N__8387\,
            I => \N__8384\
        );

    \I__1687\ : Span4Mux_v
    port map (
            O => \N__8384\,
            I => \N__8381\
        );

    \I__1686\ : Sp12to4
    port map (
            O => \N__8381\,
            I => \N__8378\
        );

    \I__1685\ : Span12Mux_h
    port map (
            O => \N__8378\,
            I => \N__8375\
        );

    \I__1684\ : Odrv12
    port map (
            O => \N__8375\,
            I => \A_c_15\
        );

    \I__1683\ : InMux
    port map (
            O => \N__8372\,
            I => \N__8365\
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__8371\,
            I => \N__8362\
        );

    \I__1681\ : InMux
    port map (
            O => \N__8370\,
            I => \N__8357\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__8369\,
            I => \N__8351\
        );

    \I__1679\ : InMux
    port map (
            O => \N__8368\,
            I => \N__8348\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__8365\,
            I => \N__8345\
        );

    \I__1677\ : InMux
    port map (
            O => \N__8362\,
            I => \N__8338\
        );

    \I__1676\ : InMux
    port map (
            O => \N__8361\,
            I => \N__8338\
        );

    \I__1675\ : InMux
    port map (
            O => \N__8360\,
            I => \N__8338\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__8357\,
            I => \N__8335\
        );

    \I__1673\ : InMux
    port map (
            O => \N__8356\,
            I => \N__8330\
        );

    \I__1672\ : InMux
    port map (
            O => \N__8355\,
            I => \N__8330\
        );

    \I__1671\ : InMux
    port map (
            O => \N__8354\,
            I => \N__8325\
        );

    \I__1670\ : InMux
    port map (
            O => \N__8351\,
            I => \N__8325\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__8348\,
            I => \N__8322\
        );

    \I__1668\ : Span4Mux_h
    port map (
            O => \N__8345\,
            I => \N__8317\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__8338\,
            I => \N__8317\
        );

    \I__1666\ : Odrv12
    port map (
            O => \N__8335\,
            I => \U712_CHIP_RAM.N_3_0\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__8330\,
            I => \U712_CHIP_RAM.N_3_0\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__8325\,
            I => \U712_CHIP_RAM.N_3_0\
        );

    \I__1663\ : Odrv4
    port map (
            O => \N__8322\,
            I => \U712_CHIP_RAM.N_3_0\
        );

    \I__1662\ : Odrv4
    port map (
            O => \N__8317\,
            I => \U712_CHIP_RAM.N_3_0\
        );

    \I__1661\ : CascadeMux
    port map (
            O => \N__8306\,
            I => \N__8300\
        );

    \I__1660\ : InMux
    port map (
            O => \N__8305\,
            I => \N__8296\
        );

    \I__1659\ : CascadeMux
    port map (
            O => \N__8304\,
            I => \N__8291\
        );

    \I__1658\ : InMux
    port map (
            O => \N__8303\,
            I => \N__8286\
        );

    \I__1657\ : InMux
    port map (
            O => \N__8300\,
            I => \N__8286\
        );

    \I__1656\ : InMux
    port map (
            O => \N__8299\,
            I => \N__8283\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__8296\,
            I => \N__8280\
        );

    \I__1654\ : InMux
    port map (
            O => \N__8295\,
            I => \N__8275\
        );

    \I__1653\ : InMux
    port map (
            O => \N__8294\,
            I => \N__8275\
        );

    \I__1652\ : InMux
    port map (
            O => \N__8291\,
            I => \N__8272\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__8286\,
            I => \N__8269\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__8283\,
            I => \N__8266\
        );

    \I__1649\ : Span4Mux_h
    port map (
            O => \N__8280\,
            I => \N__8263\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__8275\,
            I => \U712_CHIP_RAM.m186_m2_0_a2_0\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__8272\,
            I => \U712_CHIP_RAM.m186_m2_0_a2_0\
        );

    \I__1646\ : Odrv4
    port map (
            O => \N__8269\,
            I => \U712_CHIP_RAM.m186_m2_0_a2_0\
        );

    \I__1645\ : Odrv4
    port map (
            O => \N__8266\,
            I => \U712_CHIP_RAM.m186_m2_0_a2_0\
        );

    \I__1644\ : Odrv4
    port map (
            O => \N__8263\,
            I => \U712_CHIP_RAM.m186_m2_0_a2_0\
        );

    \I__1643\ : CascadeMux
    port map (
            O => \N__8252\,
            I => \U712_CHIP_RAM.m190_0_cascade_\
        );

    \I__1642\ : InMux
    port map (
            O => \N__8249\,
            I => \N__8246\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__8246\,
            I => \U712_CHIP_RAM.m190_1\
        );

    \I__1640\ : IoInMux
    port map (
            O => \N__8243\,
            I => \N__8240\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__8240\,
            I => \N__8237\
        );

    \I__1638\ : Span4Mux_s0_h
    port map (
            O => \N__8237\,
            I => \N__8234\
        );

    \I__1637\ : Sp12to4
    port map (
            O => \N__8234\,
            I => \N__8231\
        );

    \I__1636\ : Span12Mux_v
    port map (
            O => \N__8231\,
            I => \N__8228\
        );

    \I__1635\ : Span12Mux_h
    port map (
            O => \N__8228\,
            I => \N__8225\
        );

    \I__1634\ : Odrv12
    port map (
            O => \N__8225\,
            I => \CMA_c_6\
        );

    \I__1633\ : InMux
    port map (
            O => \N__8222\,
            I => \N__8219\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__8219\,
            I => \N__8216\
        );

    \I__1631\ : Odrv4
    port map (
            O => \N__8216\,
            I => \U712_CHIP_RAM.d_N_6_3\
        );

    \I__1630\ : CascadeMux
    port map (
            O => \N__8213\,
            I => \U712_CHIP_RAM.N_208_cascade_\
        );

    \I__1629\ : InMux
    port map (
            O => \N__8210\,
            I => \N__8206\
        );

    \I__1628\ : InMux
    port map (
            O => \N__8209\,
            I => \N__8203\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__8206\,
            I => \N__8199\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__8203\,
            I => \N__8196\
        );

    \I__1625\ : InMux
    port map (
            O => \N__8202\,
            I => \N__8193\
        );

    \I__1624\ : Span4Mux_h
    port map (
            O => \N__8199\,
            I => \N__8190\
        );

    \I__1623\ : Span4Mux_v
    port map (
            O => \N__8196\,
            I => \N__8187\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__8193\,
            I => \N__8184\
        );

    \I__1621\ : Odrv4
    port map (
            O => \N__8190\,
            I => \N_99_0\
        );

    \I__1620\ : Odrv4
    port map (
            O => \N__8187\,
            I => \N_99_0\
        );

    \I__1619\ : Odrv12
    port map (
            O => \N__8184\,
            I => \N_99_0\
        );

    \I__1618\ : IoInMux
    port map (
            O => \N__8177\,
            I => \N__8174\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__8174\,
            I => \N__8171\
        );

    \I__1616\ : Span12Mux_s5_v
    port map (
            O => \N__8171\,
            I => \N__8168\
        );

    \I__1615\ : Span12Mux_h
    port map (
            O => \N__8168\,
            I => \N__8164\
        );

    \I__1614\ : InMux
    port map (
            O => \N__8167\,
            I => \N__8161\
        );

    \I__1613\ : Odrv12
    port map (
            O => \N__8164\,
            I => \LDSn_c\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__8161\,
            I => \LDSn_c\
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__8156\,
            I => \N__8149\
        );

    \I__1610\ : InMux
    port map (
            O => \N__8155\,
            I => \N__8145\
        );

    \I__1609\ : InMux
    port map (
            O => \N__8154\,
            I => \N__8142\
        );

    \I__1608\ : InMux
    port map (
            O => \N__8153\,
            I => \N__8135\
        );

    \I__1607\ : InMux
    port map (
            O => \N__8152\,
            I => \N__8135\
        );

    \I__1606\ : InMux
    port map (
            O => \N__8149\,
            I => \N__8135\
        );

    \I__1605\ : CascadeMux
    port map (
            O => \N__8148\,
            I => \N__8132\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__8145\,
            I => \N__8125\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__8142\,
            I => \N__8125\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__8135\,
            I => \N__8125\
        );

    \I__1601\ : InMux
    port map (
            O => \N__8132\,
            I => \N__8122\
        );

    \I__1600\ : Span4Mux_v
    port map (
            O => \N__8125\,
            I => \N__8119\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__8122\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1598\ : Odrv4
    port map (
            O => \N__8119\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1597\ : InMux
    port map (
            O => \N__8114\,
            I => \N__8101\
        );

    \I__1596\ : InMux
    port map (
            O => \N__8113\,
            I => \N__8101\
        );

    \I__1595\ : InMux
    port map (
            O => \N__8112\,
            I => \N__8101\
        );

    \I__1594\ : InMux
    port map (
            O => \N__8111\,
            I => \N__8087\
        );

    \I__1593\ : InMux
    port map (
            O => \N__8110\,
            I => \N__8087\
        );

    \I__1592\ : InMux
    port map (
            O => \N__8109\,
            I => \N__8087\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__8108\,
            I => \N__8081\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__8101\,
            I => \N__8077\
        );

    \I__1589\ : InMux
    port map (
            O => \N__8100\,
            I => \N__8074\
        );

    \I__1588\ : InMux
    port map (
            O => \N__8099\,
            I => \N__8065\
        );

    \I__1587\ : InMux
    port map (
            O => \N__8098\,
            I => \N__8065\
        );

    \I__1586\ : InMux
    port map (
            O => \N__8097\,
            I => \N__8065\
        );

    \I__1585\ : InMux
    port map (
            O => \N__8096\,
            I => \N__8065\
        );

    \I__1584\ : InMux
    port map (
            O => \N__8095\,
            I => \N__8062\
        );

    \I__1583\ : InMux
    port map (
            O => \N__8094\,
            I => \N__8058\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__8087\,
            I => \N__8053\
        );

    \I__1581\ : InMux
    port map (
            O => \N__8086\,
            I => \N__8048\
        );

    \I__1580\ : InMux
    port map (
            O => \N__8085\,
            I => \N__8048\
        );

    \I__1579\ : InMux
    port map (
            O => \N__8084\,
            I => \N__8040\
        );

    \I__1578\ : InMux
    port map (
            O => \N__8081\,
            I => \N__8040\
        );

    \I__1577\ : InMux
    port map (
            O => \N__8080\,
            I => \N__8040\
        );

    \I__1576\ : Span4Mux_v
    port map (
            O => \N__8077\,
            I => \N__8031\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__8074\,
            I => \N__8031\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__8065\,
            I => \N__8028\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__8062\,
            I => \N__8025\
        );

    \I__1572\ : InMux
    port map (
            O => \N__8061\,
            I => \N__8022\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__8058\,
            I => \N__8019\
        );

    \I__1570\ : InMux
    port map (
            O => \N__8057\,
            I => \N__8014\
        );

    \I__1569\ : InMux
    port map (
            O => \N__8056\,
            I => \N__8014\
        );

    \I__1568\ : Span4Mux_v
    port map (
            O => \N__8053\,
            I => \N__8009\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__8048\,
            I => \N__8009\
        );

    \I__1566\ : InMux
    port map (
            O => \N__8047\,
            I => \N__8006\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__8040\,
            I => \N__8003\
        );

    \I__1564\ : InMux
    port map (
            O => \N__8039\,
            I => \N__8000\
        );

    \I__1563\ : InMux
    port map (
            O => \N__8038\,
            I => \N__7995\
        );

    \I__1562\ : InMux
    port map (
            O => \N__8037\,
            I => \N__7995\
        );

    \I__1561\ : InMux
    port map (
            O => \N__8036\,
            I => \N__7992\
        );

    \I__1560\ : Span4Mux_v
    port map (
            O => \N__8031\,
            I => \N__7989\
        );

    \I__1559\ : Span4Mux_v
    port map (
            O => \N__8028\,
            I => \N__7984\
        );

    \I__1558\ : Span4Mux_v
    port map (
            O => \N__8025\,
            I => \N__7984\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__8022\,
            I => \N__7981\
        );

    \I__1556\ : Span4Mux_v
    port map (
            O => \N__8019\,
            I => \N__7976\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__8014\,
            I => \N__7976\
        );

    \I__1554\ : Span4Mux_h
    port map (
            O => \N__8009\,
            I => \N__7971\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__8006\,
            I => \N__7971\
        );

    \I__1552\ : Span4Mux_v
    port map (
            O => \N__8003\,
            I => \N__7964\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__8000\,
            I => \N__7964\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__7995\,
            I => \N__7964\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__7992\,
            I => \N__7960\
        );

    \I__1548\ : Span4Mux_h
    port map (
            O => \N__7989\,
            I => \N__7953\
        );

    \I__1547\ : Span4Mux_h
    port map (
            O => \N__7984\,
            I => \N__7953\
        );

    \I__1546\ : Span4Mux_v
    port map (
            O => \N__7981\,
            I => \N__7953\
        );

    \I__1545\ : Span4Mux_v
    port map (
            O => \N__7976\,
            I => \N__7946\
        );

    \I__1544\ : Span4Mux_v
    port map (
            O => \N__7971\,
            I => \N__7946\
        );

    \I__1543\ : Span4Mux_v
    port map (
            O => \N__7964\,
            I => \N__7946\
        );

    \I__1542\ : InMux
    port map (
            O => \N__7963\,
            I => \N__7943\
        );

    \I__1541\ : Span12Mux_v
    port map (
            O => \N__7960\,
            I => \N__7936\
        );

    \I__1540\ : Sp12to4
    port map (
            O => \N__7953\,
            I => \N__7936\
        );

    \I__1539\ : Sp12to4
    port map (
            O => \N__7946\,
            I => \N__7936\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7943\,
            I => \N__7933\
        );

    \I__1537\ : Span12Mux_h
    port map (
            O => \N__7936\,
            I => \N__7930\
        );

    \I__1536\ : Span12Mux_h
    port map (
            O => \N__7933\,
            I => \N__7927\
        );

    \I__1535\ : Odrv12
    port map (
            O => \N__7930\,
            I => \RESETn_c\
        );

    \I__1534\ : Odrv12
    port map (
            O => \N__7927\,
            I => \RESETn_c\
        );

    \I__1533\ : IoInMux
    port map (
            O => \N__7922\,
            I => \N__7919\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__7919\,
            I => \N__7916\
        );

    \I__1531\ : Span12Mux_s7_v
    port map (
            O => \N__7916\,
            I => \N__7913\
        );

    \I__1530\ : Odrv12
    port map (
            O => \N__7913\,
            I => \RESETn_c_i\
        );

    \I__1529\ : IoInMux
    port map (
            O => \N__7910\,
            I => \N__7907\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__7907\,
            I => \N__7904\
        );

    \I__1527\ : Span4Mux_s3_v
    port map (
            O => \N__7904\,
            I => \N__7901\
        );

    \I__1526\ : Span4Mux_v
    port map (
            O => \N__7901\,
            I => \N__7898\
        );

    \I__1525\ : Span4Mux_h
    port map (
            O => \N__7898\,
            I => \N__7895\
        );

    \I__1524\ : Odrv4
    port map (
            O => \N__7895\,
            I => \RASn_c\
        );

    \I__1523\ : InMux
    port map (
            O => \N__7892\,
            I => \N__7889\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__7889\,
            I => \U712_CHIP_RAM.d_N_7\
        );

    \I__1521\ : InMux
    port map (
            O => \N__7886\,
            I => \N__7883\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__7883\,
            I => \U712_CHIP_RAM.m185_0\
        );

    \I__1519\ : InMux
    port map (
            O => \N__7880\,
            I => \N__7877\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__7877\,
            I => \N__7874\
        );

    \I__1517\ : Sp12to4
    port map (
            O => \N__7874\,
            I => \N__7871\
        );

    \I__1516\ : Span12Mux_v
    port map (
            O => \N__7871\,
            I => \N__7868\
        );

    \I__1515\ : Span12Mux_h
    port map (
            O => \N__7868\,
            I => \N__7865\
        );

    \I__1514\ : Odrv12
    port map (
            O => \N__7865\,
            I => \A_c_16\
        );

    \I__1513\ : InMux
    port map (
            O => \N__7862\,
            I => \N__7858\
        );

    \I__1512\ : InMux
    port map (
            O => \N__7861\,
            I => \N__7855\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__7858\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__7855\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\
        );

    \I__1509\ : InMux
    port map (
            O => \N__7850\,
            I => \N__7844\
        );

    \I__1508\ : InMux
    port map (
            O => \N__7849\,
            I => \N__7844\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__7844\,
            I => \N__7841\
        );

    \I__1506\ : Span4Mux_v
    port map (
            O => \N__7841\,
            I => \N__7837\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7840\,
            I => \N__7834\
        );

    \I__1504\ : Sp12to4
    port map (
            O => \N__7837\,
            I => \N__7829\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7834\,
            I => \N__7829\
        );

    \I__1502\ : Span12Mux_h
    port map (
            O => \N__7829\,
            I => \N__7826\
        );

    \I__1501\ : Odrv12
    port map (
            O => \N__7826\,
            I => \AWEn_c\
        );

    \I__1500\ : CascadeMux
    port map (
            O => \N__7823\,
            I => \N__7820\
        );

    \I__1499\ : InMux
    port map (
            O => \N__7820\,
            I => \N__7817\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__7817\,
            I => \N__7813\
        );

    \I__1497\ : CascadeMux
    port map (
            O => \N__7816\,
            I => \N__7810\
        );

    \I__1496\ : Span4Mux_v
    port map (
            O => \N__7813\,
            I => \N__7806\
        );

    \I__1495\ : InMux
    port map (
            O => \N__7810\,
            I => \N__7803\
        );

    \I__1494\ : InMux
    port map (
            O => \N__7809\,
            I => \N__7796\
        );

    \I__1493\ : Sp12to4
    port map (
            O => \N__7806\,
            I => \N__7791\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__7803\,
            I => \N__7791\
        );

    \I__1491\ : InMux
    port map (
            O => \N__7802\,
            I => \N__7786\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7801\,
            I => \N__7786\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7800\,
            I => \N__7781\
        );

    \I__1488\ : InMux
    port map (
            O => \N__7799\,
            I => \N__7781\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__7796\,
            I => \U712_CHIP_RAM.N_26_0\
        );

    \I__1486\ : Odrv12
    port map (
            O => \N__7791\,
            I => \U712_CHIP_RAM.N_26_0\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__7786\,
            I => \U712_CHIP_RAM.N_26_0\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__7781\,
            I => \U712_CHIP_RAM.N_26_0\
        );

    \I__1483\ : CascadeMux
    port map (
            O => \N__7772\,
            I => \N__7767\
        );

    \I__1482\ : InMux
    port map (
            O => \N__7771\,
            I => \N__7763\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7770\,
            I => \N__7760\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7767\,
            I => \N__7757\
        );

    \I__1479\ : CascadeMux
    port map (
            O => \N__7766\,
            I => \N__7753\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__7763\,
            I => \N__7741\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__7760\,
            I => \N__7741\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__7757\,
            I => \N__7738\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7756\,
            I => \N__7727\
        );

    \I__1474\ : InMux
    port map (
            O => \N__7753\,
            I => \N__7727\
        );

    \I__1473\ : InMux
    port map (
            O => \N__7752\,
            I => \N__7727\
        );

    \I__1472\ : InMux
    port map (
            O => \N__7751\,
            I => \N__7727\
        );

    \I__1471\ : InMux
    port map (
            O => \N__7750\,
            I => \N__7727\
        );

    \I__1470\ : InMux
    port map (
            O => \N__7749\,
            I => \N__7721\
        );

    \I__1469\ : InMux
    port map (
            O => \N__7748\,
            I => \N__7718\
        );

    \I__1468\ : InMux
    port map (
            O => \N__7747\,
            I => \N__7713\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7746\,
            I => \N__7713\
        );

    \I__1466\ : Span4Mux_h
    port map (
            O => \N__7741\,
            I => \N__7710\
        );

    \I__1465\ : Span4Mux_h
    port map (
            O => \N__7738\,
            I => \N__7705\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__7727\,
            I => \N__7705\
        );

    \I__1463\ : InMux
    port map (
            O => \N__7726\,
            I => \N__7698\
        );

    \I__1462\ : InMux
    port map (
            O => \N__7725\,
            I => \N__7698\
        );

    \I__1461\ : InMux
    port map (
            O => \N__7724\,
            I => \N__7698\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__7721\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__7718\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__7713\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1457\ : Odrv4
    port map (
            O => \N__7710\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1456\ : Odrv4
    port map (
            O => \N__7705\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__7698\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1454\ : CascadeMux
    port map (
            O => \N__7685\,
            I => \N__7682\
        );

    \I__1453\ : InMux
    port map (
            O => \N__7682\,
            I => \N__7676\
        );

    \I__1452\ : InMux
    port map (
            O => \N__7681\,
            I => \N__7673\
        );

    \I__1451\ : InMux
    port map (
            O => \N__7680\,
            I => \N__7670\
        );

    \I__1450\ : InMux
    port map (
            O => \N__7679\,
            I => \N__7667\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__7676\,
            I => \N__7663\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__7673\,
            I => \N__7660\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__7670\,
            I => \N__7655\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__7667\,
            I => \N__7655\
        );

    \I__1445\ : InMux
    port map (
            O => \N__7666\,
            I => \N__7652\
        );

    \I__1444\ : Odrv12
    port map (
            O => \N__7663\,
            I => \U712_CHIP_RAM.N_30_0\
        );

    \I__1443\ : Odrv4
    port map (
            O => \N__7660\,
            I => \U712_CHIP_RAM.N_30_0\
        );

    \I__1442\ : Odrv4
    port map (
            O => \N__7655\,
            I => \U712_CHIP_RAM.N_30_0\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__7652\,
            I => \U712_CHIP_RAM.N_30_0\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__7643\,
            I => \U712_CHIP_RAM.N_62_0_cascade_\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7640\,
            I => \N__7637\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__7637\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_RNI9THUZ0Z5\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__7634\,
            I => \U712_CHIP_RAM.CLK_EN_RNOZ0Z_2_cascade_\
        );

    \I__1436\ : InMux
    port map (
            O => \N__7631\,
            I => \N__7628\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__7628\,
            I => \N__7625\
        );

    \I__1434\ : Odrv4
    port map (
            O => \N__7625\,
            I => \U712_CHIP_RAM.CLK_EN_RNOZ0Z_3\
        );

    \I__1433\ : CascadeMux
    port map (
            O => \N__7622\,
            I => \U712_CHIP_RAM.N_174_0_cascade_\
        );

    \I__1432\ : InMux
    port map (
            O => \N__7619\,
            I => \N__7616\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__7616\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER43\
        );

    \I__1430\ : IoInMux
    port map (
            O => \N__7613\,
            I => \N__7610\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__7610\,
            I => \N__7607\
        );

    \I__1428\ : Span4Mux_s1_h
    port map (
            O => \N__7607\,
            I => \N__7604\
        );

    \I__1427\ : Sp12to4
    port map (
            O => \N__7604\,
            I => \N__7601\
        );

    \I__1426\ : Span12Mux_v
    port map (
            O => \N__7601\,
            I => \N__7598\
        );

    \I__1425\ : Span12Mux_h
    port map (
            O => \N__7598\,
            I => \N__7594\
        );

    \I__1424\ : InMux
    port map (
            O => \N__7597\,
            I => \N__7591\
        );

    \I__1423\ : Odrv12
    port map (
            O => \N__7594\,
            I => \CLK_EN_c\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__7591\,
            I => \CLK_EN_c\
        );

    \I__1421\ : CascadeMux
    port map (
            O => \N__7586\,
            I => \N__7583\
        );

    \I__1420\ : InMux
    port map (
            O => \N__7583\,
            I => \N__7575\
        );

    \I__1419\ : InMux
    port map (
            O => \N__7582\,
            I => \N__7568\
        );

    \I__1418\ : InMux
    port map (
            O => \N__7581\,
            I => \N__7568\
        );

    \I__1417\ : InMux
    port map (
            O => \N__7580\,
            I => \N__7568\
        );

    \I__1416\ : CascadeMux
    port map (
            O => \N__7579\,
            I => \N__7565\
        );

    \I__1415\ : CascadeMux
    port map (
            O => \N__7578\,
            I => \N__7561\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__7575\,
            I => \N__7558\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__7568\,
            I => \N__7555\
        );

    \I__1412\ : InMux
    port map (
            O => \N__7565\,
            I => \N__7552\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7564\,
            I => \N__7549\
        );

    \I__1410\ : InMux
    port map (
            O => \N__7561\,
            I => \N__7546\
        );

    \I__1409\ : Span4Mux_v
    port map (
            O => \N__7558\,
            I => \N__7543\
        );

    \I__1408\ : Span4Mux_v
    port map (
            O => \N__7555\,
            I => \N__7538\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__7552\,
            I => \N__7538\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__7549\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__7546\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1404\ : Odrv4
    port map (
            O => \N__7543\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1403\ : Odrv4
    port map (
            O => \N__7538\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__7529\,
            I => \N__7525\
        );

    \I__1401\ : CascadeMux
    port map (
            O => \N__7528\,
            I => \N__7521\
        );

    \I__1400\ : InMux
    port map (
            O => \N__7525\,
            I => \N__7518\
        );

    \I__1399\ : InMux
    port map (
            O => \N__7524\,
            I => \N__7515\
        );

    \I__1398\ : InMux
    port map (
            O => \N__7521\,
            I => \N__7512\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__7518\,
            I => \U712_CHIP_RAM.N_62_0\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__7515\,
            I => \U712_CHIP_RAM.N_62_0\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__7512\,
            I => \U712_CHIP_RAM.N_62_0\
        );

    \I__1394\ : InMux
    port map (
            O => \N__7505\,
            I => \N__7500\
        );

    \I__1393\ : InMux
    port map (
            O => \N__7504\,
            I => \N__7494\
        );

    \I__1392\ : InMux
    port map (
            O => \N__7503\,
            I => \N__7494\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__7500\,
            I => \N__7491\
        );

    \I__1390\ : InMux
    port map (
            O => \N__7499\,
            I => \N__7488\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__7494\,
            I => \U712_CHIP_RAM.N_52_0\
        );

    \I__1388\ : Odrv4
    port map (
            O => \N__7491\,
            I => \U712_CHIP_RAM.N_52_0\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__7488\,
            I => \U712_CHIP_RAM.N_52_0\
        );

    \I__1386\ : InMux
    port map (
            O => \N__7481\,
            I => \N__7478\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__7478\,
            I => \N__7475\
        );

    \I__1384\ : Span4Mux_v
    port map (
            O => \N__7475\,
            I => \N__7472\
        );

    \I__1383\ : Sp12to4
    port map (
            O => \N__7472\,
            I => \N__7469\
        );

    \I__1382\ : Span12Mux_h
    port map (
            O => \N__7469\,
            I => \N__7466\
        );

    \I__1381\ : Odrv12
    port map (
            O => \N__7466\,
            I => \A_c_4\
        );

    \I__1380\ : CascadeMux
    port map (
            O => \N__7463\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_\
        );

    \I__1379\ : InMux
    port map (
            O => \N__7460\,
            I => \N__7456\
        );

    \I__1378\ : InMux
    port map (
            O => \N__7459\,
            I => \N__7453\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__7456\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__7453\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\
        );

    \I__1375\ : InMux
    port map (
            O => \N__7448\,
            I => \N__7445\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__7445\,
            I => \N__7442\
        );

    \I__1373\ : Span4Mux_v
    port map (
            O => \N__7442\,
            I => \N__7439\
        );

    \I__1372\ : Sp12to4
    port map (
            O => \N__7439\,
            I => \N__7436\
        );

    \I__1371\ : Span12Mux_h
    port map (
            O => \N__7436\,
            I => \N__7433\
        );

    \I__1370\ : Odrv12
    port map (
            O => \N__7433\,
            I => \A_c_5\
        );

    \I__1369\ : InMux
    port map (
            O => \N__7430\,
            I => \N__7426\
        );

    \I__1368\ : InMux
    port map (
            O => \N__7429\,
            I => \N__7423\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__7426\,
            I => \N__7420\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__7423\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\
        );

    \I__1365\ : Odrv12
    port map (
            O => \N__7420\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\
        );

    \I__1364\ : InMux
    port map (
            O => \N__7415\,
            I => \N__7412\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__7412\,
            I => \N__7409\
        );

    \I__1362\ : Span4Mux_v
    port map (
            O => \N__7409\,
            I => \N__7406\
        );

    \I__1361\ : Sp12to4
    port map (
            O => \N__7406\,
            I => \N__7403\
        );

    \I__1360\ : Span12Mux_h
    port map (
            O => \N__7403\,
            I => \N__7400\
        );

    \I__1359\ : Odrv12
    port map (
            O => \N__7400\,
            I => \A_c_6\
        );

    \I__1358\ : InMux
    port map (
            O => \N__7397\,
            I => \N__7394\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__7394\,
            I => \N__7390\
        );

    \I__1356\ : InMux
    port map (
            O => \N__7393\,
            I => \N__7387\
        );

    \I__1355\ : Span4Mux_v
    port map (
            O => \N__7390\,
            I => \N__7384\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__7387\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\
        );

    \I__1353\ : Odrv4
    port map (
            O => \N__7384\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\
        );

    \I__1352\ : InMux
    port map (
            O => \N__7379\,
            I => \N__7376\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__7376\,
            I => \N__7373\
        );

    \I__1350\ : Span12Mux_v
    port map (
            O => \N__7373\,
            I => \N__7370\
        );

    \I__1349\ : Span12Mux_h
    port map (
            O => \N__7370\,
            I => \N__7367\
        );

    \I__1348\ : Odrv12
    port map (
            O => \N__7367\,
            I => \A_c_7\
        );

    \I__1347\ : InMux
    port map (
            O => \N__7364\,
            I => \N__7361\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__7361\,
            I => \N__7357\
        );

    \I__1345\ : InMux
    port map (
            O => \N__7360\,
            I => \N__7354\
        );

    \I__1344\ : Span4Mux_v
    port map (
            O => \N__7357\,
            I => \N__7351\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__7354\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\
        );

    \I__1342\ : Odrv4
    port map (
            O => \N__7351\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\
        );

    \I__1341\ : CascadeMux
    port map (
            O => \N__7346\,
            I => \U712_CHIP_RAM.DMA_CYCLE_START_RNIJD6OZ0Z3_cascade_\
        );

    \I__1340\ : CascadeMux
    port map (
            O => \N__7343\,
            I => \U712_CHIP_RAM.N_204_cascade_\
        );

    \I__1339\ : InMux
    port map (
            O => \N__7340\,
            I => \N__7337\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__7337\,
            I => \N__7332\
        );

    \I__1337\ : InMux
    port map (
            O => \N__7336\,
            I => \N__7329\
        );

    \I__1336\ : InMux
    port map (
            O => \N__7335\,
            I => \N__7326\
        );

    \I__1335\ : Span4Mux_v
    port map (
            O => \N__7332\,
            I => \N__7320\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__7329\,
            I => \N__7320\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__7326\,
            I => \N__7317\
        );

    \I__1332\ : InMux
    port map (
            O => \N__7325\,
            I => \N__7314\
        );

    \I__1331\ : Span4Mux_h
    port map (
            O => \N__7320\,
            I => \N__7311\
        );

    \I__1330\ : Odrv4
    port map (
            O => \N__7317\,
            I => \U712_CHIP_RAM.N_364\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__7314\,
            I => \U712_CHIP_RAM.N_364\
        );

    \I__1328\ : Odrv4
    port map (
            O => \N__7311\,
            I => \U712_CHIP_RAM.N_364\
        );

    \I__1327\ : InMux
    port map (
            O => \N__7304\,
            I => \N__7300\
        );

    \I__1326\ : InMux
    port map (
            O => \N__7303\,
            I => \N__7294\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__7300\,
            I => \N__7291\
        );

    \I__1324\ : InMux
    port map (
            O => \N__7299\,
            I => \N__7286\
        );

    \I__1323\ : InMux
    port map (
            O => \N__7298\,
            I => \N__7286\
        );

    \I__1322\ : InMux
    port map (
            O => \N__7297\,
            I => \N__7283\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__7294\,
            I => \N__7276\
        );

    \I__1320\ : Span4Mux_v
    port map (
            O => \N__7291\,
            I => \N__7273\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__7286\,
            I => \N__7268\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__7283\,
            I => \N__7268\
        );

    \I__1317\ : InMux
    port map (
            O => \N__7282\,
            I => \N__7265\
        );

    \I__1316\ : InMux
    port map (
            O => \N__7281\,
            I => \N__7262\
        );

    \I__1315\ : InMux
    port map (
            O => \N__7280\,
            I => \N__7257\
        );

    \I__1314\ : InMux
    port map (
            O => \N__7279\,
            I => \N__7257\
        );

    \I__1313\ : Span4Mux_h
    port map (
            O => \N__7276\,
            I => \N__7254\
        );

    \I__1312\ : Span4Mux_h
    port map (
            O => \N__7273\,
            I => \N__7249\
        );

    \I__1311\ : Span4Mux_h
    port map (
            O => \N__7268\,
            I => \N__7249\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__7265\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__7262\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__7257\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1307\ : Odrv4
    port map (
            O => \N__7254\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1306\ : Odrv4
    port map (
            O => \N__7249\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__7238\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_\
        );

    \I__1304\ : IoInMux
    port map (
            O => \N__7235\,
            I => \N__7232\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__7232\,
            I => \N__7229\
        );

    \I__1302\ : Span4Mux_s2_v
    port map (
            O => \N__7229\,
            I => \N__7226\
        );

    \I__1301\ : Span4Mux_v
    port map (
            O => \N__7226\,
            I => \N__7223\
        );

    \I__1300\ : Span4Mux_h
    port map (
            O => \N__7223\,
            I => \N__7220\
        );

    \I__1299\ : Sp12to4
    port map (
            O => \N__7220\,
            I => \N__7217\
        );

    \I__1298\ : Span12Mux_v
    port map (
            O => \N__7217\,
            I => \N__7213\
        );

    \I__1297\ : InMux
    port map (
            O => \N__7216\,
            I => \N__7210\
        );

    \I__1296\ : Odrv12
    port map (
            O => \N__7213\,
            I => \DBDIR_c\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__7210\,
            I => \DBDIR_c\
        );

    \I__1294\ : IoInMux
    port map (
            O => \N__7205\,
            I => \N__7202\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__7202\,
            I => \N__7199\
        );

    \I__1292\ : IoSpan4Mux
    port map (
            O => \N__7199\,
            I => \N__7196\
        );

    \I__1291\ : Span4Mux_s2_v
    port map (
            O => \N__7196\,
            I => \N__7193\
        );

    \I__1290\ : Sp12to4
    port map (
            O => \N__7193\,
            I => \N__7189\
        );

    \I__1289\ : InMux
    port map (
            O => \N__7192\,
            I => \N__7186\
        );

    \I__1288\ : Span12Mux_s8_v
    port map (
            O => \N__7189\,
            I => \N__7183\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__7186\,
            I => \N__7180\
        );

    \I__1286\ : Span12Mux_v
    port map (
            O => \N__7183\,
            I => \N__7177\
        );

    \I__1285\ : Span12Mux_v
    port map (
            O => \N__7180\,
            I => \N__7174\
        );

    \I__1284\ : Span12Mux_h
    port map (
            O => \N__7177\,
            I => \N__7171\
        );

    \I__1283\ : Span12Mux_h
    port map (
            O => \N__7174\,
            I => \N__7168\
        );

    \I__1282\ : Odrv12
    port map (
            O => \N__7171\,
            I => \A_c_11\
        );

    \I__1281\ : Odrv12
    port map (
            O => \N__7168\,
            I => \A_c_11\
        );

    \I__1280\ : CascadeMux
    port map (
            O => \N__7163\,
            I => \U712_CHIP_RAM.N_3_0_cascade_\
        );

    \I__1279\ : InMux
    port map (
            O => \N__7160\,
            I => \N__7157\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__7157\,
            I => \U712_CHIP_RAM.m187_0\
        );

    \I__1277\ : InMux
    port map (
            O => \N__7154\,
            I => \N__7151\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__7151\,
            I => \N__7148\
        );

    \I__1275\ : Span4Mux_h
    port map (
            O => \N__7148\,
            I => \N__7145\
        );

    \I__1274\ : Odrv4
    port map (
            O => \N__7145\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_1\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__7142\,
            I => \U712_CHIP_RAM.N_163_0_cascade_\
        );

    \I__1272\ : InMux
    port map (
            O => \N__7139\,
            I => \N__7133\
        );

    \I__1271\ : InMux
    port map (
            O => \N__7138\,
            I => \N__7130\
        );

    \I__1270\ : InMux
    port map (
            O => \N__7137\,
            I => \N__7125\
        );

    \I__1269\ : InMux
    port map (
            O => \N__7136\,
            I => \N__7125\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__7133\,
            I => \U712_CHIP_RAM.N_67_0\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__7130\,
            I => \U712_CHIP_RAM.N_67_0\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__7125\,
            I => \U712_CHIP_RAM.N_67_0\
        );

    \I__1265\ : SRMux
    port map (
            O => \N__7118\,
            I => \N__7115\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__7115\,
            I => \N__7112\
        );

    \I__1263\ : Span4Mux_v
    port map (
            O => \N__7112\,
            I => \N__7109\
        );

    \I__1262\ : Span4Mux_h
    port map (
            O => \N__7109\,
            I => \N__7106\
        );

    \I__1261\ : Odrv4
    port map (
            O => \N__7106\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__1260\ : InMux
    port map (
            O => \N__7103\,
            I => \N__7100\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__7100\,
            I => \N__7097\
        );

    \I__1258\ : Span4Mux_h
    port map (
            O => \N__7097\,
            I => \N__7090\
        );

    \I__1257\ : InMux
    port map (
            O => \N__7096\,
            I => \N__7087\
        );

    \I__1256\ : InMux
    port map (
            O => \N__7095\,
            I => \N__7084\
        );

    \I__1255\ : InMux
    port map (
            O => \N__7094\,
            I => \N__7079\
        );

    \I__1254\ : InMux
    port map (
            O => \N__7093\,
            I => \N__7079\
        );

    \I__1253\ : Odrv4
    port map (
            O => \N__7090\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__7087\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__7084\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__7079\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1249\ : InMux
    port map (
            O => \N__7070\,
            I => \N__7064\
        );

    \I__1248\ : InMux
    port map (
            O => \N__7069\,
            I => \N__7061\
        );

    \I__1247\ : InMux
    port map (
            O => \N__7068\,
            I => \N__7056\
        );

    \I__1246\ : InMux
    port map (
            O => \N__7067\,
            I => \N__7056\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__7064\,
            I => \N__7051\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__7061\,
            I => \N__7051\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__7056\,
            I => \U712_CHIP_RAM.N_48_0\
        );

    \I__1242\ : Odrv4
    port map (
            O => \N__7051\,
            I => \U712_CHIP_RAM.N_48_0\
        );

    \I__1241\ : InMux
    port map (
            O => \N__7046\,
            I => \N__7043\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__7043\,
            I => \N__7039\
        );

    \I__1239\ : InMux
    port map (
            O => \N__7042\,
            I => \N__7036\
        );

    \I__1238\ : Span4Mux_h
    port map (
            O => \N__7039\,
            I => \N__7033\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__7036\,
            I => \U712_CHIP_RAM.N_363\
        );

    \I__1236\ : Odrv4
    port map (
            O => \N__7033\,
            I => \U712_CHIP_RAM.N_363\
        );

    \I__1235\ : CascadeMux
    port map (
            O => \N__7028\,
            I => \U712_CHIP_RAM.N_158_0_cascade_\
        );

    \I__1234\ : InMux
    port map (
            O => \N__7025\,
            I => \N__7019\
        );

    \I__1233\ : InMux
    port map (
            O => \N__7024\,
            I => \N__7010\
        );

    \I__1232\ : InMux
    port map (
            O => \N__7023\,
            I => \N__7010\
        );

    \I__1231\ : InMux
    port map (
            O => \N__7022\,
            I => \N__7010\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__7019\,
            I => \N__7007\
        );

    \I__1229\ : InMux
    port map (
            O => \N__7018\,
            I => \N__7002\
        );

    \I__1228\ : InMux
    port map (
            O => \N__7017\,
            I => \N__7002\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__7010\,
            I => \U712_CHIP_RAM.N_58_0\
        );

    \I__1226\ : Odrv4
    port map (
            O => \N__7007\,
            I => \U712_CHIP_RAM.N_58_0\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__7002\,
            I => \U712_CHIP_RAM.N_58_0\
        );

    \I__1224\ : InMux
    port map (
            O => \N__6995\,
            I => \N__6992\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__6992\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_1\
        );

    \I__1222\ : InMux
    port map (
            O => \N__6989\,
            I => \N__6986\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__6986\,
            I => \N__6983\
        );

    \I__1220\ : Odrv4
    port map (
            O => \N__6983\,
            I => \U712_CHIP_RAM.d_N_6_0\
        );

    \I__1219\ : InMux
    port map (
            O => \N__6980\,
            I => \N__6977\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__6977\,
            I => \N__6972\
        );

    \I__1217\ : InMux
    port map (
            O => \N__6976\,
            I => \N__6969\
        );

    \I__1216\ : InMux
    port map (
            O => \N__6975\,
            I => \N__6966\
        );

    \I__1215\ : Odrv4
    port map (
            O => \N__6972\,
            I => \U712_CHIP_RAM.N_43_0\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__6969\,
            I => \U712_CHIP_RAM.N_43_0\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__6966\,
            I => \U712_CHIP_RAM.N_43_0\
        );

    \I__1212\ : CascadeMux
    port map (
            O => \N__6959\,
            I => \N__6956\
        );

    \I__1211\ : InMux
    port map (
            O => \N__6956\,
            I => \N__6953\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__6953\,
            I => \U712_CHIP_RAM.m189_0\
        );

    \I__1209\ : InMux
    port map (
            O => \N__6950\,
            I => \N__6947\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__6947\,
            I => \N__6944\
        );

    \I__1207\ : Span4Mux_h
    port map (
            O => \N__6944\,
            I => \N__6941\
        );

    \I__1206\ : Sp12to4
    port map (
            O => \N__6941\,
            I => \N__6938\
        );

    \I__1205\ : Span12Mux_v
    port map (
            O => \N__6938\,
            I => \N__6935\
        );

    \I__1204\ : Span12Mux_h
    port map (
            O => \N__6935\,
            I => \N__6932\
        );

    \I__1203\ : Odrv12
    port map (
            O => \N__6932\,
            I => \A_c_14\
        );

    \I__1202\ : IoInMux
    port map (
            O => \N__6929\,
            I => \N__6926\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__6926\,
            I => \N__6923\
        );

    \I__1200\ : IoSpan4Mux
    port map (
            O => \N__6923\,
            I => \N__6920\
        );

    \I__1199\ : Span4Mux_s0_v
    port map (
            O => \N__6920\,
            I => \N__6917\
        );

    \I__1198\ : Sp12to4
    port map (
            O => \N__6917\,
            I => \N__6914\
        );

    \I__1197\ : Odrv12
    port map (
            O => \N__6914\,
            I => \CMA_c_2\
        );

    \I__1196\ : InMux
    port map (
            O => \N__6911\,
            I => \N__6908\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__6908\,
            I => \U712_CHIP_RAM.m186_1\
        );

    \I__1194\ : IoInMux
    port map (
            O => \N__6905\,
            I => \N__6902\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__6902\,
            I => \N__6899\
        );

    \I__1192\ : Span4Mux_s1_v
    port map (
            O => \N__6899\,
            I => \N__6896\
        );

    \I__1191\ : Span4Mux_v
    port map (
            O => \N__6896\,
            I => \N__6893\
        );

    \I__1190\ : Sp12to4
    port map (
            O => \N__6893\,
            I => \N__6890\
        );

    \I__1189\ : Span12Mux_h
    port map (
            O => \N__6890\,
            I => \N__6887\
        );

    \I__1188\ : Odrv12
    port map (
            O => \N__6887\,
            I => \CMA_c_0\
        );

    \I__1187\ : IoInMux
    port map (
            O => \N__6884\,
            I => \N__6881\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__6881\,
            I => \N__6878\
        );

    \I__1185\ : Span12Mux_s7_v
    port map (
            O => \N__6878\,
            I => \N__6875\
        );

    \I__1184\ : Odrv12
    port map (
            O => \N__6875\,
            I => \CMA_c_1\
        );

    \I__1183\ : CascadeMux
    port map (
            O => \N__6872\,
            I => \U712_CHIP_RAM.N_198_cascade_\
        );

    \I__1182\ : ClkMux
    port map (
            O => \N__6869\,
            I => \N__6864\
        );

    \I__1181\ : InMux
    port map (
            O => \N__6868\,
            I => \N__6861\
        );

    \I__1180\ : ClkMux
    port map (
            O => \N__6867\,
            I => \N__6858\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__6864\,
            I => \N__6855\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__6861\,
            I => \N__6852\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__6858\,
            I => \N__6849\
        );

    \I__1176\ : Span4Mux_h
    port map (
            O => \N__6855\,
            I => \N__6842\
        );

    \I__1175\ : Span4Mux_v
    port map (
            O => \N__6852\,
            I => \N__6842\
        );

    \I__1174\ : Span4Mux_h
    port map (
            O => \N__6849\,
            I => \N__6842\
        );

    \I__1173\ : Span4Mux_v
    port map (
            O => \N__6842\,
            I => \N__6839\
        );

    \I__1172\ : Span4Mux_v
    port map (
            O => \N__6839\,
            I => \N__6836\
        );

    \I__1171\ : Odrv4
    port map (
            O => \N__6836\,
            I => \CLK40_PLL\
        );

    \I__1170\ : IoInMux
    port map (
            O => \N__6833\,
            I => \N__6828\
        );

    \I__1169\ : IoInMux
    port map (
            O => \N__6832\,
            I => \N__6825\
        );

    \I__1168\ : IoInMux
    port map (
            O => \N__6831\,
            I => \N__6822\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__6828\,
            I => \N__6819\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__6825\,
            I => \N__6816\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__6822\,
            I => \N__6813\
        );

    \I__1164\ : IoSpan4Mux
    port map (
            O => \N__6819\,
            I => \N__6810\
        );

    \I__1163\ : IoSpan4Mux
    port map (
            O => \N__6816\,
            I => \N__6807\
        );

    \I__1162\ : Span12Mux_s6_v
    port map (
            O => \N__6813\,
            I => \N__6804\
        );

    \I__1161\ : Sp12to4
    port map (
            O => \N__6810\,
            I => \N__6801\
        );

    \I__1160\ : Span4Mux_s2_h
    port map (
            O => \N__6807\,
            I => \N__6798\
        );

    \I__1159\ : Span12Mux_v
    port map (
            O => \N__6804\,
            I => \N__6795\
        );

    \I__1158\ : Span12Mux_s6_v
    port map (
            O => \N__6801\,
            I => \N__6792\
        );

    \I__1157\ : Sp12to4
    port map (
            O => \N__6798\,
            I => \N__6789\
        );

    \I__1156\ : Span12Mux_h
    port map (
            O => \N__6795\,
            I => \N__6786\
        );

    \I__1155\ : Span12Mux_v
    port map (
            O => \N__6792\,
            I => \N__6781\
        );

    \I__1154\ : Span12Mux_h
    port map (
            O => \N__6789\,
            I => \N__6781\
        );

    \I__1153\ : Odrv12
    port map (
            O => \N__6786\,
            I => \CLK40_PLL_iso_i\
        );

    \I__1152\ : Odrv12
    port map (
            O => \N__6781\,
            I => \CLK40_PLL_iso_i\
        );

    \I__1151\ : InMux
    port map (
            O => \N__6776\,
            I => \N__6773\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__6773\,
            I => \U712_CHIP_RAM.m187_1\
        );

    \I__1149\ : IoInMux
    port map (
            O => \N__6770\,
            I => \N__6767\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__6767\,
            I => \N__6764\
        );

    \I__1147\ : IoSpan4Mux
    port map (
            O => \N__6764\,
            I => \N__6761\
        );

    \I__1146\ : Span4Mux_s3_h
    port map (
            O => \N__6761\,
            I => \N__6758\
        );

    \I__1145\ : Span4Mux_v
    port map (
            O => \N__6758\,
            I => \N__6755\
        );

    \I__1144\ : Span4Mux_h
    port map (
            O => \N__6755\,
            I => \N__6752\
        );

    \I__1143\ : Sp12to4
    port map (
            O => \N__6752\,
            I => \N__6749\
        );

    \I__1142\ : Odrv12
    port map (
            O => \N__6749\,
            I => \CMA_c_4\
        );

    \I__1141\ : IoInMux
    port map (
            O => \N__6746\,
            I => \N__6743\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__6743\,
            I => \N__6740\
        );

    \I__1139\ : Span4Mux_s3_h
    port map (
            O => \N__6740\,
            I => \N__6737\
        );

    \I__1138\ : Span4Mux_v
    port map (
            O => \N__6737\,
            I => \N__6734\
        );

    \I__1137\ : Span4Mux_h
    port map (
            O => \N__6734\,
            I => \N__6731\
        );

    \I__1136\ : Span4Mux_h
    port map (
            O => \N__6731\,
            I => \N__6728\
        );

    \I__1135\ : Span4Mux_h
    port map (
            O => \N__6728\,
            I => \N__6725\
        );

    \I__1134\ : Odrv4
    port map (
            O => \N__6725\,
            I => \CMA_c_3\
        );

    \I__1133\ : IoInMux
    port map (
            O => \N__6722\,
            I => \N__6719\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__6719\,
            I => \N__6716\
        );

    \I__1131\ : Span4Mux_s2_v
    port map (
            O => \N__6716\,
            I => \N__6713\
        );

    \I__1130\ : Sp12to4
    port map (
            O => \N__6713\,
            I => \N__6710\
        );

    \I__1129\ : Span12Mux_h
    port map (
            O => \N__6710\,
            I => \N__6707\
        );

    \I__1128\ : Odrv12
    port map (
            O => \N__6707\,
            I => \CMA_c_10\
        );

    \I__1127\ : InMux
    port map (
            O => \N__6704\,
            I => \N__6701\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__6701\,
            I => \U712_CHIP_RAM.m189_1\
        );

    \I__1125\ : InMux
    port map (
            O => \N__6698\,
            I => \N__6695\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__6695\,
            I => \U712_CHIP_RAM.m188_1\
        );

    \I__1123\ : InMux
    port map (
            O => \N__6692\,
            I => \N__6689\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__6689\,
            I => \U712_CHIP_RAM.d_N_6_2\
        );

    \I__1121\ : InMux
    port map (
            O => \N__6686\,
            I => \N__6683\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__6683\,
            I => \N__6680\
        );

    \I__1119\ : Span4Mux_v
    port map (
            O => \N__6680\,
            I => \N__6677\
        );

    \I__1118\ : Sp12to4
    port map (
            O => \N__6677\,
            I => \N__6674\
        );

    \I__1117\ : Span12Mux_h
    port map (
            O => \N__6674\,
            I => \N__6671\
        );

    \I__1116\ : Odrv12
    port map (
            O => \N__6671\,
            I => \A_c_12\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6668\,
            I => \N__6665\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__6665\,
            I => \U712_CHIP_RAM.m188_0\
        );

    \I__1113\ : InMux
    port map (
            O => \N__6662\,
            I => \N__6659\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__6659\,
            I => \U712_CHIP_RAM.d_N_6\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6656\,
            I => \N__6653\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6653\,
            I => \N__6650\
        );

    \I__1109\ : Span12Mux_v
    port map (
            O => \N__6650\,
            I => \N__6647\
        );

    \I__1108\ : Span12Mux_h
    port map (
            O => \N__6647\,
            I => \N__6644\
        );

    \I__1107\ : Odrv12
    port map (
            O => \N__6644\,
            I => \A_c_13\
        );

    \I__1106\ : InMux
    port map (
            O => \N__6641\,
            I => \N__6638\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__6638\,
            I => \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\
        );

    \I__1104\ : InMux
    port map (
            O => \N__6635\,
            I => \N__6632\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__6632\,
            I => \U712_CHIP_RAM.N_213\
        );

    \I__1102\ : InMux
    port map (
            O => \N__6629\,
            I => \N__6626\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__6626\,
            I => \N__6623\
        );

    \I__1100\ : Span4Mux_v
    port map (
            O => \N__6623\,
            I => \N__6619\
        );

    \I__1099\ : InMux
    port map (
            O => \N__6622\,
            I => \N__6616\
        );

    \I__1098\ : Odrv4
    port map (
            O => \N__6619\,
            I => \CPU_TACKm\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__6616\,
            I => \CPU_TACKm\
        );

    \I__1096\ : InMux
    port map (
            O => \N__6611\,
            I => \N__6607\
        );

    \I__1095\ : InMux
    port map (
            O => \N__6610\,
            I => \N__6604\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__6607\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__6604\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1092\ : InMux
    port map (
            O => \N__6599\,
            I => \N__6595\
        );

    \I__1091\ : InMux
    port map (
            O => \N__6598\,
            I => \N__6592\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__6595\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__6592\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1088\ : CascadeMux
    port map (
            O => \N__6587\,
            I => \N__6583\
        );

    \I__1087\ : InMux
    port map (
            O => \N__6586\,
            I => \N__6580\
        );

    \I__1086\ : InMux
    port map (
            O => \N__6583\,
            I => \N__6577\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__6580\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__6577\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1083\ : InMux
    port map (
            O => \N__6572\,
            I => \N__6568\
        );

    \I__1082\ : InMux
    port map (
            O => \N__6571\,
            I => \N__6565\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__6568\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__6565\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1079\ : CascadeMux
    port map (
            O => \N__6560\,
            I => \U712_CHIP_RAM.N_333_mux_cascade_\
        );

    \I__1078\ : InMux
    port map (
            O => \N__6557\,
            I => \N__6551\
        );

    \I__1077\ : InMux
    port map (
            O => \N__6556\,
            I => \N__6546\
        );

    \I__1076\ : InMux
    port map (
            O => \N__6555\,
            I => \N__6546\
        );

    \I__1075\ : InMux
    port map (
            O => \N__6554\,
            I => \N__6541\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__6551\,
            I => \N__6538\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__6546\,
            I => \N__6535\
        );

    \I__1072\ : InMux
    port map (
            O => \N__6545\,
            I => \N__6530\
        );

    \I__1071\ : InMux
    port map (
            O => \N__6544\,
            I => \N__6530\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__6541\,
            I => \N__6527\
        );

    \I__1069\ : Odrv12
    port map (
            O => \N__6538\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1068\ : Odrv4
    port map (
            O => \N__6535\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__6530\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1066\ : Odrv4
    port map (
            O => \N__6527\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1065\ : InMux
    port map (
            O => \N__6518\,
            I => \N__6514\
        );

    \I__1064\ : InMux
    port map (
            O => \N__6517\,
            I => \N__6511\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__6514\,
            I => \N__6508\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__6511\,
            I => \U712_CHIP_RAM.N_51_0\
        );

    \I__1061\ : Odrv4
    port map (
            O => \N__6508\,
            I => \U712_CHIP_RAM.N_51_0\
        );

    \I__1060\ : CascadeMux
    port map (
            O => \N__6503\,
            I => \U712_CHIP_RAM.N_51_0_cascade_\
        );

    \I__1059\ : InMux
    port map (
            O => \N__6500\,
            I => \N__6497\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__6497\,
            I => \U712_CHIP_RAM.N_54_0\
        );

    \I__1057\ : InMux
    port map (
            O => \N__6494\,
            I => \N__6491\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__6491\,
            I => \U712_CHIP_RAM.m53_ns_1\
        );

    \I__1055\ : InMux
    port map (
            O => \N__6488\,
            I => \N__6478\
        );

    \I__1054\ : InMux
    port map (
            O => \N__6487\,
            I => \N__6471\
        );

    \I__1053\ : InMux
    port map (
            O => \N__6486\,
            I => \N__6471\
        );

    \I__1052\ : InMux
    port map (
            O => \N__6485\,
            I => \N__6471\
        );

    \I__1051\ : InMux
    port map (
            O => \N__6484\,
            I => \N__6464\
        );

    \I__1050\ : InMux
    port map (
            O => \N__6483\,
            I => \N__6464\
        );

    \I__1049\ : InMux
    port map (
            O => \N__6482\,
            I => \N__6464\
        );

    \I__1048\ : InMux
    port map (
            O => \N__6481\,
            I => \N__6461\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__6478\,
            I => \U712_CHIP_RAM.N_333_mux\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__6471\,
            I => \U712_CHIP_RAM.N_333_mux\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__6464\,
            I => \U712_CHIP_RAM.N_333_mux\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__6461\,
            I => \U712_CHIP_RAM.N_333_mux\
        );

    \I__1043\ : InMux
    port map (
            O => \N__6452\,
            I => \N__6449\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__6449\,
            I => \N__6446\
        );

    \I__1041\ : Odrv4
    port map (
            O => \N__6446\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0\
        );

    \I__1040\ : InMux
    port map (
            O => \N__6443\,
            I => \N__6434\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6442\,
            I => \N__6431\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6441\,
            I => \N__6428\
        );

    \I__1037\ : CascadeMux
    port map (
            O => \N__6440\,
            I => \N__6425\
        );

    \I__1036\ : InMux
    port map (
            O => \N__6439\,
            I => \N__6418\
        );

    \I__1035\ : InMux
    port map (
            O => \N__6438\,
            I => \N__6418\
        );

    \I__1034\ : InMux
    port map (
            O => \N__6437\,
            I => \N__6418\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__6434\,
            I => \N__6415\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__6431\,
            I => \N__6410\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__6428\,
            I => \N__6410\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6425\,
            I => \N__6407\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__6418\,
            I => \N__6399\
        );

    \I__1028\ : Span4Mux_h
    port map (
            O => \N__6415\,
            I => \N__6399\
        );

    \I__1027\ : Span4Mux_v
    port map (
            O => \N__6410\,
            I => \N__6399\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__6407\,
            I => \N__6396\
        );

    \I__1025\ : InMux
    port map (
            O => \N__6406\,
            I => \N__6393\
        );

    \I__1024\ : Odrv4
    port map (
            O => \N__6399\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1023\ : Odrv4
    port map (
            O => \N__6396\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__6393\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1021\ : InMux
    port map (
            O => \N__6386\,
            I => \N__6380\
        );

    \I__1020\ : InMux
    port map (
            O => \N__6385\,
            I => \N__6380\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__6380\,
            I => \N__6377\
        );

    \I__1018\ : Odrv4
    port map (
            O => \N__6377\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__6374\,
            I => \N__6371\
        );

    \I__1016\ : InMux
    port map (
            O => \N__6371\,
            I => \N__6368\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__6368\,
            I => \N__6364\
        );

    \I__1014\ : InMux
    port map (
            O => \N__6367\,
            I => \N__6361\
        );

    \I__1013\ : Odrv4
    port map (
            O => \N__6364\,
            I => \U712_CHIP_RAM.m41_1\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__6361\,
            I => \U712_CHIP_RAM.m41_1\
        );

    \I__1011\ : CascadeMux
    port map (
            O => \N__6356\,
            I => \U712_CHIP_RAM.N_31_0_cascade_\
        );

    \I__1010\ : CascadeMux
    port map (
            O => \N__6353\,
            I => \U712_CHIP_RAM.m217_ns_1_cascade_\
        );

    \I__1009\ : InMux
    port map (
            O => \N__6350\,
            I => \N__6347\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__6347\,
            I => \U712_CHIP_RAM.N_218\
        );

    \I__1007\ : CascadeMux
    port map (
            O => \N__6344\,
            I => \U712_CHIP_RAM.m212_ns_1_cascade_\
        );

    \I__1006\ : CascadeMux
    port map (
            O => \N__6341\,
            I => \U712_CHIP_RAM.N_30_0_cascade_\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6338\,
            I => \N__6335\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__6335\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_2\
        );

    \I__1003\ : InMux
    port map (
            O => \N__6332\,
            I => \N__6329\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__6329\,
            I => \N__6326\
        );

    \I__1001\ : Sp12to4
    port map (
            O => \N__6326\,
            I => \N__6323\
        );

    \I__1000\ : Span12Mux_v
    port map (
            O => \N__6323\,
            I => \N__6320\
        );

    \I__999\ : Span12Mux_h
    port map (
            O => \N__6320\,
            I => \N__6317\
        );

    \I__998\ : Odrv12
    port map (
            O => \N__6317\,
            I => \A_c_2\
        );

    \I__997\ : InMux
    port map (
            O => \N__6314\,
            I => \N__6310\
        );

    \I__996\ : InMux
    port map (
            O => \N__6313\,
            I => \N__6307\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__6310\,
            I => \N__6304\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__6307\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\
        );

    \I__993\ : Odrv4
    port map (
            O => \N__6304\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\
        );

    \I__992\ : InMux
    port map (
            O => \N__6299\,
            I => \N__6296\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__6296\,
            I => \N__6293\
        );

    \I__990\ : Span4Mux_v
    port map (
            O => \N__6293\,
            I => \N__6290\
        );

    \I__989\ : Span4Mux_v
    port map (
            O => \N__6290\,
            I => \N__6287\
        );

    \I__988\ : Sp12to4
    port map (
            O => \N__6287\,
            I => \N__6284\
        );

    \I__987\ : Span12Mux_h
    port map (
            O => \N__6284\,
            I => \N__6281\
        );

    \I__986\ : Odrv12
    port map (
            O => \N__6281\,
            I => \A_c_20\
        );

    \I__985\ : InMux
    port map (
            O => \N__6278\,
            I => \N__6274\
        );

    \I__984\ : InMux
    port map (
            O => \N__6277\,
            I => \N__6271\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__6274\,
            I => \N__6268\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__6271\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\
        );

    \I__981\ : Odrv4
    port map (
            O => \N__6268\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\
        );

    \I__980\ : InMux
    port map (
            O => \N__6263\,
            I => \N__6259\
        );

    \I__979\ : InMux
    port map (
            O => \N__6262\,
            I => \N__6256\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__6259\,
            I => \N__6251\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__6256\,
            I => \N__6251\
        );

    \I__976\ : Odrv4
    port map (
            O => \N__6251\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__975\ : InMux
    port map (
            O => \N__6248\,
            I => \N__6244\
        );

    \I__974\ : InMux
    port map (
            O => \N__6247\,
            I => \N__6241\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__6244\,
            I => \N__6238\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__6241\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__971\ : Odrv4
    port map (
            O => \N__6238\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__970\ : CascadeMux
    port map (
            O => \N__6233\,
            I => \N__6229\
        );

    \I__969\ : InMux
    port map (
            O => \N__6232\,
            I => \N__6226\
        );

    \I__968\ : InMux
    port map (
            O => \N__6229\,
            I => \N__6223\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__6226\,
            I => \N__6218\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__6223\,
            I => \N__6218\
        );

    \I__965\ : Odrv4
    port map (
            O => \N__6218\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__964\ : InMux
    port map (
            O => \N__6215\,
            I => \N__6212\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__6212\,
            I => \N__6209\
        );

    \I__962\ : Odrv4
    port map (
            O => \N__6209\,
            I => \U712_CHIP_RAM.REFRESH5lt7\
        );

    \I__961\ : InMux
    port map (
            O => \N__6206\,
            I => \N__6203\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__6203\,
            I => \N__6198\
        );

    \I__959\ : InMux
    port map (
            O => \N__6202\,
            I => \N__6195\
        );

    \I__958\ : InMux
    port map (
            O => \N__6201\,
            I => \N__6192\
        );

    \I__957\ : Odrv4
    port map (
            O => \N__6198\,
            I => \U712_CHIP_RAM.N_28_0\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__6195\,
            I => \U712_CHIP_RAM.N_28_0\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__6192\,
            I => \U712_CHIP_RAM.N_28_0\
        );

    \I__954\ : InMux
    port map (
            O => \N__6185\,
            I => \N__6182\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__6182\,
            I => \U712_CHIP_RAM.N_219\
        );

    \I__952\ : InMux
    port map (
            O => \N__6179\,
            I => \N__6176\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__6176\,
            I => \U712_CHIP_RAM.d_N_6_5\
        );

    \I__950\ : InMux
    port map (
            O => \N__6173\,
            I => \N__6170\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__6170\,
            I => \U712_CHIP_RAM.d_N_6_1\
        );

    \I__948\ : InMux
    port map (
            O => \N__6167\,
            I => \N__6164\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__6164\,
            I => \N__6161\
        );

    \I__946\ : Odrv4
    port map (
            O => \N__6161\,
            I => \U712_CHIP_RAM.N_353_mux\
        );

    \I__945\ : CascadeMux
    port map (
            O => \N__6158\,
            I => \U712_CHIP_RAM.N_168_0_cascade_\
        );

    \I__944\ : InMux
    port map (
            O => \N__6155\,
            I => \N__6152\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__6152\,
            I => \U712_CHIP_RAM.m64_ns_1\
        );

    \I__942\ : CascadeMux
    port map (
            O => \N__6149\,
            I => \U712_CHIP_RAM.i67_mux_cascade_\
        );

    \I__941\ : InMux
    port map (
            O => \N__6146\,
            I => \N__6143\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__6143\,
            I => \N__6140\
        );

    \I__939\ : Odrv4
    port map (
            O => \N__6140\,
            I => \U712_CHIP_RAM.m66_ns_1\
        );

    \I__938\ : InMux
    port map (
            O => \N__6137\,
            I => \N__6134\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__6134\,
            I => \U712_CHIP_RAM.N_146_0\
        );

    \I__936\ : CascadeMux
    port map (
            O => \N__6131\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_2_cascade_\
        );

    \I__935\ : CascadeMux
    port map (
            O => \N__6128\,
            I => \U712_CHIP_RAM.N_151_0_cascade_\
        );

    \I__934\ : CascadeMux
    port map (
            O => \N__6125\,
            I => \N__6122\
        );

    \I__933\ : InMux
    port map (
            O => \N__6122\,
            I => \N__6117\
        );

    \I__932\ : InMux
    port map (
            O => \N__6121\,
            I => \N__6112\
        );

    \I__931\ : InMux
    port map (
            O => \N__6120\,
            I => \N__6112\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__6117\,
            I => \N__6107\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__6112\,
            I => \N__6107\
        );

    \I__928\ : Odrv4
    port map (
            O => \N__6107\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\
        );

    \I__927\ : InMux
    port map (
            O => \N__6104\,
            I => \N__6101\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__6101\,
            I => \U712_REG_SM_UDSn_6_0\
        );

    \I__925\ : IoInMux
    port map (
            O => \N__6098\,
            I => \N__6095\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__6095\,
            I => \N__6092\
        );

    \I__923\ : Span4Mux_s3_v
    port map (
            O => \N__6092\,
            I => \N__6089\
        );

    \I__922\ : Span4Mux_v
    port map (
            O => \N__6089\,
            I => \N__6086\
        );

    \I__921\ : Span4Mux_v
    port map (
            O => \N__6086\,
            I => \N__6083\
        );

    \I__920\ : Sp12to4
    port map (
            O => \N__6083\,
            I => \N__6079\
        );

    \I__919\ : InMux
    port map (
            O => \N__6082\,
            I => \N__6076\
        );

    \I__918\ : Odrv12
    port map (
            O => \N__6079\,
            I => \UDSn_c\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__6076\,
            I => \UDSn_c\
        );

    \I__916\ : InMux
    port map (
            O => \N__6071\,
            I => \N__6068\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__6068\,
            I => \N__6065\
        );

    \I__914\ : Span4Mux_v
    port map (
            O => \N__6065\,
            I => \N__6061\
        );

    \I__913\ : InMux
    port map (
            O => \N__6064\,
            I => \N__6058\
        );

    \I__912\ : Span4Mux_v
    port map (
            O => \N__6061\,
            I => \N__6055\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__6058\,
            I => \N__6052\
        );

    \I__910\ : Sp12to4
    port map (
            O => \N__6055\,
            I => \N__6049\
        );

    \I__909\ : Span4Mux_h
    port map (
            O => \N__6052\,
            I => \N__6046\
        );

    \I__908\ : Odrv12
    port map (
            O => \N__6049\,
            I => \DBRn_c_i\
        );

    \I__907\ : Odrv4
    port map (
            O => \N__6046\,
            I => \DBRn_c_i\
        );

    \I__906\ : IoInMux
    port map (
            O => \N__6041\,
            I => \N__6038\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__6038\,
            I => \N__6035\
        );

    \I__904\ : IoSpan4Mux
    port map (
            O => \N__6035\,
            I => \N__6032\
        );

    \I__903\ : Span4Mux_s3_h
    port map (
            O => \N__6032\,
            I => \N__6029\
        );

    \I__902\ : Sp12to4
    port map (
            O => \N__6029\,
            I => \N__6026\
        );

    \I__901\ : Span12Mux_h
    port map (
            O => \N__6026\,
            I => \N__6023\
        );

    \I__900\ : Odrv12
    port map (
            O => \N__6023\,
            I => \CMA_c_8\
        );

    \I__899\ : IoInMux
    port map (
            O => \N__6020\,
            I => \N__6016\
        );

    \I__898\ : InMux
    port map (
            O => \N__6019\,
            I => \N__6013\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__6016\,
            I => \N__6010\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__6013\,
            I => \N__6007\
        );

    \I__895\ : Span12Mux_s4_v
    port map (
            O => \N__6010\,
            I => \N__6004\
        );

    \I__894\ : Span4Mux_v
    port map (
            O => \N__6007\,
            I => \N__6001\
        );

    \I__893\ : Span12Mux_v
    port map (
            O => \N__6004\,
            I => \N__5998\
        );

    \I__892\ : Span4Mux_h
    port map (
            O => \N__6001\,
            I => \N__5995\
        );

    \I__891\ : Span12Mux_h
    port map (
            O => \N__5998\,
            I => \N__5992\
        );

    \I__890\ : Sp12to4
    port map (
            O => \N__5995\,
            I => \N__5989\
        );

    \I__889\ : Odrv12
    port map (
            O => \N__5992\,
            I => \A_c_9\
        );

    \I__888\ : Odrv12
    port map (
            O => \N__5989\,
            I => \A_c_9\
        );

    \I__887\ : CascadeMux
    port map (
            O => \N__5984\,
            I => \U712_CHIP_RAM.m186_0_cascade_\
        );

    \I__886\ : InMux
    port map (
            O => \N__5981\,
            I => \N__5978\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5978\,
            I => \N__5975\
        );

    \I__884\ : Sp12to4
    port map (
            O => \N__5975\,
            I => \N__5972\
        );

    \I__883\ : Span12Mux_v
    port map (
            O => \N__5972\,
            I => \N__5969\
        );

    \I__882\ : Span12Mux_h
    port map (
            O => \N__5969\,
            I => \N__5966\
        );

    \I__881\ : Odrv12
    port map (
            O => \N__5966\,
            I => \A_c_17\
        );

    \I__880\ : CascadeMux
    port map (
            O => \N__5963\,
            I => \U712_CHIP_RAM.m192_0_cascade_\
        );

    \I__879\ : InMux
    port map (
            O => \N__5960\,
            I => \N__5956\
        );

    \I__878\ : InMux
    port map (
            O => \N__5959\,
            I => \N__5953\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__5956\,
            I => \N__5950\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__5953\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__875\ : Odrv4
    port map (
            O => \N__5950\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__874\ : InMux
    port map (
            O => \N__5945\,
            I => \N__5942\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__5942\,
            I => \U712_CHIP_RAM.m192_1\
        );

    \I__872\ : CascadeMux
    port map (
            O => \N__5939\,
            I => \N__5936\
        );

    \I__871\ : InMux
    port map (
            O => \N__5936\,
            I => \N__5933\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__5933\,
            I => \N__5930\
        );

    \I__869\ : Odrv4
    port map (
            O => \N__5930\,
            I => \U712_CHIP_RAM.N_215\
        );

    \I__868\ : InMux
    port map (
            O => \N__5927\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__867\ : InMux
    port map (
            O => \N__5924\,
            I => \N__5921\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__5921\,
            I => \N__5918\
        );

    \I__865\ : Odrv4
    port map (
            O => \N__5918\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__864\ : InMux
    port map (
            O => \N__5915\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__863\ : InMux
    port map (
            O => \N__5912\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__862\ : InMux
    port map (
            O => \N__5909\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__861\ : InMux
    port map (
            O => \N__5906\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__860\ : InMux
    port map (
            O => \N__5903\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__859\ : CascadeMux
    port map (
            O => \N__5900\,
            I => \N__5897\
        );

    \I__858\ : InMux
    port map (
            O => \N__5897\,
            I => \N__5894\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__5894\,
            I => \N__5884\
        );

    \I__856\ : InMux
    port map (
            O => \N__5893\,
            I => \N__5881\
        );

    \I__855\ : InMux
    port map (
            O => \N__5892\,
            I => \N__5872\
        );

    \I__854\ : InMux
    port map (
            O => \N__5891\,
            I => \N__5872\
        );

    \I__853\ : InMux
    port map (
            O => \N__5890\,
            I => \N__5872\
        );

    \I__852\ : InMux
    port map (
            O => \N__5889\,
            I => \N__5872\
        );

    \I__851\ : InMux
    port map (
            O => \N__5888\,
            I => \N__5867\
        );

    \I__850\ : InMux
    port map (
            O => \N__5887\,
            I => \N__5867\
        );

    \I__849\ : Odrv4
    port map (
            O => \N__5884\,
            I => \U712_CHIP_RAM.N_56_0_i\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__5881\,
            I => \U712_CHIP_RAM.N_56_0_i\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__5872\,
            I => \U712_CHIP_RAM.N_56_0_i\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__5867\,
            I => \U712_CHIP_RAM.N_56_0_i\
        );

    \I__845\ : InMux
    port map (
            O => \N__5858\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__844\ : CEMux
    port map (
            O => \N__5855\,
            I => \N__5851\
        );

    \I__843\ : CEMux
    port map (
            O => \N__5854\,
            I => \N__5847\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__5851\,
            I => \N__5844\
        );

    \I__841\ : CEMux
    port map (
            O => \N__5850\,
            I => \N__5841\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__5847\,
            I => \N__5838\
        );

    \I__839\ : Span4Mux_v
    port map (
            O => \N__5844\,
            I => \N__5835\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__5841\,
            I => \N__5832\
        );

    \I__837\ : Odrv4
    port map (
            O => \N__5838\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__836\ : Odrv4
    port map (
            O => \N__5835\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__835\ : Odrv4
    port map (
            O => \N__5832\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__834\ : InMux
    port map (
            O => \N__5825\,
            I => \N__5822\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__5822\,
            I => \U712_CHIP_RAM.N_330\
        );

    \I__832\ : InMux
    port map (
            O => \N__5819\,
            I => \N__5816\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__5816\,
            I => \N__5813\
        );

    \I__830\ : Odrv4
    port map (
            O => \N__5813\,
            I => \U712_CHIP_RAM.m38_1\
        );

    \I__829\ : CascadeMux
    port map (
            O => \N__5810\,
            I => \U712_CHIP_RAM.N_34_0_cascade_\
        );

    \I__828\ : CascadeMux
    port map (
            O => \N__5807\,
            I => \N__5804\
        );

    \I__827\ : InMux
    port map (
            O => \N__5804\,
            I => \N__5801\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__5801\,
            I => \U712_CHIP_RAM.N_359\
        );

    \I__825\ : InMux
    port map (
            O => \N__5798\,
            I => \N__5792\
        );

    \I__824\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5785\
        );

    \I__823\ : InMux
    port map (
            O => \N__5796\,
            I => \N__5785\
        );

    \I__822\ : InMux
    port map (
            O => \N__5795\,
            I => \N__5785\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__5792\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__5785\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__819\ : InMux
    port map (
            O => \N__5780\,
            I => \N__5776\
        );

    \I__818\ : InMux
    port map (
            O => \N__5779\,
            I => \N__5773\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__5776\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__5773\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__815\ : CascadeMux
    port map (
            O => \N__5768\,
            I => \U712_CHIP_RAM.N_28_0_cascade_\
        );

    \I__814\ : CascadeMux
    port map (
            O => \N__5765\,
            I => \U712_CHIP_RAM.N_47_0_cascade_\
        );

    \I__813\ : CascadeMux
    port map (
            O => \N__5762\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_cascade_\
        );

    \I__812\ : CEMux
    port map (
            O => \N__5759\,
            I => \N__5756\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__5756\,
            I => \N__5753\
        );

    \I__810\ : Span4Mux_v
    port map (
            O => \N__5753\,
            I => \N__5750\
        );

    \I__809\ : Odrv4
    port map (
            O => \N__5750\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0\
        );

    \I__808\ : CascadeMux
    port map (
            O => \N__5747\,
            I => \U712_CHIP_RAM.N_146_0_cascade_\
        );

    \I__807\ : CascadeMux
    port map (
            O => \N__5744\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_3_cascade_\
        );

    \I__806\ : InMux
    port map (
            O => \N__5741\,
            I => \N__5738\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__5738\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_3\
        );

    \I__804\ : CascadeMux
    port map (
            O => \N__5735\,
            I => \U712_CHIP_RAM.N_154_0_cascade_\
        );

    \I__803\ : InMux
    port map (
            O => \N__5732\,
            I => \N__5729\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__5729\,
            I => \N__5726\
        );

    \I__801\ : Odrv4
    port map (
            O => \N__5726\,
            I => \U712_CHIP_RAM.N_7_0\
        );

    \I__800\ : InMux
    port map (
            O => \N__5723\,
            I => \N__5719\
        );

    \I__799\ : InMux
    port map (
            O => \N__5722\,
            I => \N__5716\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__5719\,
            I => \N_86_0\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5716\,
            I => \N_86_0\
        );

    \I__796\ : CascadeMux
    port map (
            O => \N__5711\,
            I => \N__5706\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__5710\,
            I => \N__5702\
        );

    \I__794\ : InMux
    port map (
            O => \N__5709\,
            I => \N__5696\
        );

    \I__793\ : InMux
    port map (
            O => \N__5706\,
            I => \N__5693\
        );

    \I__792\ : InMux
    port map (
            O => \N__5705\,
            I => \N__5690\
        );

    \I__791\ : InMux
    port map (
            O => \N__5702\,
            I => \N__5687\
        );

    \I__790\ : CascadeMux
    port map (
            O => \N__5701\,
            I => \N__5684\
        );

    \I__789\ : InMux
    port map (
            O => \N__5700\,
            I => \N__5678\
        );

    \I__788\ : InMux
    port map (
            O => \N__5699\,
            I => \N__5675\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5696\,
            I => \N__5668\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__5693\,
            I => \N__5668\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__5690\,
            I => \N__5668\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__5687\,
            I => \N__5662\
        );

    \I__783\ : InMux
    port map (
            O => \N__5684\,
            I => \N__5659\
        );

    \I__782\ : InMux
    port map (
            O => \N__5683\,
            I => \N__5656\
        );

    \I__781\ : InMux
    port map (
            O => \N__5682\,
            I => \N__5651\
        );

    \I__780\ : InMux
    port map (
            O => \N__5681\,
            I => \N__5651\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__5678\,
            I => \N__5646\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__5675\,
            I => \N__5646\
        );

    \I__777\ : Span4Mux_v
    port map (
            O => \N__5668\,
            I => \N__5643\
        );

    \I__776\ : InMux
    port map (
            O => \N__5667\,
            I => \N__5636\
        );

    \I__775\ : InMux
    port map (
            O => \N__5666\,
            I => \N__5636\
        );

    \I__774\ : InMux
    port map (
            O => \N__5665\,
            I => \N__5636\
        );

    \I__773\ : Span4Mux_h
    port map (
            O => \N__5662\,
            I => \N__5633\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__5659\,
            I => \U712_REG_SM_C3_SYNC_1\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__5656\,
            I => \U712_REG_SM_C3_SYNC_1\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__5651\,
            I => \U712_REG_SM_C3_SYNC_1\
        );

    \I__769\ : Odrv4
    port map (
            O => \N__5646\,
            I => \U712_REG_SM_C3_SYNC_1\
        );

    \I__768\ : Odrv4
    port map (
            O => \N__5643\,
            I => \U712_REG_SM_C3_SYNC_1\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__5636\,
            I => \U712_REG_SM_C3_SYNC_1\
        );

    \I__766\ : Odrv4
    port map (
            O => \N__5633\,
            I => \U712_REG_SM_C3_SYNC_1\
        );

    \I__765\ : IoInMux
    port map (
            O => \N__5618\,
            I => \N__5615\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__5615\,
            I => \N__5611\
        );

    \I__763\ : IoInMux
    port map (
            O => \N__5614\,
            I => \N__5608\
        );

    \I__762\ : IoSpan4Mux
    port map (
            O => \N__5611\,
            I => \N__5605\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__5608\,
            I => \N__5602\
        );

    \I__760\ : Sp12to4
    port map (
            O => \N__5605\,
            I => \N__5599\
        );

    \I__759\ : Span4Mux_s1_v
    port map (
            O => \N__5602\,
            I => \N__5596\
        );

    \I__758\ : Span12Mux_s7_h
    port map (
            O => \N__5599\,
            I => \N__5593\
        );

    \I__757\ : Sp12to4
    port map (
            O => \N__5596\,
            I => \N__5590\
        );

    \I__756\ : Span12Mux_h
    port map (
            O => \N__5593\,
            I => \N__5585\
        );

    \I__755\ : Span12Mux_h
    port map (
            O => \N__5590\,
            I => \N__5585\
        );

    \I__754\ : Odrv12
    port map (
            O => \N__5585\,
            I => \BLSn_c\
        );

    \I__753\ : CEMux
    port map (
            O => \N__5582\,
            I => \N__5579\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__5579\,
            I => \N__5576\
        );

    \I__751\ : Span4Mux_v
    port map (
            O => \N__5576\,
            I => \N__5573\
        );

    \I__750\ : Span4Mux_h
    port map (
            O => \N__5573\,
            I => \N__5570\
        );

    \I__749\ : Odrv4
    port map (
            O => \N__5570\,
            I => \U712_REG_SM.N_86_0_0\
        );

    \I__748\ : CascadeMux
    port map (
            O => \N__5567\,
            I => \U712_CYCLE_TERM.N_36_0_cascade_\
        );

    \I__747\ : IoInMux
    port map (
            O => \N__5564\,
            I => \N__5559\
        );

    \I__746\ : IoInMux
    port map (
            O => \N__5563\,
            I => \N__5556\
        );

    \I__745\ : IoInMux
    port map (
            O => \N__5562\,
            I => \N__5553\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__5559\,
            I => \N__5550\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__5556\,
            I => \N__5547\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__5553\,
            I => \N__5544\
        );

    \I__741\ : Span4Mux_s1_h
    port map (
            O => \N__5550\,
            I => \N__5541\
        );

    \I__740\ : Span4Mux_s0_v
    port map (
            O => \N__5547\,
            I => \N__5538\
        );

    \I__739\ : Span4Mux_s3_v
    port map (
            O => \N__5544\,
            I => \N__5535\
        );

    \I__738\ : Sp12to4
    port map (
            O => \N__5541\,
            I => \N__5532\
        );

    \I__737\ : Span4Mux_h
    port map (
            O => \N__5538\,
            I => \N__5529\
        );

    \I__736\ : Span4Mux_v
    port map (
            O => \N__5535\,
            I => \N__5526\
        );

    \I__735\ : Span12Mux_s11_v
    port map (
            O => \N__5532\,
            I => \N__5523\
        );

    \I__734\ : Sp12to4
    port map (
            O => \N__5529\,
            I => \N__5520\
        );

    \I__733\ : Span4Mux_h
    port map (
            O => \N__5526\,
            I => \N__5517\
        );

    \I__732\ : Span12Mux_h
    port map (
            O => \N__5523\,
            I => \N__5513\
        );

    \I__731\ : Span12Mux_h
    port map (
            O => \N__5520\,
            I => \N__5510\
        );

    \I__730\ : Span4Mux_h
    port map (
            O => \N__5517\,
            I => \N__5507\
        );

    \I__729\ : InMux
    port map (
            O => \N__5516\,
            I => \N__5504\
        );

    \I__728\ : Odrv12
    port map (
            O => \N__5513\,
            I => \TACK_OUT\
        );

    \I__727\ : Odrv12
    port map (
            O => \N__5510\,
            I => \TACK_OUT\
        );

    \I__726\ : Odrv4
    port map (
            O => \N__5507\,
            I => \TACK_OUT\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__5504\,
            I => \TACK_OUT\
        );

    \I__724\ : InMux
    port map (
            O => \N__5495\,
            I => \N__5490\
        );

    \I__723\ : InMux
    port map (
            O => \N__5494\,
            I => \N__5485\
        );

    \I__722\ : InMux
    port map (
            O => \N__5493\,
            I => \N__5485\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__5490\,
            I => \N__5480\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__5485\,
            I => \N__5480\
        );

    \I__719\ : Span4Mux_h
    port map (
            O => \N__5480\,
            I => \N__5476\
        );

    \I__718\ : InMux
    port map (
            O => \N__5479\,
            I => \N__5473\
        );

    \I__717\ : Span4Mux_v
    port map (
            O => \N__5476\,
            I => \N__5470\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__5473\,
            I => \U712_CYCLE_TERM.TACK_STARTZ0\
        );

    \I__715\ : Odrv4
    port map (
            O => \N__5470\,
            I => \U712_CYCLE_TERM.TACK_STARTZ0\
        );

    \I__714\ : InMux
    port map (
            O => \N__5465\,
            I => \N__5458\
        );

    \I__713\ : InMux
    port map (
            O => \N__5464\,
            I => \N__5449\
        );

    \I__712\ : InMux
    port map (
            O => \N__5463\,
            I => \N__5449\
        );

    \I__711\ : InMux
    port map (
            O => \N__5462\,
            I => \N__5449\
        );

    \I__710\ : InMux
    port map (
            O => \N__5461\,
            I => \N__5449\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__5458\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__5449\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__707\ : CascadeMux
    port map (
            O => \N__5444\,
            I => \N__5441\
        );

    \I__706\ : InMux
    port map (
            O => \N__5441\,
            I => \N__5436\
        );

    \I__705\ : InMux
    port map (
            O => \N__5440\,
            I => \N__5431\
        );

    \I__704\ : InMux
    port map (
            O => \N__5439\,
            I => \N__5431\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__5436\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__5431\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__701\ : InMux
    port map (
            O => \N__5426\,
            I => \N__5423\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__5423\,
            I => \U712_CHIP_RAM.N_83_0\
        );

    \I__699\ : CascadeMux
    port map (
            O => \N__5420\,
            I => \U712_CHIP_RAM.N_94_0_cascade_\
        );

    \I__698\ : InMux
    port map (
            O => \N__5417\,
            I => \N__5412\
        );

    \I__697\ : InMux
    port map (
            O => \N__5416\,
            I => \N__5405\
        );

    \I__696\ : InMux
    port map (
            O => \N__5415\,
            I => \N__5405\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__5412\,
            I => \N__5402\
        );

    \I__694\ : InMux
    port map (
            O => \N__5411\,
            I => \N__5399\
        );

    \I__693\ : InMux
    port map (
            O => \N__5410\,
            I => \N__5396\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__5405\,
            I => \U712_REG_SM_STATE_COUNT_1\
        );

    \I__691\ : Odrv4
    port map (
            O => \N__5402\,
            I => \U712_REG_SM_STATE_COUNT_1\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__5399\,
            I => \U712_REG_SM_STATE_COUNT_1\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__5396\,
            I => \U712_REG_SM_STATE_COUNT_1\
        );

    \I__688\ : InMux
    port map (
            O => \N__5387\,
            I => \N__5383\
        );

    \I__687\ : InMux
    port map (
            O => \N__5386\,
            I => \N__5380\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__5383\,
            I => \U712_REG_SM_STATE_COUNT_2\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__5380\,
            I => \U712_REG_SM_STATE_COUNT_2\
        );

    \I__684\ : InMux
    port map (
            O => \N__5375\,
            I => \N__5371\
        );

    \I__683\ : CascadeMux
    port map (
            O => \N__5374\,
            I => \N__5368\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__5371\,
            I => \N__5365\
        );

    \I__681\ : InMux
    port map (
            O => \N__5368\,
            I => \N__5362\
        );

    \I__680\ : Odrv4
    port map (
            O => \N__5365\,
            I => \DBR_SYNC_i_1\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__5362\,
            I => \DBR_SYNC_i_1\
        );

    \I__678\ : InMux
    port map (
            O => \N__5357\,
            I => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\
        );

    \I__677\ : InMux
    port map (
            O => \N__5354\,
            I => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\
        );

    \I__676\ : InMux
    port map (
            O => \N__5351\,
            I => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2\
        );

    \I__675\ : InMux
    port map (
            O => \N__5348\,
            I => \N__5345\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__5345\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1\
        );

    \I__673\ : CascadeMux
    port map (
            O => \N__5342\,
            I => \N__5339\
        );

    \I__672\ : InMux
    port map (
            O => \N__5339\,
            I => \N__5336\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__5336\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2\
        );

    \I__670\ : InMux
    port map (
            O => \N__5333\,
            I => \N__5327\
        );

    \I__669\ : InMux
    port map (
            O => \N__5332\,
            I => \N__5327\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__5327\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\
        );

    \I__667\ : CascadeMux
    port map (
            O => \N__5324\,
            I => \N__5321\
        );

    \I__666\ : InMux
    port map (
            O => \N__5321\,
            I => \N__5315\
        );

    \I__665\ : InMux
    port map (
            O => \N__5320\,
            I => \N__5315\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__5315\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_1\
        );

    \I__663\ : CascadeMux
    port map (
            O => \N__5312\,
            I => \N__5309\
        );

    \I__662\ : InMux
    port map (
            O => \N__5309\,
            I => \N__5306\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__5306\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3\
        );

    \I__660\ : InMux
    port map (
            O => \N__5303\,
            I => \N__5297\
        );

    \I__659\ : InMux
    port map (
            O => \N__5302\,
            I => \N__5297\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__5297\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\
        );

    \I__657\ : InMux
    port map (
            O => \N__5294\,
            I => \N__5290\
        );

    \I__656\ : IoInMux
    port map (
            O => \N__5293\,
            I => \N__5287\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__5290\,
            I => \N__5284\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__5287\,
            I => \N__5281\
        );

    \I__653\ : Span4Mux_v
    port map (
            O => \N__5284\,
            I => \N__5278\
        );

    \I__652\ : IoSpan4Mux
    port map (
            O => \N__5281\,
            I => \N__5275\
        );

    \I__651\ : Sp12to4
    port map (
            O => \N__5278\,
            I => \N__5272\
        );

    \I__650\ : IoSpan4Mux
    port map (
            O => \N__5275\,
            I => \N__5269\
        );

    \I__649\ : Span12Mux_h
    port map (
            O => \N__5272\,
            I => \N__5266\
        );

    \I__648\ : IoSpan4Mux
    port map (
            O => \N__5269\,
            I => \N__5263\
        );

    \I__647\ : Odrv12
    port map (
            O => \N__5266\,
            I => \C1_c\
        );

    \I__646\ : Odrv4
    port map (
            O => \N__5263\,
            I => \C1_c\
        );

    \I__645\ : InMux
    port map (
            O => \N__5258\,
            I => \N__5255\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__5255\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__643\ : InMux
    port map (
            O => \N__5252\,
            I => \N__5249\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__5249\,
            I => \U712_CHIP_RAM.m231_0\
        );

    \I__641\ : InMux
    port map (
            O => \N__5246\,
            I => \N__5243\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__5243\,
            I => \U712_CHIP_RAM.N_236\
        );

    \I__639\ : InMux
    port map (
            O => \N__5240\,
            I => \N__5235\
        );

    \I__638\ : InMux
    port map (
            O => \N__5239\,
            I => \N__5232\
        );

    \I__637\ : InMux
    port map (
            O => \N__5238\,
            I => \N__5229\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__5235\,
            I => \N__5224\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__5232\,
            I => \N__5224\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__5229\,
            I => \U712_REG_SM_STATE_COUNT_0_sqmuxa_1\
        );

    \I__633\ : Odrv4
    port map (
            O => \N__5224\,
            I => \U712_REG_SM_STATE_COUNT_0_sqmuxa_1\
        );

    \I__632\ : CascadeMux
    port map (
            O => \N__5219\,
            I => \U712_CHIP_RAM.N_83_0_cascade_\
        );

    \I__631\ : CascadeMux
    port map (
            O => \N__5216\,
            I => \N__5212\
        );

    \I__630\ : CascadeMux
    port map (
            O => \N__5215\,
            I => \N__5209\
        );

    \I__629\ : InMux
    port map (
            O => \N__5212\,
            I => \N__5204\
        );

    \I__628\ : InMux
    port map (
            O => \N__5209\,
            I => \N__5201\
        );

    \I__627\ : InMux
    port map (
            O => \N__5208\,
            I => \N__5196\
        );

    \I__626\ : InMux
    port map (
            O => \N__5207\,
            I => \N__5196\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__5204\,
            I => \U712_REG_SM_REG_CYCLE_START\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__5201\,
            I => \U712_REG_SM_REG_CYCLE_START\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__5196\,
            I => \U712_REG_SM_REG_CYCLE_START\
        );

    \I__622\ : InMux
    port map (
            O => \N__5189\,
            I => \N__5183\
        );

    \I__621\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5183\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__5183\,
            I => \U712_REG_SM_START_RST\
        );

    \I__619\ : InMux
    port map (
            O => \N__5180\,
            I => \N__5177\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__5177\,
            I => \N__5174\
        );

    \I__617\ : Odrv4
    port map (
            O => \N__5174\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_3\
        );

    \I__616\ : InMux
    port map (
            O => \N__5171\,
            I => \N__5168\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__5168\,
            I => \N__5165\
        );

    \I__614\ : Span4Mux_h
    port map (
            O => \N__5165\,
            I => \N__5162\
        );

    \I__613\ : Span4Mux_v
    port map (
            O => \N__5162\,
            I => \N__5158\
        );

    \I__612\ : IoInMux
    port map (
            O => \N__5161\,
            I => \N__5155\
        );

    \I__611\ : Span4Mux_v
    port map (
            O => \N__5158\,
            I => \N__5152\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__5155\,
            I => \N__5149\
        );

    \I__609\ : Span4Mux_v
    port map (
            O => \N__5152\,
            I => \N__5146\
        );

    \I__608\ : IoSpan4Mux
    port map (
            O => \N__5149\,
            I => \N__5143\
        );

    \I__607\ : Odrv4
    port map (
            O => \N__5146\,
            I => \RAMENn_c\
        );

    \I__606\ : Odrv4
    port map (
            O => \N__5143\,
            I => \RAMENn_c\
        );

    \I__605\ : CascadeMux
    port map (
            O => \N__5138\,
            I => \N__5134\
        );

    \I__604\ : InMux
    port map (
            O => \N__5137\,
            I => \N__5129\
        );

    \I__603\ : InMux
    port map (
            O => \N__5134\,
            I => \N__5129\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__5129\,
            I => \N__5126\
        );

    \I__601\ : Span4Mux_v
    port map (
            O => \N__5126\,
            I => \N__5123\
        );

    \I__600\ : Sp12to4
    port map (
            O => \N__5123\,
            I => \N__5120\
        );

    \I__599\ : Span12Mux_h
    port map (
            O => \N__5120\,
            I => \N__5117\
        );

    \I__598\ : Span12Mux_v
    port map (
            O => \N__5117\,
            I => \N__5114\
        );

    \I__597\ : Odrv12
    port map (
            O => \N__5114\,
            I => \TSn_c\
        );

    \I__596\ : CascadeMux
    port map (
            O => \N__5111\,
            I => \U712_CHIP_RAM.m223_ns_1_cascade_\
        );

    \I__595\ : InMux
    port map (
            O => \N__5108\,
            I => \N__5105\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__5105\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_5\
        );

    \I__593\ : InMux
    port map (
            O => \N__5102\,
            I => \N__5098\
        );

    \I__592\ : InMux
    port map (
            O => \N__5101\,
            I => \N__5095\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__5098\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__5095\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\
        );

    \I__589\ : InMux
    port map (
            O => \N__5090\,
            I => \N__5087\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__5087\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__587\ : InMux
    port map (
            O => \N__5084\,
            I => \bfn_9_11_0_\
        );

    \I__586\ : InMux
    port map (
            O => \N__5081\,
            I => \N__5077\
        );

    \I__585\ : InMux
    port map (
            O => \N__5080\,
            I => \N__5074\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__5077\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__5074\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__582\ : InMux
    port map (
            O => \N__5069\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__581\ : InMux
    port map (
            O => \N__5066\,
            I => \N__5062\
        );

    \I__580\ : InMux
    port map (
            O => \N__5065\,
            I => \N__5059\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__5062\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__5059\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__577\ : InMux
    port map (
            O => \N__5054\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__576\ : InMux
    port map (
            O => \N__5051\,
            I => \N__5047\
        );

    \I__575\ : InMux
    port map (
            O => \N__5050\,
            I => \N__5044\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__5047\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__5044\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__572\ : InMux
    port map (
            O => \N__5039\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__571\ : CascadeMux
    port map (
            O => \N__5036\,
            I => \N__5032\
        );

    \I__570\ : InMux
    port map (
            O => \N__5035\,
            I => \N__5029\
        );

    \I__569\ : InMux
    port map (
            O => \N__5032\,
            I => \N__5026\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__5029\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__5026\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__566\ : InMux
    port map (
            O => \N__5021\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__565\ : InMux
    port map (
            O => \N__5018\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__564\ : InMux
    port map (
            O => \N__5015\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__563\ : InMux
    port map (
            O => \N__5012\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__562\ : ClkMux
    port map (
            O => \N__5009\,
            I => \N__4982\
        );

    \I__561\ : ClkMux
    port map (
            O => \N__5008\,
            I => \N__4982\
        );

    \I__560\ : ClkMux
    port map (
            O => \N__5007\,
            I => \N__4982\
        );

    \I__559\ : ClkMux
    port map (
            O => \N__5006\,
            I => \N__4982\
        );

    \I__558\ : ClkMux
    port map (
            O => \N__5005\,
            I => \N__4982\
        );

    \I__557\ : ClkMux
    port map (
            O => \N__5004\,
            I => \N__4982\
        );

    \I__556\ : ClkMux
    port map (
            O => \N__5003\,
            I => \N__4982\
        );

    \I__555\ : ClkMux
    port map (
            O => \N__5002\,
            I => \N__4982\
        );

    \I__554\ : ClkMux
    port map (
            O => \N__5001\,
            I => \N__4982\
        );

    \I__553\ : GlobalMux
    port map (
            O => \N__4982\,
            I => \N__4979\
        );

    \I__552\ : gio2CtrlBuf
    port map (
            O => \N__4979\,
            I => \C1_c_g\
        );

    \I__551\ : InMux
    port map (
            O => \N__4976\,
            I => \N__4973\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__4973\,
            I => \N__4970\
        );

    \I__549\ : Span4Mux_v
    port map (
            O => \N__4970\,
            I => \N__4967\
        );

    \I__548\ : Span4Mux_v
    port map (
            O => \N__4967\,
            I => \N__4964\
        );

    \I__547\ : Sp12to4
    port map (
            O => \N__4964\,
            I => \N__4961\
        );

    \I__546\ : Span12Mux_h
    port map (
            O => \N__4961\,
            I => \N__4958\
        );

    \I__545\ : Odrv12
    port map (
            O => \N__4958\,
            I => \REGSPACEn_c\
        );

    \I__544\ : InMux
    port map (
            O => \N__4955\,
            I => \N__4950\
        );

    \I__543\ : InMux
    port map (
            O => \N__4954\,
            I => \N__4944\
        );

    \I__542\ : InMux
    port map (
            O => \N__4953\,
            I => \N__4944\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__4950\,
            I => \N__4941\
        );

    \I__540\ : InMux
    port map (
            O => \N__4949\,
            I => \N__4938\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__4944\,
            I => \U712_REG_SM_WRITE_CYCLE\
        );

    \I__538\ : Odrv4
    port map (
            O => \N__4941\,
            I => \U712_REG_SM_WRITE_CYCLE\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__4938\,
            I => \U712_REG_SM_WRITE_CYCLE\
        );

    \I__536\ : IoInMux
    port map (
            O => \N__4931\,
            I => \N__4928\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__4928\,
            I => \N__4925\
        );

    \I__534\ : IoSpan4Mux
    port map (
            O => \N__4925\,
            I => \N__4922\
        );

    \I__533\ : Span4Mux_s3_v
    port map (
            O => \N__4922\,
            I => \N__4919\
        );

    \I__532\ : Sp12to4
    port map (
            O => \N__4919\,
            I => \N__4916\
        );

    \I__531\ : Span12Mux_s11_v
    port map (
            O => \N__4916\,
            I => \N__4912\
        );

    \I__530\ : InMux
    port map (
            O => \N__4915\,
            I => \N__4909\
        );

    \I__529\ : Odrv12
    port map (
            O => \N__4912\,
            I => \PRnW_c\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__4909\,
            I => \PRnW_c\
        );

    \I__527\ : InMux
    port map (
            O => \N__4904\,
            I => \N__4901\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__4901\,
            I => \N__4898\
        );

    \I__525\ : Odrv4
    port map (
            O => \N__4898\,
            I => \U712_CHIP_RAM.N_332\
        );

    \I__524\ : InMux
    port map (
            O => \N__4895\,
            I => \N__4892\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__4892\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\
        );

    \I__522\ : InMux
    port map (
            O => \N__4889\,
            I => \N__4886\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__4886\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_2\
        );

    \I__520\ : IoInMux
    port map (
            O => \N__4883\,
            I => \N__4879\
        );

    \I__519\ : IoInMux
    port map (
            O => \N__4882\,
            I => \N__4875\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__4879\,
            I => \N__4872\
        );

    \I__517\ : IoInMux
    port map (
            O => \N__4878\,
            I => \N__4869\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__4875\,
            I => \N__4866\
        );

    \I__515\ : IoSpan4Mux
    port map (
            O => \N__4872\,
            I => \N__4863\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__4869\,
            I => \N__4860\
        );

    \I__513\ : Span4Mux_s0_h
    port map (
            O => \N__4866\,
            I => \N__4857\
        );

    \I__512\ : Span4Mux_s0_v
    port map (
            O => \N__4863\,
            I => \N__4854\
        );

    \I__511\ : IoSpan4Mux
    port map (
            O => \N__4860\,
            I => \N__4851\
        );

    \I__510\ : Sp12to4
    port map (
            O => \N__4857\,
            I => \N__4848\
        );

    \I__509\ : Span4Mux_v
    port map (
            O => \N__4854\,
            I => \N__4845\
        );

    \I__508\ : IoSpan4Mux
    port map (
            O => \N__4851\,
            I => \N__4842\
        );

    \I__507\ : Span12Mux_v
    port map (
            O => \N__4848\,
            I => \N__4837\
        );

    \I__506\ : Sp12to4
    port map (
            O => \N__4845\,
            I => \N__4834\
        );

    \I__505\ : Span4Mux_s2_v
    port map (
            O => \N__4842\,
            I => \N__4831\
        );

    \I__504\ : InMux
    port map (
            O => \N__4841\,
            I => \N__4828\
        );

    \I__503\ : InMux
    port map (
            O => \N__4840\,
            I => \N__4825\
        );

    \I__502\ : Span12Mux_h
    port map (
            O => \N__4837\,
            I => \N__4816\
        );

    \I__501\ : Span12Mux_h
    port map (
            O => \N__4834\,
            I => \N__4816\
        );

    \I__500\ : Sp12to4
    port map (
            O => \N__4831\,
            I => \N__4816\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__4828\,
            I => \N__4816\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__4825\,
            I => \TACK_EN\
        );

    \I__497\ : Odrv12
    port map (
            O => \N__4816\,
            I => \TACK_EN\
        );

    \I__496\ : SRMux
    port map (
            O => \N__4811\,
            I => \N__4808\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__4808\,
            I => \U712_CYCLE_TERM.TACK_RST_0_i\
        );

    \I__494\ : InMux
    port map (
            O => \N__4805\,
            I => \N__4802\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__4802\,
            I => \U712_REG_SM_STATE_COUNT_7\
        );

    \I__492\ : InMux
    port map (
            O => \N__4799\,
            I => \N__4791\
        );

    \I__491\ : InMux
    port map (
            O => \N__4798\,
            I => \N__4791\
        );

    \I__490\ : InMux
    port map (
            O => \N__4797\,
            I => \N__4786\
        );

    \I__489\ : InMux
    port map (
            O => \N__4796\,
            I => \N__4786\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__4791\,
            I => \U712_REG_SM_STATE_COUNT_0\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__4786\,
            I => \U712_REG_SM_STATE_COUNT_0\
        );

    \I__486\ : InMux
    port map (
            O => \N__4781\,
            I => \N__4778\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__4778\,
            I => \U712_CHIP_RAM.N_79_0\
        );

    \I__484\ : InMux
    port map (
            O => \N__4775\,
            I => \N__4771\
        );

    \I__483\ : InMux
    port map (
            O => \N__4774\,
            I => \N__4768\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__4771\,
            I => \U712_REG_SM_STATE_COUNT_5\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__4768\,
            I => \U712_REG_SM_STATE_COUNT_5\
        );

    \I__480\ : InMux
    port map (
            O => \N__4763\,
            I => \N__4760\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4760\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__478\ : InMux
    port map (
            O => \N__4757\,
            I => \N__4754\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__4754\,
            I => \U712_CHIP_RAM.N_103_0\
        );

    \I__476\ : InMux
    port map (
            O => \N__4751\,
            I => \N__4741\
        );

    \I__475\ : InMux
    port map (
            O => \N__4750\,
            I => \N__4741\
        );

    \I__474\ : InMux
    port map (
            O => \N__4749\,
            I => \N__4736\
        );

    \I__473\ : InMux
    port map (
            O => \N__4748\,
            I => \N__4736\
        );

    \I__472\ : InMux
    port map (
            O => \N__4747\,
            I => \N__4731\
        );

    \I__471\ : InMux
    port map (
            O => \N__4746\,
            I => \N__4731\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__4741\,
            I => \U712_REG_SM_STATE_COUNT_8\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__4736\,
            I => \U712_REG_SM_STATE_COUNT_8\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__4731\,
            I => \U712_REG_SM_STATE_COUNT_8\
        );

    \I__467\ : CascadeMux
    port map (
            O => \N__4724\,
            I => \U712_CHIP_RAM.N_103_0_cascade_\
        );

    \I__466\ : InMux
    port map (
            O => \N__4721\,
            I => \N__4718\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__4718\,
            I => \U712_CHIP_RAM.m106_nsZ0Z_1\
        );

    \I__464\ : InMux
    port map (
            O => \N__4715\,
            I => \N__4712\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__4712\,
            I => i62_mux
        );

    \I__462\ : InMux
    port map (
            O => \N__4709\,
            I => \N__4706\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__4706\,
            I => \N__4702\
        );

    \I__460\ : InMux
    port map (
            O => \N__4705\,
            I => \N__4699\
        );

    \I__459\ : Span12Mux_h
    port map (
            O => \N__4702\,
            I => \N__4696\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__4699\,
            I => \N__4693\
        );

    \I__457\ : Span12Mux_v
    port map (
            O => \N__4696\,
            I => \N__4690\
        );

    \I__456\ : Span12Mux_h
    port map (
            O => \N__4693\,
            I => \N__4687\
        );

    \I__455\ : Odrv12
    port map (
            O => \N__4690\,
            I => \DBRn_c\
        );

    \I__454\ : Odrv12
    port map (
            O => \N__4687\,
            I => \DBRn_c\
        );

    \I__453\ : InMux
    port map (
            O => \N__4682\,
            I => \N__4679\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__4679\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__451\ : IoInMux
    port map (
            O => \N__4676\,
            I => \N__4673\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__4673\,
            I => \N__4670\
        );

    \I__449\ : Odrv12
    port map (
            O => \N__4670\,
            I => \VBENn_c\
        );

    \I__448\ : InMux
    port map (
            O => \N__4667\,
            I => \N__4663\
        );

    \I__447\ : InMux
    port map (
            O => \N__4666\,
            I => \N__4660\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__4663\,
            I => \REG_TACK\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__4660\,
            I => \REG_TACK\
        );

    \I__444\ : InMux
    port map (
            O => \N__4655\,
            I => \N__4652\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__4652\,
            I => \U712_CHIP_RAM_m113_0\
        );

    \I__442\ : CascadeMux
    port map (
            O => \N__4649\,
            I => \N__4646\
        );

    \I__441\ : InMux
    port map (
            O => \N__4646\,
            I => \N__4643\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__4643\,
            I => \U712_CHIP_RAM.N_87_0\
        );

    \I__439\ : CascadeMux
    port map (
            O => \N__4640\,
            I => \U712_CHIP_RAM.N_87_0_cascade_\
        );

    \I__438\ : CascadeMux
    port map (
            O => \N__4637\,
            I => \U712_CHIP_RAM.N_97_0_cascade_\
        );

    \I__437\ : CascadeMux
    port map (
            O => \N__4634\,
            I => \N__4631\
        );

    \I__436\ : InMux
    port map (
            O => \N__4631\,
            I => \N__4628\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__4628\,
            I => \N_112_0\
        );

    \I__434\ : InMux
    port map (
            O => \N__4625\,
            I => \N__4622\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__4622\,
            I => \U712_REG_SM_REG_TACK_7_0\
        );

    \I__432\ : CascadeMux
    port map (
            O => \N__4619\,
            I => \N_19_0_cascade_\
        );

    \I__431\ : InMux
    port map (
            O => \N__4616\,
            I => \N__4608\
        );

    \I__430\ : InMux
    port map (
            O => \N__4615\,
            I => \N__4608\
        );

    \I__429\ : InMux
    port map (
            O => \N__4614\,
            I => \N__4603\
        );

    \I__428\ : InMux
    port map (
            O => \N__4613\,
            I => \N__4603\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__4608\,
            I => \U712_REG_SM_STATE_COUNT_3\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__4603\,
            I => \U712_REG_SM_STATE_COUNT_3\
        );

    \I__425\ : InMux
    port map (
            O => \N__4598\,
            I => \N__4595\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__4595\,
            I => \N_19_0\
        );

    \I__423\ : InMux
    port map (
            O => \N__4592\,
            I => \N__4589\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__4589\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__421\ : IoInMux
    port map (
            O => \N__4586\,
            I => \N__4583\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__4583\,
            I => \N__4580\
        );

    \I__419\ : IoSpan4Mux
    port map (
            O => \N__4580\,
            I => \N__4577\
        );

    \I__418\ : Span4Mux_s3_h
    port map (
            O => \N__4577\,
            I => \N__4574\
        );

    \I__417\ : Span4Mux_v
    port map (
            O => \N__4574\,
            I => \N__4570\
        );

    \I__416\ : InMux
    port map (
            O => \N__4573\,
            I => \N__4567\
        );

    \I__415\ : Span4Mux_h
    port map (
            O => \N__4570\,
            I => \N__4564\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__4567\,
            I => \N__4561\
        );

    \I__413\ : Sp12to4
    port map (
            O => \N__4564\,
            I => \N__4558\
        );

    \I__412\ : Span4Mux_v
    port map (
            O => \N__4561\,
            I => \N__4555\
        );

    \I__411\ : Span12Mux_h
    port map (
            O => \N__4558\,
            I => \N__4550\
        );

    \I__410\ : Sp12to4
    port map (
            O => \N__4555\,
            I => \N__4550\
        );

    \I__409\ : Span12Mux_h
    port map (
            O => \N__4550\,
            I => \N__4547\
        );

    \I__408\ : Odrv12
    port map (
            O => \N__4547\,
            I => \C3_c\
        );

    \I__407\ : InMux
    port map (
            O => \N__4544\,
            I => \N__4541\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__4541\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__405\ : IoInMux
    port map (
            O => \N__4538\,
            I => \N__4535\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__4535\,
            I => \N__4532\
        );

    \I__403\ : Span4Mux_s3_h
    port map (
            O => \N__4532\,
            I => \N__4529\
        );

    \I__402\ : Odrv4
    port map (
            O => \N__4529\,
            I => \DBRn_c_i_0\
        );

    \I__401\ : IoInMux
    port map (
            O => \N__4526\,
            I => \N__4523\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__4523\,
            I => \N__4520\
        );

    \I__399\ : Span4Mux_s2_v
    port map (
            O => \N__4520\,
            I => \N__4517\
        );

    \I__398\ : Span4Mux_v
    port map (
            O => \N__4517\,
            I => \N__4514\
        );

    \I__397\ : Odrv4
    port map (
            O => \N__4514\,
            I => \CLK80_PLL_i_i\
        );

    \I__396\ : IoInMux
    port map (
            O => \N__4511\,
            I => \N__4508\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__4508\,
            I => \N__4505\
        );

    \I__394\ : IoSpan4Mux
    port map (
            O => \N__4505\,
            I => \N__4502\
        );

    \I__393\ : Span4Mux_s2_v
    port map (
            O => \N__4502\,
            I => \N__4499\
        );

    \I__392\ : Sp12to4
    port map (
            O => \N__4499\,
            I => \N__4496\
        );

    \I__391\ : Span12Mux_v
    port map (
            O => \N__4496\,
            I => \N__4493\
        );

    \I__390\ : Odrv12
    port map (
            O => \N__4493\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__5001\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__5004\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            I => \N__5006\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            I => \N__5008\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            I => \N__5009\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            I => \N__5003\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            I => \N__5005\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\,
            I => \N__5007\
        );

    \INVU712_CYCLE_TERM.TACK_OUTC\ : INV
    port map (
            O => \INVU712_CYCLE_TERM.TACK_OUTC_net\,
            I => \N__6867\
        );

    \INVU712_CYCLE_TERM.TACK_ENC\ : INV
    port map (
            O => \INVU712_CYCLE_TERM.TACK_ENC_net\,
            I => \N__6869\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_10_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_14_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_16_0_\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5293\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7922\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4538\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4586\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6064\,
            in2 => \_gnd_net_\,
            in3 => \N__11327\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_3_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11474\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBRn_ibuf_RNIBAB_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4709\,
            lcout => \DBRn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110101010001"
        )
    port map (
            in0 => \N__4625\,
            in1 => \N__4655\,
            in2 => \N__4634\,
            in3 => \N__4666\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11454\,
            ce => 'H',
            sr => \N__11281\
        );

    \U712_CHIP_RAM.m111_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110000100000"
        )
    port map (
            in0 => \N__4748\,
            in1 => \N__5700\,
            in2 => \N__9458\,
            in3 => \N__4613\,
            lcout => \N_112_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m101_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__4749\,
            in1 => \N__4614\,
            in2 => \_gnd_net_\,
            in3 => \N__4955\,
            lcout => \U712_REG_SM_REG_TACK_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m18_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5683\,
            in2 => \_gnd_net_\,
            in3 => \N__9452\,
            lcout => \N_19_0\,
            ltout => \N_19_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110000001000"
        )
    port map (
            in0 => \N__4616\,
            in1 => \N__8109\,
            in2 => \N__4619\,
            in3 => \N__4757\,
            lcout => \U712_REG_SM_STATE_COUNT_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11461\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8110\,
            in1 => \N__4615\,
            in2 => \_gnd_net_\,
            in3 => \N__4598\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11461\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_5_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8111\,
            in2 => \_gnd_net_\,
            in3 => \N__4592\,
            lcout => \U712_REG_SM_STATE_COUNT_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11461\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_0_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4573\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11464\,
            ce => 'H',
            sr => \N__11267\
        );

    \U712_REG_SM.C3_SYNC_1_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4544\,
            lcout => \U712_REG_SM_C3_SYNC_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11464\,
            ce => 'H',
            sr => \N__11267\
        );

    \DBR_SYNC_1_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4682\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11468\,
            ce => 'H',
            sr => \N__11262\
        );

    \DBR_SYNC_0_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4705\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11470\,
            ce => 'H',
            sr => \N__11258\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNI59L8_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__11076\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11122\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_START_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4667\,
            in1 => \N__6629\,
            in2 => \_gnd_net_\,
            in3 => \N__5479\,
            lcout => \U712_CYCLE_TERM.TACK_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11446\,
            ce => 'H',
            sr => \N__4811\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__5050\,
            in1 => \N__5065\,
            in2 => \N__5036\,
            in3 => \N__5080\,
            lcout => \U712_CHIP_RAM.REFRESH5lt7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m113_0_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4774\,
            in2 => \_gnd_net_\,
            in3 => \N__4799\,
            lcout => \U712_CHIP_RAM_m113_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m79_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__9440\,
            in1 => \N__4798\,
            in2 => \N__5215\,
            in3 => \N__5699\,
            lcout => \U712_REG_SM_STATE_COUNT_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_8_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110010001000"
        )
    port map (
            in0 => \N__4805\,
            in1 => \N__8099\,
            in2 => \N__4649\,
            in3 => \N__4751\,
            lcout => \U712_REG_SM_STATE_COUNT_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m86_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__5682\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9425\,
            lcout => \U712_CHIP_RAM.N_87_0\,
            ltout => \U712_CHIP_RAM.N_87_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m96_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4640\,
            in3 => \N__4750\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_97_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011111110101"
        )
    port map (
            in0 => \N__8096\,
            in1 => \N__4781\,
            in2 => \N__4637\,
            in3 => \N__4797\,
            lcout => \U712_REG_SM_STATE_COUNT_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_7_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8098\,
            in2 => \_gnd_net_\,
            in3 => \N__4763\,
            lcout => \U712_REG_SM_STATE_COUNT_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m20_e_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4796\,
            in2 => \_gnd_net_\,
            in3 => \N__5207\,
            lcout => \U712_CHIP_RAM.N_332\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m78_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__5208\,
            in1 => \N__5681\,
            in2 => \_gnd_net_\,
            in3 => \N__9431\,
            lcout => \U712_CHIP_RAM.N_79_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_6_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8097\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4775\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m106_ns_1_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100110011"
        )
    port map (
            in0 => \N__5666\,
            in1 => \N__4949\,
            in2 => \_gnd_net_\,
            in3 => \N__9414\,
            lcout => \U712_CHIP_RAM.m106_nsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__11109\,
            in1 => \N__8100\,
            in2 => \_gnd_net_\,
            in3 => \N__4715\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11462\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m98_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__5665\,
            in1 => \N__5410\,
            in2 => \N__9439\,
            in3 => \N__4746\,
            lcout => \N_99_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m102_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5667\,
            in1 => \N__9415\,
            in2 => \N__6440\,
            in3 => \N__5386\,
            lcout => \U712_CHIP_RAM.N_103_0\,
            ltout => \U712_CHIP_RAM.N_103_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m106_ns_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101100000001"
        )
    port map (
            in0 => \N__4747\,
            in1 => \N__11108\,
            in2 => \N__4724\,
            in3 => \N__4721\,
            lcout => i62_mux,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.WRITE_CYCLE_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__10792\,
            in1 => \N__5239\,
            in2 => \_gnd_net_\,
            in3 => \N__4953\,
            lcout => \U712_REG_SM_WRITE_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11465\,
            ce => 'H',
            sr => \N__11263\
        );

    \U712_REG_SM.PRnW_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111010111001100"
        )
    port map (
            in0 => \N__4954\,
            in1 => \N__4915\,
            in2 => \N__5701\,
            in3 => \N__5723\,
            lcout => \PRnW_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11465\,
            ce => 'H',
            sr => \N__11263\
        );

    \DBR_SYNC_RNITKK4_1_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6406\,
            lcout => \DBR_SYNC_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m85_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__9435\,
            in1 => \N__5411\,
            in2 => \N__5710\,
            in3 => \N__4904\,
            lcout => \N_86_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001100"
        )
    port map (
            in0 => \N__5465\,
            in1 => \N__4840\,
            in2 => \N__5444\,
            in3 => \N__5495\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CYCLE_TERM.TACK_ENC_net\,
            ce => 'H',
            sr => \N__11297\
        );

    \U712_CHIP_RAM.RAS_SYNC_1_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11486\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11439\,
            ce => 'H',
            sr => \N__11282\
        );

    \U712_CHIP_RAM.RAS_SYNC_2_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4895\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11439\,
            ce => 'H',
            sr => \N__11282\
        );

    \U712_CHIP_RAM.RAS_SYNC_3_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4889\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11439\,
            ce => 'H',
            sr => \N__11282\
        );

    \U712_CYCLE_TERM.TACK_START_RNO_0_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8095\,
            in2 => \_gnd_net_\,
            in3 => \N__4841\,
            lcout => \U712_CYCLE_TERM.TACK_RST_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5090\,
            in2 => \_gnd_net_\,
            in3 => \N__5084\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__5002\,
            ce => 'H',
            sr => \N__7118\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5081\,
            in2 => \_gnd_net_\,
            in3 => \N__5069\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__5002\,
            ce => 'H',
            sr => \N__7118\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5066\,
            in2 => \_gnd_net_\,
            in3 => \N__5054\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__5002\,
            ce => 'H',
            sr => \N__7118\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5051\,
            in2 => \_gnd_net_\,
            in3 => \N__5039\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__5002\,
            ce => 'H',
            sr => \N__7118\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5035\,
            in2 => \_gnd_net_\,
            in3 => \N__5021\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__5002\,
            ce => 'H',
            sr => \N__7118\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6247\,
            in2 => \_gnd_net_\,
            in3 => \N__5018\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__5002\,
            ce => 'H',
            sr => \N__7118\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6263\,
            in2 => \_gnd_net_\,
            in3 => \N__5015\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__5002\,
            ce => 'H',
            sr => \N__7118\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6232\,
            in2 => \_gnd_net_\,
            in3 => \N__5012\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5002\,
            ce => 'H',
            sr => \N__7118\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001110011"
        )
    port map (
            in0 => \N__5189\,
            in1 => \N__4976\,
            in2 => \N__5216\,
            in3 => \N__5137\,
            lcout => \U712_REG_SM_REG_CYCLE_START\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11450\,
            ce => 'H',
            sr => \N__11268\
        );

    \U712_REG_SM.START_RST_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__5238\,
            in1 => \N__5188\,
            in2 => \_gnd_net_\,
            in3 => \N__5417\,
            lcout => \U712_REG_SM_START_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11450\,
            ce => 'H',
            sr => \N__11268\
        );

    \U712_CHIP_RAM.RAS_SYNC_5_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5102\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11450\,
            ce => 'H',
            sr => \N__11268\
        );

    \U712_CHIP_RAM.RAS_SYNC_4_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5180\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11450\,
            ce => 'H',
            sr => \N__11268\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011100000101"
        )
    port map (
            in0 => \N__5171\,
            in1 => \N__10992\,
            in2 => \N__5138\,
            in3 => \N__5798\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11450\,
            ce => 'H',
            sr => \N__11268\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIBFJU_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__7279\,
            in1 => \_gnd_net_\,
            in2 => \N__8882\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_363\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIPMTA2_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110100"
        )
    port map (
            in0 => \N__8664\,
            in1 => \N__7280\,
            in2 => \N__6374\,
            in3 => \N__7103\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m223_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRTQU5_3_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__7325\,
            in1 => \N__7748\,
            in2 => \N__5111\,
            in3 => \N__7681\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5108\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5101\,
            lcout => \U712_CHIP_RAM.m231_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__8841\,
            in1 => \N__9124\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_364\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_1_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5258\,
            lcout => \U712_REG_SM_C1_SYNC_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11458\,
            ce => 'H',
            sr => \N__11264\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__5246\,
            in1 => \N__5779\,
            in2 => \_gnd_net_\,
            in3 => \N__7564\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11458\,
            ce => 'H',
            sr => \N__11264\
        );

    \U712_REG_SM.C1_SYNC_0_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5294\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11458\,
            ce => 'H',
            sr => \N__11264\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001100"
        )
    port map (
            in0 => \N__8155\,
            in1 => \N__7282\,
            in2 => \N__10352\,
            in3 => \N__5252\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11458\,
            ce => 'H',
            sr => \N__11264\
        );

    \U712_CHIP_RAM.m77_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001101"
        )
    port map (
            in0 => \N__10155\,
            in1 => \N__10794\,
            in2 => \N__9450\,
            in3 => \N__5732\,
            lcout => \U712_REG_SM_UDSn_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7840\,
            in1 => \N__10793\,
            in2 => \_gnd_net_\,
            in3 => \N__7281\,
            lcout => \U712_CHIP_RAM.N_236\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m82_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5705\,
            in2 => \_gnd_net_\,
            in3 => \N__9426\,
            lcout => \U712_CHIP_RAM.N_83_0\,
            ltout => \U712_CHIP_RAM.N_83_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101010001000"
        )
    port map (
            in0 => \N__8085\,
            in1 => \N__5240\,
            in2 => \N__5219\,
            in3 => \N__5415\,
            lcout => \U712_REG_SM_STATE_COUNT_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11463\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m93_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__5387\,
            in1 => \N__9430\,
            in2 => \N__5711\,
            in3 => \N__6441\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_94_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__8086\,
            in1 => \N__5426\,
            in2 => \N__5420\,
            in3 => \N__5416\,
            lcout => \U712_REG_SM_STATE_COUNT_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11463\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6385\,
            in2 => \N__5374\,
            in3 => \N__5375\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5320\,
            in2 => \_gnd_net_\,
            in3 => \N__5357\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5332\,
            in2 => \_gnd_net_\,
            in3 => \N__5354\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5302\,
            in2 => \_gnd_net_\,
            in3 => \N__5351\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_1_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__8112\,
            in1 => \N__5348\,
            in2 => \N__8156\,
            in3 => \N__6439\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11466\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_2_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__6437\,
            in1 => \N__8113\,
            in2 => \N__5342\,
            in3 => \N__8152\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11466\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__5303\,
            in1 => \N__5333\,
            in2 => \N__5324\,
            in3 => \N__6386\,
            lcout => \U712_CHIP_RAM.N_330\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_3_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__6438\,
            in1 => \N__8114\,
            in2 => \N__5312\,
            in3 => \N__8153\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11466\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m6_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__10077\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9987\,
            lcout => \U712_CHIP_RAM.N_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_ess_RNO_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11324\,
            in2 => \_gnd_net_\,
            in3 => \N__5722\,
            lcout => \U712_REG_SM.N_86_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_ess_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5709\,
            in2 => \_gnd_net_\,
            in3 => \N__9451\,
            lcout => \BLSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11469\,
            ce => \N__5582\,
            sr => \N__11246\
        );

    \U712_CYCLE_TERM.TACK_OUT_RNO_0_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__5439\,
            in1 => \N__5461\,
            in2 => \_gnd_net_\,
            in3 => \N__5493\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_36_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_OUT_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110110011"
        )
    port map (
            in0 => \N__5464\,
            in1 => \N__8080\,
            in2 => \N__5567\,
            in3 => \N__5516\,
            lcout => \TACK_OUT\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CYCLE_TERM.TACK_OUTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__5440\,
            in1 => \N__5463\,
            in2 => \N__8108\,
            in3 => \N__5494\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CYCLE_TERM.TACK_OUTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5462\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8084\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CYCLE_TERM.TACK_OUTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIEG6A1_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__8039\,
            in1 => \N__9130\,
            in2 => \_gnd_net_\,
            in3 => \N__8640\,
            lcout => \U712_CHIP_RAM.m38_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7335\,
            in2 => \_gnd_net_\,
            in3 => \N__6980\,
            lcout => \U712_CHIP_RAM.CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11440\,
            ce => \N__5759\,
            sr => \N__11275\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__8886\,
            in1 => \N__6975\,
            in2 => \N__5939\,
            in3 => \N__9086\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__11325\,
            in1 => \_gnd_net_\,
            in2 => \N__5762\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIIHAH6_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000111111011"
        )
    port map (
            in0 => \N__7303\,
            in1 => \N__7067\,
            in2 => \N__5807\,
            in3 => \N__7018\,
            lcout => \U712_CHIP_RAM.m64_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__7068\,
            in1 => \N__8887\,
            in2 => \N__7823\,
            in3 => \N__8666\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIFK326_0_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8665\,
            in1 => \N__8772\,
            in2 => \_gnd_net_\,
            in3 => \N__7017\,
            lcout => \U712_CHIP_RAM.N_146_0\,
            ltout => \U712_CHIP_RAM.N_146_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__7680\,
            in1 => \N__8888\,
            in2 => \N__5747\,
            in3 => \N__8667\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9087\,
            in2 => \N__5744\,
            in3 => \N__5741\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_154_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111101010111"
        )
    port map (
            in0 => \N__7963\,
            in1 => \N__7139\,
            in2 => \N__5735\,
            in3 => \N__11984\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11444\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIRHVM3_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100000000"
        )
    port map (
            in0 => \N__7094\,
            in1 => \N__5797\,
            in2 => \N__6125\,
            in3 => \N__8771\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_34_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIKHPV5_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111111111"
        )
    port map (
            in0 => \N__5819\,
            in1 => \_gnd_net_\,
            in2 => \N__5810\,
            in3 => \N__7042\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__7093\,
            in1 => \N__6121\,
            in2 => \_gnd_net_\,
            in3 => \N__5795\,
            lcout => \U712_CHIP_RAM.N_359\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNI1EAT_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__8585\,
            in1 => \N__6120\,
            in2 => \_gnd_net_\,
            in3 => \N__5796\,
            lcout => \U712_CHIP_RAM.m41_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__5924\,
            in1 => \N__8047\,
            in2 => \N__5900\,
            in3 => \N__5780\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11447\,
            ce => \N__5850\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__8057\,
            in1 => \N__6185\,
            in2 => \N__8702\,
            in3 => \N__5893\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11451\,
            ce => \N__5855\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_3_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8593\,
            in1 => \N__7746\,
            in2 => \_gnd_net_\,
            in3 => \N__7799\,
            lcout => \U712_CHIP_RAM.N_28_0\,
            ltout => \U712_CHIP_RAM.N_28_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIBDIU5_3_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011111001111"
        )
    port map (
            in0 => \N__7747\,
            in1 => \N__9125\,
            in2 => \N__5768\,
            in3 => \N__6488\,
            lcout => \U712_CHIP_RAM.m66_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__8594\,
            in1 => \N__8873\,
            in2 => \N__7578\,
            in3 => \N__7800\,
            lcout => \U712_CHIP_RAM.N_353_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIA1VV6_1_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__8595\,
            in1 => \N__8874\,
            in2 => \N__8784\,
            in3 => \N__6201\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_47_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIAEA2H_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110101110101"
        )
    port map (
            in0 => \N__8056\,
            in1 => \N__9126\,
            in2 => \N__5765\,
            in3 => \N__6500\,
            lcout => \U712_CHIP_RAM.N_56_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8589\,
            in2 => \_gnd_net_\,
            in3 => \N__6517\,
            lcout => \U712_CHIP_RAM.N_215\,
            ltout => OPEN,
            carryin => \bfn_10_14_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5889\,
            in1 => \N__8872\,
            in2 => \_gnd_net_\,
            in3 => \N__5927\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__11455\,
            ce => \N__5854\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6557\,
            in2 => \_gnd_net_\,
            in3 => \N__5915\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5890\,
            in1 => \N__7749\,
            in2 => \_gnd_net_\,
            in3 => \N__5912\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__11455\,
            ce => \N__5854\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5887\,
            in1 => \N__6586\,
            in2 => \_gnd_net_\,
            in3 => \N__5909\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__11455\,
            ce => \N__5854\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5891\,
            in1 => \N__6599\,
            in2 => \_gnd_net_\,
            in3 => \N__5906\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__11455\,
            ce => \N__5854\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5888\,
            in1 => \N__6611\,
            in2 => \_gnd_net_\,
            in3 => \N__5903\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__11455\,
            ce => \N__5854\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5892\,
            in1 => \N__6572\,
            in2 => \_gnd_net_\,
            in3 => \N__5858\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11455\,
            ce => \N__5854\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001110111"
        )
    port map (
            in0 => \N__8154\,
            in1 => \N__5825\,
            in2 => \_gnd_net_\,
            in3 => \N__6442\,
            lcout => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11459\,
            ce => 'H',
            sr => \N__11255\
        );

    \U712_REG_SM.UDSn_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__6082\,
            in1 => \N__6104\,
            in2 => \_gnd_net_\,
            in3 => \N__8209\,
            lcout => \UDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11459\,
            ce => 'H',
            sr => \N__11255\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__6071\,
            in1 => \N__11845\,
            in2 => \N__11789\,
            in3 => \N__5959\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\,
            ce => 'H',
            sr => \N__11286\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101100000000"
        )
    port map (
            in0 => \N__9617\,
            in1 => \N__12214\,
            in2 => \N__11044\,
            in3 => \N__5945\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11428\,
            ce => \N__9646\,
            sr => \N__11283\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__6019\,
            in1 => \N__12123\,
            in2 => \N__8369\,
            in3 => \N__10939\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m186_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000010000"
        )
    port map (
            in0 => \N__8294\,
            in1 => \N__6173\,
            in2 => \N__5984\,
            in3 => \N__10478\,
            lcout => \U712_CHIP_RAM.m186_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10937\,
            in2 => \_gnd_net_\,
            in3 => \N__12122\,
            lcout => \U712_CHIP_RAM.m186_m2_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011111"
        )
    port map (
            in0 => \N__10938\,
            in1 => \N__5981\,
            in2 => \N__12182\,
            in3 => \N__8354\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m192_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000000010000"
        )
    port map (
            in0 => \N__6179\,
            in1 => \N__8295\,
            in2 => \N__5963\,
            in3 => \N__5960\,
            lcout => \U712_CHIP_RAM.m192_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_8_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__12120\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6278\,
            lcout => \U712_CHIP_RAM.d_N_6_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_0_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__12121\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6314\,
            lcout => \U712_CHIP_RAM.d_N_6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNILLSM_0_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__9221\,
            in1 => \N__12119\,
            in2 => \N__9873\,
            in3 => \N__10915\,
            lcout => \U712_CHIP_RAM.m184_m2_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110100000"
        )
    port map (
            in0 => \N__6167\,
            in1 => \N__8671\,
            in2 => \N__9120\,
            in3 => \N__8786\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_168_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111101010111"
        )
    port map (
            in0 => \N__8037\,
            in1 => \N__7136\,
            in2 => \N__6158\,
            in3 => \N__9884\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11437\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIO6RP9_3_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000100010001"
        )
    port map (
            in0 => \N__8668\,
            in1 => \N__6155\,
            in2 => \N__7772\,
            in3 => \N__7679\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.i67_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNISRNIG_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011101010"
        )
    port map (
            in0 => \N__8914\,
            in1 => \N__9088\,
            in2 => \N__6149\,
            in3 => \N__6146\,
            lcout => \U712_CHIP_RAM.N_67_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__8670\,
            in1 => \N__6137\,
            in2 => \N__7685\,
            in3 => \N__8915\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9089\,
            in2 => \N__6131\,
            in3 => \N__6338\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_151_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111100110111"
        )
    port map (
            in0 => \N__7137\,
            in1 => \N__8038\,
            in2 => \N__6128\,
            in3 => \N__9233\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11437\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000001000100"
        )
    port map (
            in0 => \N__8913\,
            in1 => \N__7070\,
            in2 => \N__7816\,
            in3 => \N__8669\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_0_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6332\,
            in1 => \N__6313\,
            in2 => \_gnd_net_\,
            in3 => \N__8977\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11441\,
            ce => 'H',
            sr => \N__11265\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__8978\,
            in1 => \N__6299\,
            in2 => \N__11782\,
            in3 => \N__6277\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11441\,
            ce => 'H',
            sr => \N__11265\
        );

    \U712_CHIP_RAM.REFRESH_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6262\,
            in1 => \N__6248\,
            in2 => \N__6233\,
            in3 => \N__6215\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11441\,
            ce => 'H',
            sr => \N__11265\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__9102\,
            in1 => \N__8923\,
            in2 => \_gnd_net_\,
            in3 => \N__6206\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11441\,
            ce => 'H',
            sr => \N__11265\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011000000"
        )
    port map (
            in0 => \N__8885\,
            in1 => \N__6350\,
            in2 => \N__9121\,
            in3 => \N__6202\,
            lcout => \U712_CHIP_RAM.N_219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIA7LA2_3_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__6483\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7750\,
            lcout => \U712_CHIP_RAM.N_48_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_2_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__7752\,
            in1 => \N__6556\,
            in2 => \_gnd_net_\,
            in3 => \N__6484\,
            lcout => \U712_CHIP_RAM.N_31_0\,
            ltout => \U712_CHIP_RAM.N_31_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNI50JL4_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__7297\,
            in1 => \N__6367\,
            in2 => \N__6356\,
            in3 => \N__7096\,
            lcout => \U712_CHIP_RAM.N_43_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_0_2_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__7751\,
            in1 => \N__6555\,
            in2 => \_gnd_net_\,
            in3 => \N__6482\,
            lcout => \U712_CHIP_RAM.N_58_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_3_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7802\,
            in1 => \N__8639\,
            in2 => \_gnd_net_\,
            in3 => \N__7756\,
            lcout => \U712_CHIP_RAM.CLK_EN_RNOZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_3_0_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100100010"
        )
    port map (
            in0 => \N__8883\,
            in1 => \N__6518\,
            in2 => \N__7766\,
            in3 => \N__7801\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m217_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110000010100"
        )
    port map (
            in0 => \N__8625\,
            in1 => \N__8884\,
            in2 => \N__6353\,
            in3 => \N__7505\,
            lcout => \U712_CHIP_RAM.N_218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100001111"
        )
    port map (
            in0 => \N__10994\,
            in1 => \N__8628\,
            in2 => \N__8899\,
            in3 => \N__7024\,
            lcout => \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000000100"
        )
    port map (
            in0 => \N__8627\,
            in1 => \N__8867\,
            in2 => \N__7586\,
            in3 => \N__10993\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m212_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000001000"
        )
    port map (
            in0 => \N__8871\,
            in1 => \N__7023\,
            in2 => \N__6344\,
            in3 => \N__7524\,
            lcout => \U712_CHIP_RAM.N_213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI96LA2_0_2_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6545\,
            in2 => \_gnd_net_\,
            in3 => \N__6481\,
            lcout => \U712_CHIP_RAM.N_30_0\,
            ltout => \U712_CHIP_RAM.N_30_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010000100000"
        )
    port map (
            in0 => \N__8866\,
            in1 => \N__8626\,
            in2 => \N__6341\,
            in3 => \N__7022\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__6622\,
            in1 => \N__6641\,
            in2 => \N__9131\,
            in3 => \N__6635\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11448\,
            ce => 'H',
            sr => \N__11259\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6610\,
            in1 => \N__6598\,
            in2 => \N__6587\,
            in3 => \N__6571\,
            lcout => \U712_CHIP_RAM.N_333_mux\,
            ltout => \U712_CHIP_RAM.N_333_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI96LA2_2_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6560\,
            in3 => \N__6544\,
            lcout => \U712_CHIP_RAM.N_26_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNI2E2T2_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__7724\,
            in1 => \N__6554\,
            in2 => \N__7579\,
            in3 => \N__6485\,
            lcout => \U712_CHIP_RAM.N_51_0\,
            ltout => \U712_CHIP_RAM.N_51_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIFI279_1_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011011000100"
        )
    port map (
            in0 => \N__8846\,
            in1 => \N__6494\,
            in2 => \N__6503\,
            in3 => \N__7499\,
            lcout => \U712_CHIP_RAM.N_54_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001100"
        )
    port map (
            in0 => \N__7726\,
            in1 => \N__8845\,
            in2 => \N__8641\,
            in3 => \N__6487\,
            lcout => \U712_CHIP_RAM.m53_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_RNIAPHI2_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6486\,
            in1 => \N__10337\,
            in2 => \_gnd_net_\,
            in3 => \N__7725\,
            lcout => \U712_CHIP_RAM.N_52_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_0_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__8094\,
            in1 => \N__6452\,
            in2 => \N__8148\,
            in3 => \N__6443\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11460\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__11071\,
            in1 => \N__9803\,
            in2 => \N__12228\,
            in3 => \N__6704\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11424\,
            ce => \N__9666\,
            sr => \N__11291\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__11070\,
            in1 => \N__9308\,
            in2 => \N__12227\,
            in3 => \N__6698\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11424\,
            ce => \N__9666\,
            sr => \N__11291\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__8370\,
            in1 => \N__12014\,
            in2 => \_gnd_net_\,
            in3 => \N__12199\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11424\,
            ce => \N__9666\,
            sr => \N__11291\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000000010000"
        )
    port map (
            in0 => \N__6662\,
            in1 => \N__8303\,
            in2 => \N__6959\,
            in3 => \N__9707\,
            lcout => \U712_CHIP_RAM.m189_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010000000100"
        )
    port map (
            in0 => \N__6692\,
            in1 => \N__6668\,
            in2 => \N__8306\,
            in3 => \N__9752\,
            lcout => \U712_CHIP_RAM.m188_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__9242\,
            in1 => \N__12183\,
            in2 => \N__9892\,
            in3 => \N__7364\,
            lcout => \U712_CHIP_RAM.d_N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_3_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__12185\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7430\,
            lcout => \U712_CHIP_RAM.d_N_6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011111"
        )
    port map (
            in0 => \N__11045\,
            in1 => \N__6686\,
            in2 => \N__12225\,
            in3 => \N__8360\,
            lcout => \U712_CHIP_RAM.m188_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_4_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12184\,
            in2 => \_gnd_net_\,
            in3 => \N__7397\,
            lcout => \U712_CHIP_RAM.d_N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111111"
        )
    port map (
            in0 => \N__6656\,
            in1 => \N__11060\,
            in2 => \N__12226\,
            in3 => \N__8361\,
            lcout => \U712_CHIP_RAM.m189_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__6950\,
            in1 => \N__12186\,
            in2 => \N__8371\,
            in3 => \N__11046\,
            lcout => \U712_CHIP_RAM.m185_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__11000\,
            in1 => \N__9608\,
            in2 => \N__12242\,
            in3 => \N__6776\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11427\,
            ce => \N__9645\,
            sr => \N__11278\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__10998\,
            in1 => \N__10463\,
            in2 => \N__12240\,
            in3 => \N__6911\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11427\,
            ce => \N__9645\,
            sr => \N__11278\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101111"
        )
    port map (
            in0 => \N__10999\,
            in1 => \N__10589\,
            in2 => \N__12241\,
            in3 => \N__8399\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11427\,
            ce => \N__9645\,
            sr => \N__11278\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000000111"
        )
    port map (
            in0 => \N__9234\,
            in1 => \N__12148\,
            in2 => \N__12006\,
            in3 => \N__9880\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_198_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__11326\,
            in1 => \_gnd_net_\,
            in2 => \N__6872\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_198_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK40_PLL_derived_clock_RNIIOT_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6868\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_PLL_iso_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010000000100"
        )
    port map (
            in0 => \N__6989\,
            in1 => \N__7160\,
            in2 => \N__8304\,
            in3 => \N__9599\,
            lcout => \U712_CHIP_RAM.m187_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9220\,
            in2 => \_gnd_net_\,
            in3 => \N__9855\,
            lcout => \U712_CHIP_RAM.N_3_0\,
            ltout => \U712_CHIP_RAM.N_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__11004\,
            in1 => \N__7192\,
            in2 => \N__7163\,
            in3 => \N__12163\,
            lcout => \U712_CHIP_RAM.m187_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9122\,
            in1 => \N__7154\,
            in2 => \_gnd_net_\,
            in3 => \N__6995\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_163_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100111111"
        )
    port map (
            in0 => \N__12164\,
            in1 => \N__8061\,
            in2 => \N__7142\,
            in3 => \N__7138\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9228\,
            in1 => \N__9854\,
            in2 => \N__12181\,
            in3 => \N__11996\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__7304\,
            in1 => \N__7095\,
            in2 => \_gnd_net_\,
            in3 => \N__7069\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_158_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__7046\,
            in1 => \N__8676\,
            in2 => \N__7028\,
            in3 => \N__7025\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_2_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12118\,
            in2 => \_gnd_net_\,
            in3 => \N__7459\,
            lcout => \U712_CHIP_RAM.d_N_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIU7TF5_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7336\,
            in2 => \_gnd_net_\,
            in3 => \N__6976\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_2_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7481\,
            in2 => \N__7463\,
            in3 => \N__7460\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11436\,
            ce => 'H',
            sr => \N__11261\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_3_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7448\,
            in1 => \N__7429\,
            in2 => \_gnd_net_\,
            in3 => \N__8974\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11436\,
            ce => 'H',
            sr => \N__11261\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_4_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8975\,
            in1 => \N__7415\,
            in2 => \_gnd_net_\,
            in3 => \N__7393\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11436\,
            ce => 'H',
            sr => \N__11261\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_5_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7379\,
            in1 => \N__7360\,
            in2 => \_gnd_net_\,
            in3 => \N__8976\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11436\,
            ce => 'H',
            sr => \N__11261\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIJD6O3_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7298\,
            in1 => \N__8681\,
            in2 => \_gnd_net_\,
            in3 => \N__8779\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.DMA_CYCLE_START_RNIJD6OZ0Z3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ1M5A_1_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8922\,
            in2 => \N__7346\,
            in3 => \N__7640\,
            lcout => \U712_CHIP_RAM.N_204\,
            ltout => \U712_CHIP_RAM.N_204_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__9103\,
            in1 => \N__7861\,
            in2 => \N__7343\,
            in3 => \N__10331\,
            lcout => \U712_CHIP_RAM.DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11438\,
            ce => 'H',
            sr => \N__11257\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8780\,
            in1 => \N__7340\,
            in2 => \N__8687\,
            in3 => \N__7299\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBDIR_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011111100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7849\,
            in2 => \N__7238\,
            in3 => \N__7216\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11438\,
            ce => 'H',
            sr => \N__11257\
        );

    \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__7862\,
            in1 => \N__10723\,
            in2 => \_gnd_net_\,
            in3 => \N__7850\,
            lcout => \U712_CHIP_RAM.DMA_WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11438\,
            ce => 'H',
            sr => \N__11257\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_1_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8920\,
            in1 => \N__7771\,
            in2 => \N__8680\,
            in3 => \N__7809\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_3_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7770\,
            in2 => \_gnd_net_\,
            in3 => \N__7666\,
            lcout => \U712_CHIP_RAM.N_62_0\,
            ltout => \U712_CHIP_RAM.N_62_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNI9THU5_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__8653\,
            in1 => \N__7580\,
            in2 => \N__7643\,
            in3 => \N__7503\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_RNI9THUZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_2_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7582\,
            in1 => \N__11030\,
            in2 => \N__7529\,
            in3 => \N__8658\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CLK_EN_RNOZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__8921\,
            in1 => \_gnd_net_\,
            in2 => \N__7634\,
            in3 => \N__7631\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_174_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__7597\,
            in1 => \N__9119\,
            in2 => \N__7622\,
            in3 => \N__7619\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11443\,
            ce => 'H',
            sr => \N__11254\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__8654\,
            in1 => \N__7581\,
            in2 => \N__7528\,
            in3 => \N__7504\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_208_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8919\,
            in2 => \N__8213\,
            in3 => \N__9118\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_ess_RNO_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11323\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8202\,
            lcout => \U712_REG_SM.N_99_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__8167\,
            in1 => \N__9341\,
            in2 => \_gnd_net_\,
            in3 => \N__8210\,
            lcout => \LDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11453\,
            ce => 'H',
            sr => \N__11245\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10289\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11456\,
            ce => 'H',
            sr => \N__11244\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8036\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RASn_LC_13_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9241\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11423\,
            ce => 'H',
            sr => \N__11301\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011111110"
        )
    port map (
            in0 => \N__7892\,
            in1 => \N__7886\,
            in2 => \N__8429\,
            in3 => \N__10601\,
            lcout => \U712_CHIP_RAM.m185_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8372\,
            in2 => \_gnd_net_\,
            in3 => \N__12230\,
            lcout => \U712_CHIP_RAM.m194_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__11846\,
            in1 => \N__11942\,
            in2 => \_gnd_net_\,
            in3 => \N__11746\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__11564\,
            sr => \N__11287\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010011"
        )
    port map (
            in0 => \N__11022\,
            in1 => \N__8368\,
            in2 => \N__12229\,
            in3 => \N__7880\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m191_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000000010000"
        )
    port map (
            in0 => \N__8477\,
            in1 => \N__8305\,
            in2 => \N__8486\,
            in3 => \N__8483\,
            lcout => \U712_CHIP_RAM.m191_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_7_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9146\,
            in2 => \_gnd_net_\,
            in3 => \N__12151\,
            lcout => \U712_CHIP_RAM.d_N_6_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100000"
        )
    port map (
            in0 => \N__12152\,
            in1 => \N__8461\,
            in2 => \N__11061\,
            in3 => \N__8355\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m184_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011111110"
        )
    port map (
            in0 => \N__8425\,
            in1 => \N__9176\,
            in2 => \N__8402\,
            in3 => \N__10538\,
            lcout => \U712_CHIP_RAM.m184_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011111"
        )
    port map (
            in0 => \N__12153\,
            in1 => \N__8393\,
            in2 => \N__11062\,
            in3 => \N__8356\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m190_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000010000"
        )
    port map (
            in0 => \N__8299\,
            in1 => \N__8222\,
            in2 => \N__8252\,
            in3 => \N__9590\,
            lcout => \U712_CHIP_RAM.m190_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__9584\,
            in1 => \N__11029\,
            in2 => \N__12224\,
            in3 => \N__8249\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11435\,
            ce => \N__9647\,
            sr => \N__11276\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_6_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8935\,
            in2 => \_gnd_net_\,
            in3 => \N__12150\,
            lcout => \U712_CHIP_RAM.d_N_6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__9232\,
            in1 => \N__12149\,
            in2 => \N__9891\,
            in3 => \N__8992\,
            lcout => \U712_CHIP_RAM.d_N_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_7_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8981\,
            in1 => \N__9167\,
            in2 => \_gnd_net_\,
            in3 => \N__9145\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11442\,
            ce => 'H',
            sr => \N__11266\
        );

    \U712_CHIP_RAM.DBENn_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010111010101010"
        )
    port map (
            in0 => \N__10235\,
            in1 => \N__9123\,
            in2 => \N__8738\,
            in3 => \N__9020\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11442\,
            ce => 'H',
            sr => \N__11266\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_1_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9014\,
            in1 => \N__8993\,
            in2 => \_gnd_net_\,
            in3 => \N__8979\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11442\,
            ce => 'H',
            sr => \N__11266\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_6_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8980\,
            in1 => \N__8948\,
            in2 => \_gnd_net_\,
            in3 => \N__8936\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11442\,
            ce => 'H',
            sr => \N__11266\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__8924\,
            in1 => \N__8785\,
            in2 => \N__8685\,
            in3 => \N__10364\,
            lcout => \U712_CHIP_RAM.DBENn_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__8719\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8672\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__10330\,
            in1 => \N__8497\,
            in2 => \N__8686\,
            in3 => \N__8513\,
            lcout => \LATCH_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11449\,
            ce => 'H',
            sr => \N__11260\
        );

    \U712_REG_SM.ASn_ess_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9457\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11452\,
            ce => \N__9470\,
            sr => \N__11256\
        );

    \U712_CHIP_RAM.m74_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__9938\,
            in1 => \N__10801\,
            in2 => \_gnd_net_\,
            in3 => \N__9453\,
            lcout => \U712_REG_SM_LDSn_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m8_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__9989\,
            in1 => \_gnd_net_\,
            in2 => \N__10097\,
            in3 => \N__10167\,
            lcout => \U712_CHIP_RAM.N_325_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m11_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000111000100"
        )
    port map (
            in0 => \N__10034\,
            in1 => \N__10090\,
            in2 => \N__10169\,
            in3 => \N__9988\,
            lcout => \LMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101111"
        )
    port map (
            in0 => \N__9296\,
            in1 => \N__11043\,
            in2 => \N__12248\,
            in3 => \N__9335\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11426\,
            ce => \N__9667\,
            sr => \N__11298\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11779\,
            in1 => \N__10572\,
            in2 => \_gnd_net_\,
            in3 => \N__9793\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11602\,
            ce => \N__11568\,
            sr => \N__11294\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9743\,
            in1 => \N__11780\,
            in2 => \_gnd_net_\,
            in3 => \N__10630\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11602\,
            ce => \N__11568\,
            sr => \N__11294\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__9290\,
            in1 => \N__9269\,
            in2 => \N__11080\,
            in3 => \N__11615\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11429\,
            ce => \N__9671\,
            sr => \N__11292\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__11855\,
            in1 => \N__11072\,
            in2 => \N__12243\,
            in3 => \N__9698\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11429\,
            ce => \N__9671\,
            sr => \N__11292\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__11828\,
            in1 => \N__11937\,
            in2 => \_gnd_net_\,
            in3 => \N__11706\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11601\,
            ce => \N__11565\,
            sr => \N__11288\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10529\,
            in1 => \N__10571\,
            in2 => \_gnd_net_\,
            in3 => \N__11705\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11601\,
            ce => \N__11565\,
            sr => \N__11288\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10580\,
            in1 => \N__9782\,
            in2 => \_gnd_net_\,
            in3 => \N__11751\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__11562\,
            sr => \N__11284\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__11886\,
            in1 => \N__11936\,
            in2 => \_gnd_net_\,
            in3 => \N__11752\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__11562\,
            sr => \N__11284\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10629\,
            in1 => \N__11750\,
            in2 => \_gnd_net_\,
            in3 => \N__11885\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11597\,
            ce => \N__11560\,
            sr => \N__11279\
        );

    \U712_CHIP_RAM.DBENn_RNI6U6F1_0_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001011111"
        )
    port map (
            in0 => \N__10280\,
            in1 => \N__9910\,
            in2 => \N__10262\,
            in3 => \N__11063\,
            lcout => \CUMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNI8DDB1_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011110101"
        )
    port map (
            in0 => \N__10298\,
            in1 => \N__9547\,
            in2 => \N__10263\,
            in3 => \N__11066\,
            lcout => \CLMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNI8DDB1_0_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111011101"
        )
    port map (
            in0 => \N__11065\,
            in1 => \N__10114\,
            in2 => \N__10264\,
            in3 => \N__10297\,
            lcout => \CUUBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_RNIMKV8_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__10856\,
            in1 => \N__10350\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_346\,
            ltout => \U712_CHIP_RAM.N_346_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNI6U6F1_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101000101"
        )
    port map (
            in0 => \N__11064\,
            in1 => \N__10252\,
            in2 => \N__10217\,
            in3 => \N__10186\,
            lcout => \CLLBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m9_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111000010010"
        )
    port map (
            in0 => \N__10096\,
            in1 => \N__10037\,
            in2 => \N__10000\,
            in3 => \N__9937\,
            lcout => \LLBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m13_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011100000"
        )
    port map (
            in0 => \N__10036\,
            in1 => \N__10168\,
            in2 => \N__10001\,
            in3 => \N__10095\,
            lcout => \UUBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m12_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101101001000"
        )
    port map (
            in0 => \N__10094\,
            in1 => \N__10035\,
            in2 => \N__9999\,
            in3 => \N__9936\,
            lcout => \UMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WEn_LC_15_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9896\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11425\,
            ce => 'H',
            sr => \N__11307\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__9742\,
            in1 => \N__9794\,
            in2 => \_gnd_net_\,
            in3 => \N__11781\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11603\,
            ce => \N__11573\,
            sr => \N__11302\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__9740\,
            in1 => \N__9792\,
            in2 => \_gnd_net_\,
            in3 => \N__11777\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            ce => \N__11571\,
            sr => \N__11299\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11778\,
            in1 => \N__10646\,
            in2 => \_gnd_net_\,
            in3 => \N__9741\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            ce => \N__11571\,
            sr => \N__11299\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11776\,
            in1 => \N__10642\,
            in2 => \_gnd_net_\,
            in3 => \N__11894\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__11569\,
            sr => \N__11295\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11701\,
            in1 => \N__10418\,
            in2 => \_gnd_net_\,
            in3 => \N__10528\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11599\,
            ce => \N__11567\,
            sr => \N__11293\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10579\,
            in1 => \N__10527\,
            in2 => \_gnd_net_\,
            in3 => \N__11749\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__11566\,
            sr => \N__11289\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10413\,
            in1 => \N__10517\,
            in2 => \_gnd_net_\,
            in3 => \N__11748\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__11563\,
            sr => \N__11285\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11747\,
            in1 => \N__10450\,
            in2 => \_gnd_net_\,
            in3 => \N__10417\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11596\,
            ce => \N__11561\,
            sr => \N__11280\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__10451\,
            in1 => \_gnd_net_\,
            in2 => \N__11710\,
            in3 => \N__10409\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__11559\,
            sr => \N__11277\
        );

    \U712_CHIP_RAM.DMA_CYCLE_RNIVA8H_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__10351\,
            in1 => \N__10712\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_345\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__10708\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10852\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11467\,
            ce => 'H',
            sr => \N__11250\
        );

    \U712_CHIP_RAM.DMA_WRITE_CYCLE_RNIVHJN_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__10735\,
            in1 => \N__10707\,
            in2 => \_gnd_net_\,
            in3 => \N__10845\,
            lcout => \DMA_LATCH_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CASn_LC_16_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12247\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11430\,
            ce => 'H',
            sr => \N__11306\
        );

    \U712_CHIP_RAM.CRCSn_LC_16_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12013\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11430\,
            ce => 'H',
            sr => \N__11306\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__11938\,
            in1 => \N__11893\,
            in2 => \_gnd_net_\,
            in3 => \N__11775\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11600\,
            ce => \N__11572\,
            sr => \N__11300\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__11841\,
            in1 => \N__11521\,
            in2 => \_gnd_net_\,
            in3 => \N__11700\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11598\,
            ce => \N__11570\,
            sr => \N__11296\
        );

    \U712_CHIP_RAM.RAS_SYNC_0_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11522\,
            in2 => \_gnd_net_\,
            in3 => \N__11498\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11445\,
            ce => 'H',
            sr => \N__11290\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNIQ44J_LC_24_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000000"
        )
    port map (
            in0 => \N__11129\,
            in1 => \N__10683\,
            in2 => \N__10836\,
            in3 => \N__11087\,
            lcout => \N_338_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_WRITE_CYCLE_RNIRVG61_LC_24_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100001111"
        )
    port map (
            in0 => \N__10830\,
            in1 => \N__10802\,
            in2 => \N__10742\,
            in3 => \N__10684\,
            lcout => \N_328_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jun 13 2025 15:27:47

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U400_TOP" view "INTERFACE"

module U400_TOP (
    SIZ,
    MA,
    A,
    LBENn,
    CS0n,
    UUBEn,
    TAn,
    CLK40,
    RnW,
    BANK1,
    UMBEn,
    WEn,
    LLBEn,
    TSn,
    LMBEn,
    RASn,
    CS1n,
    RESETn,
    CLK_EN,
    CASn,
    BANK0);

    input [1:0] SIZ;
    output [12:0] MA;
    input [31:0] A;
    output LBENn;
    output CS0n;
    output UUBEn;
    output TAn;
    input CLK40;
    input RnW;
    output BANK1;
    output UMBEn;
    output WEn;
    output LLBEn;
    input TSn;
    output LMBEn;
    output RASn;
    output CS1n;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;

    wire N__7125;
    wire N__7124;
    wire N__7123;
    wire N__7116;
    wire N__7115;
    wire N__7114;
    wire N__7107;
    wire N__7106;
    wire N__7105;
    wire N__7098;
    wire N__7097;
    wire N__7096;
    wire N__7089;
    wire N__7088;
    wire N__7087;
    wire N__7080;
    wire N__7079;
    wire N__7078;
    wire N__7071;
    wire N__7070;
    wire N__7069;
    wire N__7062;
    wire N__7061;
    wire N__7060;
    wire N__7053;
    wire N__7052;
    wire N__7051;
    wire N__7044;
    wire N__7043;
    wire N__7042;
    wire N__7035;
    wire N__7034;
    wire N__7033;
    wire N__7026;
    wire N__7025;
    wire N__7024;
    wire N__7017;
    wire N__7016;
    wire N__7015;
    wire N__7008;
    wire N__7007;
    wire N__7006;
    wire N__6999;
    wire N__6998;
    wire N__6997;
    wire N__6990;
    wire N__6989;
    wire N__6988;
    wire N__6981;
    wire N__6980;
    wire N__6979;
    wire N__6972;
    wire N__6971;
    wire N__6970;
    wire N__6963;
    wire N__6962;
    wire N__6961;
    wire N__6954;
    wire N__6953;
    wire N__6952;
    wire N__6945;
    wire N__6944;
    wire N__6943;
    wire N__6936;
    wire N__6935;
    wire N__6934;
    wire N__6927;
    wire N__6926;
    wire N__6925;
    wire N__6918;
    wire N__6917;
    wire N__6916;
    wire N__6909;
    wire N__6908;
    wire N__6907;
    wire N__6900;
    wire N__6899;
    wire N__6898;
    wire N__6891;
    wire N__6890;
    wire N__6889;
    wire N__6882;
    wire N__6881;
    wire N__6880;
    wire N__6873;
    wire N__6872;
    wire N__6871;
    wire N__6864;
    wire N__6863;
    wire N__6862;
    wire N__6855;
    wire N__6854;
    wire N__6853;
    wire N__6846;
    wire N__6845;
    wire N__6844;
    wire N__6837;
    wire N__6836;
    wire N__6835;
    wire N__6828;
    wire N__6827;
    wire N__6826;
    wire N__6819;
    wire N__6818;
    wire N__6817;
    wire N__6810;
    wire N__6809;
    wire N__6808;
    wire N__6801;
    wire N__6800;
    wire N__6799;
    wire N__6792;
    wire N__6791;
    wire N__6790;
    wire N__6783;
    wire N__6782;
    wire N__6781;
    wire N__6774;
    wire N__6773;
    wire N__6772;
    wire N__6765;
    wire N__6764;
    wire N__6763;
    wire N__6756;
    wire N__6755;
    wire N__6754;
    wire N__6747;
    wire N__6746;
    wire N__6745;
    wire N__6738;
    wire N__6737;
    wire N__6736;
    wire N__6729;
    wire N__6728;
    wire N__6727;
    wire N__6720;
    wire N__6719;
    wire N__6718;
    wire N__6711;
    wire N__6710;
    wire N__6709;
    wire N__6702;
    wire N__6701;
    wire N__6700;
    wire N__6693;
    wire N__6692;
    wire N__6691;
    wire N__6684;
    wire N__6683;
    wire N__6682;
    wire N__6675;
    wire N__6674;
    wire N__6673;
    wire N__6666;
    wire N__6665;
    wire N__6664;
    wire N__6657;
    wire N__6656;
    wire N__6655;
    wire N__6648;
    wire N__6647;
    wire N__6646;
    wire N__6639;
    wire N__6638;
    wire N__6637;
    wire N__6630;
    wire N__6629;
    wire N__6628;
    wire N__6621;
    wire N__6620;
    wire N__6619;
    wire N__6612;
    wire N__6611;
    wire N__6610;
    wire N__6603;
    wire N__6602;
    wire N__6601;
    wire N__6594;
    wire N__6593;
    wire N__6592;
    wire N__6585;
    wire N__6584;
    wire N__6583;
    wire N__6576;
    wire N__6575;
    wire N__6574;
    wire N__6567;
    wire N__6566;
    wire N__6565;
    wire N__6558;
    wire N__6557;
    wire N__6556;
    wire N__6549;
    wire N__6548;
    wire N__6547;
    wire N__6530;
    wire N__6527;
    wire N__6524;
    wire N__6521;
    wire N__6518;
    wire N__6515;
    wire N__6512;
    wire N__6509;
    wire N__6506;
    wire N__6503;
    wire N__6502;
    wire N__6501;
    wire N__6500;
    wire N__6499;
    wire N__6498;
    wire N__6497;
    wire N__6496;
    wire N__6495;
    wire N__6492;
    wire N__6491;
    wire N__6490;
    wire N__6489;
    wire N__6486;
    wire N__6485;
    wire N__6482;
    wire N__6479;
    wire N__6476;
    wire N__6475;
    wire N__6474;
    wire N__6469;
    wire N__6466;
    wire N__6463;
    wire N__6462;
    wire N__6459;
    wire N__6454;
    wire N__6451;
    wire N__6450;
    wire N__6447;
    wire N__6444;
    wire N__6437;
    wire N__6432;
    wire N__6427;
    wire N__6426;
    wire N__6425;
    wire N__6422;
    wire N__6419;
    wire N__6412;
    wire N__6409;
    wire N__6400;
    wire N__6397;
    wire N__6394;
    wire N__6391;
    wire N__6386;
    wire N__6379;
    wire N__6368;
    wire N__6365;
    wire N__6362;
    wire N__6359;
    wire N__6356;
    wire N__6353;
    wire N__6350;
    wire N__6347;
    wire N__6344;
    wire N__6341;
    wire N__6338;
    wire N__6337;
    wire N__6336;
    wire N__6335;
    wire N__6334;
    wire N__6333;
    wire N__6332;
    wire N__6331;
    wire N__6328;
    wire N__6325;
    wire N__6316;
    wire N__6311;
    wire N__6310;
    wire N__6307;
    wire N__6304;
    wire N__6301;
    wire N__6298;
    wire N__6295;
    wire N__6290;
    wire N__6287;
    wire N__6278;
    wire N__6275;
    wire N__6272;
    wire N__6269;
    wire N__6268;
    wire N__6267;
    wire N__6266;
    wire N__6265;
    wire N__6262;
    wire N__6259;
    wire N__6258;
    wire N__6255;
    wire N__6254;
    wire N__6251;
    wire N__6248;
    wire N__6245;
    wire N__6242;
    wire N__6241;
    wire N__6238;
    wire N__6237;
    wire N__6234;
    wire N__6231;
    wire N__6228;
    wire N__6225;
    wire N__6220;
    wire N__6217;
    wire N__6214;
    wire N__6211;
    wire N__6206;
    wire N__6191;
    wire N__6188;
    wire N__6187;
    wire N__6184;
    wire N__6181;
    wire N__6180;
    wire N__6179;
    wire N__6178;
    wire N__6177;
    wire N__6174;
    wire N__6173;
    wire N__6172;
    wire N__6171;
    wire N__6170;
    wire N__6169;
    wire N__6166;
    wire N__6165;
    wire N__6164;
    wire N__6163;
    wire N__6162;
    wire N__6161;
    wire N__6160;
    wire N__6159;
    wire N__6158;
    wire N__6157;
    wire N__6116;
    wire N__6113;
    wire N__6110;
    wire N__6107;
    wire N__6104;
    wire N__6101;
    wire N__6098;
    wire N__6095;
    wire N__6092;
    wire N__6089;
    wire N__6086;
    wire N__6083;
    wire N__6080;
    wire N__6077;
    wire N__6076;
    wire N__6075;
    wire N__6074;
    wire N__6071;
    wire N__6070;
    wire N__6069;
    wire N__6068;
    wire N__6067;
    wire N__6064;
    wire N__6063;
    wire N__6062;
    wire N__6059;
    wire N__6056;
    wire N__6053;
    wire N__6050;
    wire N__6047;
    wire N__6044;
    wire N__6041;
    wire N__6040;
    wire N__6037;
    wire N__6032;
    wire N__6031;
    wire N__6022;
    wire N__6017;
    wire N__6014;
    wire N__6011;
    wire N__6006;
    wire N__6003;
    wire N__6000;
    wire N__5991;
    wire N__5984;
    wire N__5981;
    wire N__5978;
    wire N__5975;
    wire N__5972;
    wire N__5969;
    wire N__5968;
    wire N__5967;
    wire N__5964;
    wire N__5961;
    wire N__5960;
    wire N__5959;
    wire N__5958;
    wire N__5957;
    wire N__5956;
    wire N__5955;
    wire N__5954;
    wire N__5951;
    wire N__5948;
    wire N__5945;
    wire N__5942;
    wire N__5939;
    wire N__5936;
    wire N__5933;
    wire N__5930;
    wire N__5925;
    wire N__5924;
    wire N__5921;
    wire N__5918;
    wire N__5913;
    wire N__5906;
    wire N__5901;
    wire N__5898;
    wire N__5895;
    wire N__5890;
    wire N__5885;
    wire N__5876;
    wire N__5873;
    wire N__5870;
    wire N__5867;
    wire N__5866;
    wire N__5861;
    wire N__5858;
    wire N__5857;
    wire N__5854;
    wire N__5853;
    wire N__5850;
    wire N__5847;
    wire N__5844;
    wire N__5841;
    wire N__5838;
    wire N__5833;
    wire N__5828;
    wire N__5825;
    wire N__5824;
    wire N__5823;
    wire N__5822;
    wire N__5819;
    wire N__5816;
    wire N__5813;
    wire N__5812;
    wire N__5811;
    wire N__5808;
    wire N__5805;
    wire N__5800;
    wire N__5795;
    wire N__5790;
    wire N__5787;
    wire N__5784;
    wire N__5781;
    wire N__5776;
    wire N__5771;
    wire N__5770;
    wire N__5767;
    wire N__5762;
    wire N__5759;
    wire N__5758;
    wire N__5757;
    wire N__5756;
    wire N__5755;
    wire N__5752;
    wire N__5749;
    wire N__5748;
    wire N__5745;
    wire N__5742;
    wire N__5739;
    wire N__5736;
    wire N__5731;
    wire N__5728;
    wire N__5725;
    wire N__5718;
    wire N__5715;
    wire N__5712;
    wire N__5709;
    wire N__5704;
    wire N__5701;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5687;
    wire N__5684;
    wire N__5681;
    wire N__5678;
    wire N__5675;
    wire N__5672;
    wire N__5669;
    wire N__5666;
    wire N__5663;
    wire N__5660;
    wire N__5657;
    wire N__5654;
    wire N__5651;
    wire N__5648;
    wire N__5645;
    wire N__5642;
    wire N__5639;
    wire N__5636;
    wire N__5633;
    wire N__5630;
    wire N__5627;
    wire N__5624;
    wire N__5621;
    wire N__5618;
    wire N__5615;
    wire N__5612;
    wire N__5609;
    wire N__5606;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5594;
    wire N__5591;
    wire N__5588;
    wire N__5585;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5570;
    wire N__5567;
    wire N__5564;
    wire N__5561;
    wire N__5558;
    wire N__5555;
    wire N__5552;
    wire N__5551;
    wire N__5550;
    wire N__5549;
    wire N__5548;
    wire N__5547;
    wire N__5546;
    wire N__5545;
    wire N__5544;
    wire N__5539;
    wire N__5534;
    wire N__5533;
    wire N__5530;
    wire N__5529;
    wire N__5528;
    wire N__5527;
    wire N__5524;
    wire N__5523;
    wire N__5522;
    wire N__5521;
    wire N__5520;
    wire N__5517;
    wire N__5516;
    wire N__5513;
    wire N__5510;
    wire N__5505;
    wire N__5500;
    wire N__5497;
    wire N__5494;
    wire N__5491;
    wire N__5484;
    wire N__5477;
    wire N__5474;
    wire N__5471;
    wire N__5468;
    wire N__5465;
    wire N__5458;
    wire N__5457;
    wire N__5456;
    wire N__5449;
    wire N__5446;
    wire N__5441;
    wire N__5436;
    wire N__5431;
    wire N__5428;
    wire N__5423;
    wire N__5414;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5398;
    wire N__5397;
    wire N__5396;
    wire N__5395;
    wire N__5394;
    wire N__5393;
    wire N__5392;
    wire N__5391;
    wire N__5388;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5370;
    wire N__5367;
    wire N__5354;
    wire N__5351;
    wire N__5350;
    wire N__5349;
    wire N__5346;
    wire N__5341;
    wire N__5336;
    wire N__5333;
    wire N__5330;
    wire N__5327;
    wire N__5324;
    wire N__5321;
    wire N__5318;
    wire N__5315;
    wire N__5312;
    wire N__5309;
    wire N__5306;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5294;
    wire N__5291;
    wire N__5288;
    wire N__5285;
    wire N__5282;
    wire N__5279;
    wire N__5276;
    wire N__5273;
    wire N__5270;
    wire N__5267;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5255;
    wire N__5252;
    wire N__5249;
    wire N__5246;
    wire N__5245;
    wire N__5242;
    wire N__5239;
    wire N__5238;
    wire N__5235;
    wire N__5232;
    wire N__5229;
    wire N__5226;
    wire N__5223;
    wire N__5220;
    wire N__5217;
    wire N__5214;
    wire N__5211;
    wire N__5208;
    wire N__5203;
    wire N__5198;
    wire N__5195;
    wire N__5194;
    wire N__5193;
    wire N__5190;
    wire N__5187;
    wire N__5184;
    wire N__5183;
    wire N__5180;
    wire N__5177;
    wire N__5174;
    wire N__5171;
    wire N__5168;
    wire N__5159;
    wire N__5156;
    wire N__5153;
    wire N__5150;
    wire N__5147;
    wire N__5144;
    wire N__5143;
    wire N__5140;
    wire N__5137;
    wire N__5134;
    wire N__5131;
    wire N__5128;
    wire N__5123;
    wire N__5120;
    wire N__5117;
    wire N__5116;
    wire N__5113;
    wire N__5110;
    wire N__5107;
    wire N__5104;
    wire N__5101;
    wire N__5098;
    wire N__5095;
    wire N__5090;
    wire N__5087;
    wire N__5084;
    wire N__5083;
    wire N__5080;
    wire N__5077;
    wire N__5072;
    wire N__5069;
    wire N__5066;
    wire N__5063;
    wire N__5060;
    wire N__5057;
    wire N__5054;
    wire N__5051;
    wire N__5048;
    wire N__5047;
    wire N__5046;
    wire N__5045;
    wire N__5044;
    wire N__5043;
    wire N__5040;
    wire N__5039;
    wire N__5036;
    wire N__5031;
    wire N__5028;
    wire N__5025;
    wire N__5022;
    wire N__5019;
    wire N__5016;
    wire N__5003;
    wire N__5002;
    wire N__5001;
    wire N__5000;
    wire N__4999;
    wire N__4998;
    wire N__4997;
    wire N__4996;
    wire N__4995;
    wire N__4990;
    wire N__4987;
    wire N__4984;
    wire N__4975;
    wire N__4972;
    wire N__4961;
    wire N__4958;
    wire N__4955;
    wire N__4952;
    wire N__4949;
    wire N__4948;
    wire N__4947;
    wire N__4946;
    wire N__4943;
    wire N__4942;
    wire N__4941;
    wire N__4940;
    wire N__4937;
    wire N__4932;
    wire N__4931;
    wire N__4930;
    wire N__4927;
    wire N__4926;
    wire N__4925;
    wire N__4920;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4910;
    wire N__4909;
    wire N__4908;
    wire N__4907;
    wire N__4902;
    wire N__4901;
    wire N__4900;
    wire N__4899;
    wire N__4898;
    wire N__4895;
    wire N__4892;
    wire N__4889;
    wire N__4884;
    wire N__4881;
    wire N__4878;
    wire N__4871;
    wire N__4868;
    wire N__4865;
    wire N__4862;
    wire N__4857;
    wire N__4854;
    wire N__4845;
    wire N__4826;
    wire N__4823;
    wire N__4820;
    wire N__4819;
    wire N__4818;
    wire N__4817;
    wire N__4814;
    wire N__4813;
    wire N__4810;
    wire N__4809;
    wire N__4808;
    wire N__4807;
    wire N__4806;
    wire N__4803;
    wire N__4800;
    wire N__4799;
    wire N__4798;
    wire N__4797;
    wire N__4796;
    wire N__4795;
    wire N__4794;
    wire N__4791;
    wire N__4790;
    wire N__4789;
    wire N__4786;
    wire N__4785;
    wire N__4782;
    wire N__4775;
    wire N__4774;
    wire N__4773;
    wire N__4770;
    wire N__4765;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4748;
    wire N__4745;
    wire N__4742;
    wire N__4739;
    wire N__4734;
    wire N__4731;
    wire N__4728;
    wire N__4725;
    wire N__4722;
    wire N__4717;
    wire N__4688;
    wire N__4687;
    wire N__4684;
    wire N__4681;
    wire N__4680;
    wire N__4679;
    wire N__4678;
    wire N__4675;
    wire N__4672;
    wire N__4671;
    wire N__4668;
    wire N__4665;
    wire N__4664;
    wire N__4663;
    wire N__4660;
    wire N__4659;
    wire N__4656;
    wire N__4653;
    wire N__4650;
    wire N__4647;
    wire N__4640;
    wire N__4635;
    wire N__4630;
    wire N__4619;
    wire N__4618;
    wire N__4617;
    wire N__4616;
    wire N__4615;
    wire N__4612;
    wire N__4611;
    wire N__4610;
    wire N__4609;
    wire N__4608;
    wire N__4605;
    wire N__4602;
    wire N__4599;
    wire N__4598;
    wire N__4597;
    wire N__4596;
    wire N__4593;
    wire N__4592;
    wire N__4591;
    wire N__4590;
    wire N__4589;
    wire N__4588;
    wire N__4587;
    wire N__4580;
    wire N__4575;
    wire N__4574;
    wire N__4573;
    wire N__4572;
    wire N__4569;
    wire N__4566;
    wire N__4561;
    wire N__4558;
    wire N__4555;
    wire N__4550;
    wire N__4547;
    wire N__4540;
    wire N__4537;
    wire N__4532;
    wire N__4529;
    wire N__4524;
    wire N__4517;
    wire N__4514;
    wire N__4493;
    wire N__4492;
    wire N__4491;
    wire N__4490;
    wire N__4489;
    wire N__4488;
    wire N__4485;
    wire N__4482;
    wire N__4479;
    wire N__4474;
    wire N__4473;
    wire N__4470;
    wire N__4469;
    wire N__4468;
    wire N__4463;
    wire N__4462;
    wire N__4461;
    wire N__4456;
    wire N__4453;
    wire N__4450;
    wire N__4445;
    wire N__4444;
    wire N__4443;
    wire N__4442;
    wire N__4441;
    wire N__4438;
    wire N__4435;
    wire N__4432;
    wire N__4429;
    wire N__4426;
    wire N__4421;
    wire N__4414;
    wire N__4411;
    wire N__4394;
    wire N__4393;
    wire N__4390;
    wire N__4387;
    wire N__4382;
    wire N__4381;
    wire N__4380;
    wire N__4377;
    wire N__4374;
    wire N__4371;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire N__4357;
    wire N__4356;
    wire N__4353;
    wire N__4350;
    wire N__4349;
    wire N__4346;
    wire N__4341;
    wire N__4338;
    wire N__4337;
    wire N__4336;
    wire N__4335;
    wire N__4334;
    wire N__4333;
    wire N__4332;
    wire N__4331;
    wire N__4328;
    wire N__4325;
    wire N__4322;
    wire N__4317;
    wire N__4308;
    wire N__4305;
    wire N__4292;
    wire N__4289;
    wire N__4288;
    wire N__4285;
    wire N__4284;
    wire N__4281;
    wire N__4280;
    wire N__4279;
    wire N__4278;
    wire N__4273;
    wire N__4270;
    wire N__4263;
    wire N__4256;
    wire N__4255;
    wire N__4254;
    wire N__4253;
    wire N__4250;
    wire N__4249;
    wire N__4246;
    wire N__4243;
    wire N__4240;
    wire N__4237;
    wire N__4230;
    wire N__4223;
    wire N__4222;
    wire N__4219;
    wire N__4218;
    wire N__4217;
    wire N__4214;
    wire N__4213;
    wire N__4212;
    wire N__4207;
    wire N__4204;
    wire N__4197;
    wire N__4190;
    wire N__4189;
    wire N__4186;
    wire N__4183;
    wire N__4178;
    wire N__4177;
    wire N__4174;
    wire N__4173;
    wire N__4172;
    wire N__4171;
    wire N__4168;
    wire N__4163;
    wire N__4158;
    wire N__4151;
    wire N__4150;
    wire N__4149;
    wire N__4148;
    wire N__4147;
    wire N__4146;
    wire N__4143;
    wire N__4138;
    wire N__4135;
    wire N__4130;
    wire N__4121;
    wire N__4118;
    wire N__4117;
    wire N__4112;
    wire N__4109;
    wire N__4108;
    wire N__4107;
    wire N__4106;
    wire N__4105;
    wire N__4104;
    wire N__4103;
    wire N__4102;
    wire N__4095;
    wire N__4092;
    wire N__4083;
    wire N__4076;
    wire N__4075;
    wire N__4074;
    wire N__4073;
    wire N__4072;
    wire N__4071;
    wire N__4070;
    wire N__4069;
    wire N__4068;
    wire N__4067;
    wire N__4066;
    wire N__4065;
    wire N__4064;
    wire N__4063;
    wire N__4062;
    wire N__4061;
    wire N__4060;
    wire N__4059;
    wire N__4058;
    wire N__4057;
    wire N__4056;
    wire N__4055;
    wire N__4054;
    wire N__4053;
    wire N__4052;
    wire N__4051;
    wire N__4050;
    wire N__3995;
    wire N__3992;
    wire N__3989;
    wire N__3986;
    wire N__3983;
    wire N__3982;
    wire N__3981;
    wire N__3980;
    wire N__3977;
    wire N__3974;
    wire N__3971;
    wire N__3970;
    wire N__3969;
    wire N__3968;
    wire N__3967;
    wire N__3966;
    wire N__3965;
    wire N__3962;
    wire N__3959;
    wire N__3956;
    wire N__3953;
    wire N__3952;
    wire N__3943;
    wire N__3942;
    wire N__3941;
    wire N__3940;
    wire N__3937;
    wire N__3936;
    wire N__3933;
    wire N__3932;
    wire N__3931;
    wire N__3930;
    wire N__3927;
    wire N__3920;
    wire N__3917;
    wire N__3914;
    wire N__3911;
    wire N__3908;
    wire N__3903;
    wire N__3896;
    wire N__3893;
    wire N__3890;
    wire N__3887;
    wire N__3882;
    wire N__3877;
    wire N__3870;
    wire N__3865;
    wire N__3860;
    wire N__3857;
    wire N__3854;
    wire N__3851;
    wire N__3848;
    wire N__3845;
    wire N__3842;
    wire N__3833;
    wire N__3830;
    wire N__3829;
    wire N__3826;
    wire N__3823;
    wire N__3818;
    wire N__3815;
    wire N__3814;
    wire N__3811;
    wire N__3808;
    wire N__3803;
    wire N__3800;
    wire N__3799;
    wire N__3796;
    wire N__3793;
    wire N__3792;
    wire N__3789;
    wire N__3786;
    wire N__3783;
    wire N__3778;
    wire N__3773;
    wire N__3770;
    wire N__3769;
    wire N__3766;
    wire N__3763;
    wire N__3760;
    wire N__3757;
    wire N__3752;
    wire N__3749;
    wire N__3746;
    wire N__3743;
    wire N__3740;
    wire N__3739;
    wire N__3738;
    wire N__3735;
    wire N__3732;
    wire N__3729;
    wire N__3722;
    wire N__3719;
    wire N__3716;
    wire N__3713;
    wire N__3710;
    wire N__3707;
    wire N__3706;
    wire N__3703;
    wire N__3700;
    wire N__3695;
    wire N__3692;
    wire N__3689;
    wire N__3686;
    wire N__3683;
    wire N__3680;
    wire N__3677;
    wire N__3674;
    wire N__3671;
    wire N__3668;
    wire N__3665;
    wire N__3662;
    wire N__3661;
    wire N__3658;
    wire N__3655;
    wire N__3650;
    wire N__3649;
    wire N__3644;
    wire N__3641;
    wire N__3638;
    wire N__3635;
    wire N__3632;
    wire N__3631;
    wire N__3628;
    wire N__3625;
    wire N__3622;
    wire N__3619;
    wire N__3614;
    wire N__3611;
    wire N__3608;
    wire N__3605;
    wire N__3602;
    wire N__3599;
    wire N__3596;
    wire N__3593;
    wire N__3590;
    wire N__3587;
    wire N__3584;
    wire N__3581;
    wire N__3578;
    wire N__3575;
    wire N__3572;
    wire N__3571;
    wire N__3570;
    wire N__3563;
    wire N__3560;
    wire N__3557;
    wire N__3554;
    wire N__3551;
    wire N__3550;
    wire N__3545;
    wire N__3542;
    wire N__3539;
    wire N__3536;
    wire N__3533;
    wire N__3530;
    wire N__3527;
    wire N__3524;
    wire N__3521;
    wire N__3520;
    wire N__3515;
    wire N__3512;
    wire N__3511;
    wire N__3508;
    wire N__3503;
    wire N__3500;
    wire N__3499;
    wire N__3498;
    wire N__3497;
    wire N__3496;
    wire N__3493;
    wire N__3492;
    wire N__3491;
    wire N__3490;
    wire N__3487;
    wire N__3480;
    wire N__3475;
    wire N__3470;
    wire N__3467;
    wire N__3458;
    wire N__3455;
    wire N__3452;
    wire N__3449;
    wire N__3446;
    wire N__3445;
    wire N__3444;
    wire N__3441;
    wire N__3438;
    wire N__3435;
    wire N__3428;
    wire N__3425;
    wire N__3422;
    wire N__3421;
    wire N__3420;
    wire N__3419;
    wire N__3416;
    wire N__3413;
    wire N__3410;
    wire N__3407;
    wire N__3398;
    wire N__3395;
    wire N__3392;
    wire N__3389;
    wire N__3386;
    wire N__3383;
    wire N__3380;
    wire N__3377;
    wire N__3374;
    wire N__3371;
    wire N__3368;
    wire N__3367;
    wire N__3364;
    wire N__3361;
    wire N__3356;
    wire N__3353;
    wire N__3350;
    wire N__3347;
    wire N__3344;
    wire N__3341;
    wire N__3340;
    wire N__3337;
    wire N__3334;
    wire N__3329;
    wire N__3326;
    wire N__3323;
    wire N__3320;
    wire N__3317;
    wire N__3316;
    wire N__3313;
    wire N__3310;
    wire N__3305;
    wire N__3302;
    wire N__3299;
    wire N__3296;
    wire N__3293;
    wire N__3290;
    wire N__3287;
    wire N__3284;
    wire N__3281;
    wire N__3278;
    wire N__3275;
    wire N__3272;
    wire N__3271;
    wire N__3268;
    wire N__3265;
    wire N__3260;
    wire N__3259;
    wire N__3258;
    wire N__3251;
    wire N__3248;
    wire N__3245;
    wire N__3242;
    wire N__3239;
    wire N__3236;
    wire N__3233;
    wire N__3230;
    wire N__3227;
    wire N__3224;
    wire N__3221;
    wire N__3218;
    wire N__3215;
    wire N__3212;
    wire N__3209;
    wire N__3206;
    wire N__3203;
    wire N__3200;
    wire N__3197;
    wire N__3194;
    wire N__3191;
    wire N__3188;
    wire N__3185;
    wire N__3182;
    wire N__3181;
    wire N__3178;
    wire N__3175;
    wire N__3170;
    wire N__3169;
    wire N__3166;
    wire N__3163;
    wire N__3158;
    wire N__3155;
    wire N__3152;
    wire N__3149;
    wire N__3146;
    wire N__3143;
    wire N__3140;
    wire N__3137;
    wire N__3134;
    wire N__3131;
    wire N__3128;
    wire N__3125;
    wire N__3122;
    wire N__3119;
    wire N__3116;
    wire N__3113;
    wire N__3110;
    wire N__3107;
    wire N__3106;
    wire N__3103;
    wire N__3100;
    wire N__3097;
    wire N__3092;
    wire N__3091;
    wire N__3088;
    wire N__3085;
    wire N__3080;
    wire N__3079;
    wire N__3076;
    wire N__3073;
    wire N__3070;
    wire N__3065;
    wire N__3064;
    wire N__3063;
    wire N__3060;
    wire N__3055;
    wire N__3050;
    wire N__3049;
    wire N__3046;
    wire N__3043;
    wire N__3038;
    wire N__3037;
    wire N__3034;
    wire N__3031;
    wire N__3028;
    wire N__3023;
    wire N__3022;
    wire N__3019;
    wire N__3016;
    wire N__3013;
    wire N__3008;
    wire N__3007;
    wire N__3004;
    wire N__3001;
    wire N__3000;
    wire N__2999;
    wire N__2996;
    wire N__2989;
    wire N__2984;
    wire N__2981;
    wire N__2980;
    wire N__2977;
    wire N__2974;
    wire N__2971;
    wire N__2966;
    wire N__2963;
    wire N__2960;
    wire N__2957;
    wire N__2954;
    wire N__2951;
    wire N__2948;
    wire N__2945;
    wire N__2942;
    wire N__2939;
    wire N__2936;
    wire N__2933;
    wire N__2930;
    wire N__2927;
    wire N__2924;
    wire N__2921;
    wire N__2920;
    wire N__2917;
    wire N__2914;
    wire N__2909;
    wire N__2906;
    wire N__2903;
    wire N__2900;
    wire N__2897;
    wire N__2894;
    wire N__2891;
    wire N__2888;
    wire N__2885;
    wire N__2882;
    wire N__2879;
    wire N__2876;
    wire N__2873;
    wire N__2870;
    wire N__2867;
    wire N__2864;
    wire N__2861;
    wire N__2858;
    wire N__2855;
    wire N__2852;
    wire N__2849;
    wire N__2846;
    wire N__2843;
    wire N__2840;
    wire N__2837;
    wire N__2834;
    wire N__2831;
    wire N__2828;
    wire N__2825;
    wire N__2822;
    wire N__2819;
    wire N__2816;
    wire N__2813;
    wire N__2810;
    wire N__2807;
    wire N__2804;
    wire N__2801;
    wire N__2798;
    wire N__2795;
    wire N__2792;
    wire N__2789;
    wire N__2786;
    wire N__2783;
    wire N__2780;
    wire N__2777;
    wire N__2774;
    wire N__2771;
    wire N__2768;
    wire N__2765;
    wire N__2762;
    wire N__2759;
    wire N__2756;
    wire N__2753;
    wire N__2750;
    wire N__2747;
    wire N__2744;
    wire N__2741;
    wire N__2740;
    wire N__2737;
    wire N__2734;
    wire N__2729;
    wire N__2728;
    wire N__2725;
    wire N__2722;
    wire N__2717;
    wire N__2716;
    wire N__2713;
    wire N__2710;
    wire N__2707;
    wire N__2702;
    wire N__2701;
    wire N__2698;
    wire N__2695;
    wire N__2690;
    wire N__2687;
    wire N__2684;
    wire N__2681;
    wire N__2680;
    wire N__2677;
    wire N__2674;
    wire N__2669;
    wire N__2666;
    wire N__2663;
    wire N__2660;
    wire N__2657;
    wire N__2654;
    wire N__2651;
    wire N__2648;
    wire N__2645;
    wire N__2642;
    wire N__2639;
    wire N__2636;
    wire N__2633;
    wire N__2630;
    wire N__2627;
    wire N__2624;
    wire N__2621;
    wire N__2618;
    wire N__2615;
    wire N__2612;
    wire N__2609;
    wire N__2606;
    wire N__2603;
    wire N__2600;
    wire N__2597;
    wire N__2594;
    wire N__2591;
    wire N__2588;
    wire N__2585;
    wire N__2582;
    wire CLK40_ibuf_gb_io_gb_input;
    wire GNDG0;
    wire VCCG0;
    wire RESETn_c_i;
    wire CONSTANT_ONE_NET;
    wire A_c_27;
    wire A_c_28;
    wire \INVU400_SDRAM.SDRAM_CONFIGUREDC_net ;
    wire \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_a2_1_0_0_cascade_ ;
    wire bfn_4_5_0_;
    wire \U400_SDRAM.un2_REFRESH_COUNTER_cry_1 ;
    wire \U400_SDRAM.un2_REFRESH_COUNTER_cry_2 ;
    wire \U400_SDRAM.un2_REFRESH_COUNTER_cry_3 ;
    wire \U400_SDRAM.un2_REFRESH_COUNTER_cry_4 ;
    wire \U400_SDRAM.un2_REFRESH_COUNTER_cry_5 ;
    wire \U400_SDRAM.un2_REFRESH_COUNTER_cry_6 ;
    wire \U400_SDRAM.un2_REFRESH_COUNTER_cry_7 ;
    wire \INVU400_SDRAM.REFRESH_COUNTER_2C_net ;
    wire bfn_4_6_0_;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_0 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_1 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_2 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_3 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_4 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_5 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_6 ;
    wire \INVU400_SDRAM.SDRAM_COUNTER_2C_net ;
    wire \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_0_0 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_a2_1_0_cascade_ ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U400_SDRAM.N_97_cascade_ ;
    wire \U400_SDRAM.N_256_cascade_ ;
    wire \U400_SDRAM.SDRAM_CMD_3_sqmuxa ;
    wire CS0n_c;
    wire \INVU400_SDRAM.CS0nC_net ;
    wire CASn_c;
    wire WEn_c;
    wire \INVU400_SDRAM.CASnC_net ;
    wire RASn_c;
    wire \INVU400_SDRAM.RASnC_net ;
    wire A_c_24;
    wire A_c_18;
    wire MA_c_8;
    wire A_c_9;
    wire A_c_17;
    wire MA_c_7;
    wire \INVU400_SDRAM.MA_nesr_8C_net ;
    wire A_c_8;
    wire A_c_16;
    wire MA_c_6;
    wire \INVU400_SDRAM.MA_nesr_6C_net ;
    wire \U400_SDRAM.N_216 ;
    wire \U400_SDRAM.N_187 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_2_0 ;
    wire \U400_SDRAM.SDRAM_COUNTER_s_0 ;
    wire \INVU400_SDRAM.SDRAM_COUNTER_0C_net ;
    wire \U400_SDRAM.TACK_7_iv_i_i_2 ;
    wire \U400_SDRAM.TACK_7_iv_i_i_1_0_cascade_ ;
    wire \U400_SDRAM.N_258 ;
    wire \U400_SDRAM.un1_SDRAM_COUNTER52_4_i_0_1 ;
    wire \U400_SDRAM.N_258_cascade_ ;
    wire \U400_SDRAM.un1_SDRAM_COUNTER52_4_i_0_0 ;
    wire \U400_SDRAM.N_240_cascade_ ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_2 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_0 ;
    wire \INVU400_SDRAM.REFRESH_COUNTER_1C_net ;
    wire \U400_SDRAM.SDRAM_CONFIGURED_RNIJKCAZ0Z2 ;
    wire \U400_SDRAM.CS0_EN_0_cascade_ ;
    wire \U400_SDRAM.CS0_ENZ0 ;
    wire A_c_23;
    wire \U400_SDRAM.CS1_EN_0_cascade_ ;
    wire \INVU400_SDRAM.CS0_ENC_net ;
    wire \U400_SDRAM.N_114_cascade_ ;
    wire \U400_SDRAM.N_220 ;
    wire \U400_SDRAM.SDRAM_CONFIGURED_RNI5POA3Z0Z_0 ;
    wire \U400_SDRAM.N_230_cascade_ ;
    wire A_c_19;
    wire MA_c_9;
    wire \INVU400_SDRAM.MA_nesr_9C_net ;
    wire A_c_30;
    wire A_c_29;
    wire \U400_SDRAM.TA_COUNTER_0_sqmuxa_cascade_ ;
    wire \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en ;
    wire \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en_0 ;
    wire A_c_21;
    wire BANK0_c;
    wire A_c_22;
    wire \U400_SDRAM.N_240 ;
    wire BANK1_c;
    wire RnW_c;
    wire \U400_SDRAM.N_82 ;
    wire \U400_SDRAM.N_34 ;
    wire \INVU400_SDRAM.BANK0C_net ;
    wire \U400_SDRAM.N_118_cascade_ ;
    wire \U400_SDRAM.N_215 ;
    wire \U400_SDRAM.RAM_CYCLEZ0 ;
    wire \U400_SDRAM.N_236_cascade_ ;
    wire \U400_SDRAM.N_23_i ;
    wire \U400_SDRAM.N_23_i_cascade_ ;
    wire \U400_SDRAM.N_242 ;
    wire \U400_SDRAM.N_139 ;
    wire \U400_SDRAM.SDRAM_COUNTER_s_1 ;
    wire \U400_SDRAM.N_198 ;
    wire \U400_SDRAM.N_259 ;
    wire \U400_SDRAM.N_118 ;
    wire \U400_SDRAM.N_39 ;
    wire \U400_SDRAM.SDRAM_COUNTER_s_3 ;
    wire \INVU400_SDRAM.SDRAM_COUNTER_1C_net ;
    wire \U400_SDRAM.N_219_i ;
    wire \U400_SDRAM.N_239 ;
    wire \U400_SDRAM.N_207 ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_5_1_cascade_ ;
    wire \U400_SDRAM.N_250 ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_0_31_i_i_i_2_cascade_ ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_0_31_i_i_i_3_cascade_ ;
    wire \INVU400_SDRAM.SDRAM_CMD_1C_net ;
    wire \U400_SDRAM.N_261 ;
    wire \U400_SDRAM.N_140 ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_4_1 ;
    wire \U400_SDRAM.CS1_ENZ0 ;
    wire CS1n_c;
    wire \INVU400_SDRAM.CS1nC_net ;
    wire A_c_26;
    wire MA_c_12;
    wire \INVU400_SDRAM.MA_nesr_12C_net ;
    wire TA_OUT;
    wire N_66;
    wire \U400_SDRAM.BURSTZ0 ;
    wire \U400_SDRAM.TA_EN11_m ;
    wire \U400_SDRAM.un1_TA_COUNTER26_0_cascade_ ;
    wire \U400_SDRAM.un1_TA_COUNTER26_2_0 ;
    wire \U400_SDRAM.TA_COUNTER27 ;
    wire \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0 ;
    wire \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0_cascade_ ;
    wire \U400_SDRAM.TA_COUNTERZ0Z_2 ;
    wire \U400_SDRAM.TA_COUNTERZ0Z_3 ;
    wire \U400_SDRAM.TA_COUNTERZ0Z_1 ;
    wire \U400_SDRAM.CO1 ;
    wire \U400_SDRAM.TA_COUNTER23 ;
    wire \U400_SDRAM.TACKZ0 ;
    wire \U400_SDRAM.TA_COUNTER_7_f1_0_0_cascade_ ;
    wire \U400_SDRAM.TA_COUNTER_0_sqmuxa ;
    wire \U400_SDRAM.TA_COUNTERZ0Z_0 ;
    wire CLK40_c_g;
    wire \U400_SDRAM.N_189 ;
    wire RESETn_c;
    wire \U400_SDRAM.un1_REFRESH_COUNTERlto7_5 ;
    wire \U400_SDRAM.un1_REFRESH_COUNTERlto7_4 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_8 ;
    wire \U400_SDRAM.un1_SDRAM_COUNTER52_2_0_i_1 ;
    wire \U400_SDRAM.N_195_cascade_ ;
    wire \U400_SDRAM.N_94 ;
    wire U400_ADDRESS_DECODE_RAM_SPACE_i_o3_0_o2_1;
    wire A_c_31;
    wire U400_ADDRESS_DECODE_RAM_SPACE_i_o3_0_o2_2;
    wire TSn_c;
    wire \U400_SDRAM.N_225 ;
    wire \U400_SDRAM.N_236 ;
    wire \U400_SDRAM.RAM_CYCLE_STARTZ0 ;
    wire \U400_SDRAM.N_228 ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_a2_2_0_1_cascade_ ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_1_1_cascade_ ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_2_1 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U400_SDRAM.WRITE_CYCLEZ0 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U400_SDRAM.N_256 ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_a2_0_1_0_cascade_ ;
    wire \U400_SDRAM.N_97 ;
    wire \U400_SDRAM.SDRAM_CONFIGUREDZ0 ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_0_0 ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_1_0_cascade_ ;
    wire \U400_SDRAM.N_114 ;
    wire \INVU400_SDRAM.SDRAM_CMD_ne_0C_net ;
    wire \U400_SDRAM.N_71 ;
    wire A_c_25;
    wire MA_c_11;
    wire \INVU400_SDRAM.MA_nesr_11C_net ;
    wire A_c_7;
    wire A_c_15;
    wire \U400_SDRAM.MA_5_iv_0_5 ;
    wire MA_c_5;
    wire \INVU400_SDRAM.MA_nesr_5C_net ;
    wire \U400_BYTE_ENABLE.N_101_i ;
    wire \U400_BYTE_ENABLE.N_101_i_cascade_ ;
    wire un1_LMBEn_i_0_0;
    wire A_c_0;
    wire RAM_SPACE_i_o3_0_o2dup;
    wire A_c_20;
    wire MA_c_10;
    wire \INVU400_SDRAM.MA_nesr_10C_net ;
    wire \U400_SDRAM.SDRAM_CMDZ0Z_1 ;
    wire A_c_3;
    wire \U400_SDRAM.SDRAM_CMDZ0Z_0 ;
    wire N_63;
    wire A_c_1;
    wire SIZ_c_1;
    wire \U400_BYTE_ENABLE.N_168 ;
    wire SIZ_c_0;
    wire un1_LLBEn_i_0_0;
    wire TA_EN_i_ess;
    wire N_526_i;
    wire A_c_5;
    wire A_c_13;
    wire MA_c_3;
    wire \INVU400_SDRAM.MA_nesr_3C_net ;
    wire A_c_4;
    wire A_c_12;
    wire MA_c_2;
    wire A_c_2;
    wire A_c_10;
    wire MA_c_0;
    wire A_c_6;
    wire A_c_14;
    wire \U400_SDRAM.SDRAM_CMDZ0Z_2 ;
    wire MA_c_4;
    wire \U400_SDRAM.MA_5_iv_0_1 ;
    wire A_c_11;
    wire \U400_SDRAM.MA19 ;
    wire MA_c_1;
    wire _gnd_net_;
    wire \INVU400_SDRAM.MA_nesr_2C_net ;
    wire \U400_SDRAM.un1_MA20_0_i_0 ;
    wire RESETn_c_i_g;

    IO_PAD MA_obuf_7_iopad (
            .OE(N__7125),
            .DIN(N__7124),
            .DOUT(N__7123),
            .PACKAGEPIN(MA[7]));
    defparam MA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_7_preio (
            .PADOEN(N__7125),
            .PADOUT(N__7124),
            .PADIN(N__7123),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2774),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__7116),
            .DIN(N__7115),
            .DOUT(N__7114),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__7116),
            .PADOUT(N__7115),
            .PADIN(N__7114),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__7107),
            .DIN(N__7106),
            .DOUT(N__7105),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__7107),
            .PADOUT(N__7106),
            .PADIN(N__7105),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2870),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__7098),
            .DIN(N__7097),
            .DOUT(N__7096),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__7098),
            .PADOUT(N__7097),
            .PADIN(N__7096),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3329),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_8_iopad (
            .OE(N__7089),
            .DIN(N__7088),
            .DOUT(N__7087),
            .PACKAGEPIN(MA[8]));
    defparam MA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_8_preio (
            .PADOEN(N__7089),
            .PADOUT(N__7088),
            .PADIN(N__7087),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2810),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_10_iopad (
            .OE(N__7080),
            .DIN(N__7079),
            .DOUT(N__7078),
            .PACKAGEPIN(MA[10]));
    defparam MA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_10_preio (
            .PADOEN(N__7080),
            .PADOUT(N__7079),
            .PADIN(N__7078),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6086),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_23_iopad (
            .OE(N__7071),
            .DIN(N__7070),
            .DOUT(N__7069),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__7071),
            .PADOUT(N__7070),
            .PADIN(N__7069),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_2_iopad (
            .OE(N__7062),
            .DIN(N__7061),
            .DOUT(N__7060),
            .PACKAGEPIN(MA[2]));
    defparam MA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_2_preio (
            .PADOEN(N__7062),
            .PADOUT(N__7061),
            .PADIN(N__7060),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5597),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__7053),
            .DIN(N__7052),
            .DOUT(N__7051),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__7053),
            .PADOUT(N__7052),
            .PADIN(N__7051),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__7044),
            .DIN(N__7043),
            .DOUT(N__7042),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__7044),
            .PADOUT(N__7043),
            .PADIN(N__7042),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__7035),
            .DIN(N__7034),
            .DOUT(N__7033),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__7035),
            .PADOUT(N__7034),
            .PADIN(N__7033),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3752),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_24_iopad (
            .OE(N__7026),
            .DIN(N__7025),
            .DOUT(N__7024),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__7026),
            .PADOUT(N__7025),
            .PADIN(N__7024),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_31_iopad (
            .OE(N__7017),
            .DIN(N__7016),
            .DOUT(N__7015),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__7017),
            .PADOUT(N__7016),
            .PADIN(N__7015),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__7008),
            .DIN(N__7007),
            .DOUT(N__7006),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__7008),
            .PADOUT(N__7007),
            .PADIN(N__7006),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_12_iopad (
            .OE(N__6999),
            .DIN(N__6998),
            .DOUT(N__6997),
            .PACKAGEPIN(MA[12]));
    defparam MA_obuf_12_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_12_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_12_preio (
            .PADOEN(N__6999),
            .PADOUT(N__6998),
            .PADIN(N__6997),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3584),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_1_iopad (
            .OE(N__6990),
            .DIN(N__6989),
            .DOUT(N__6988),
            .PACKAGEPIN(MA[1]));
    defparam MA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_1_preio (
            .PADOEN(N__6990),
            .PADOUT(N__6989),
            .PADIN(N__6988),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6278),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__6981),
            .DIN(N__6980),
            .DOUT(N__6979),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__6981),
            .PADOUT(N__6980),
            .PADIN(N__6979),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__6972),
            .DIN(N__6971),
            .DOUT(N__6970),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__6972),
            .PADOUT(N__6971),
            .PADIN(N__6970),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_21_iopad (
            .OE(N__6963),
            .DIN(N__6962),
            .DOUT(N__6961),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__6963),
            .PADOUT(N__6962),
            .PADIN(N__6961),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_4_iopad (
            .OE(N__6954),
            .DIN(N__6953),
            .DOUT(N__6952),
            .PACKAGEPIN(MA[4]));
    defparam MA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_4_preio (
            .PADOEN(N__6954),
            .PADOUT(N__6953),
            .PADIN(N__6952),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6368),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__6945),
            .DIN(N__6944),
            .DOUT(N__6943),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__6945),
            .PADOUT(N__6944),
            .PADIN(N__6943),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__6936),
            .DIN(N__6935),
            .DOUT(N__6934),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__6936),
            .PADOUT(N__6935),
            .PADIN(N__6934),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__6927),
            .DIN(N__6926),
            .DOUT(N__6925),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__6927),
            .PADOUT(N__6926),
            .PADIN(N__6925),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5696),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__6918),
            .DIN(N__6917),
            .DOUT(N__6916),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__6918),
            .PADOUT(N__6917),
            .PADIN(N__6916),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_9_iopad (
            .OE(N__6909),
            .DIN(N__6908),
            .DOUT(N__6907),
            .PACKAGEPIN(MA[9]));
    defparam MA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_9_preio (
            .PADOEN(N__6909),
            .PADOUT(N__6908),
            .PADIN(N__6907),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3227),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__6900),
            .DIN(N__6899),
            .DOUT(N__6898),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__6900),
            .PADOUT(N__6899),
            .PADIN(N__6898),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5876),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__6891),
            .DIN(N__6890),
            .DOUT(N__6889),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__6891),
            .PADOUT(N__6890),
            .PADIN(N__6889),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_29_iopad (
            .OE(N__6882),
            .DIN(N__6881),
            .DOUT(N__6880),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__6882),
            .PADOUT(N__6881),
            .PADIN(N__6880),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__6873),
            .DIN(N__6872),
            .DOUT(N__6871),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__6873),
            .PADOUT(N__6872),
            .PADIN(N__6871),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2636),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__6864),
            .DIN(N__6863),
            .DOUT(N__6862),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__6864),
            .PADOUT(N__6863),
            .PADIN(N__6862),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_22_iopad (
            .OE(N__6855),
            .DIN(N__6854),
            .DOUT(N__6853),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__6855),
            .PADOUT(N__6854),
            .PADIN(N__6853),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_3_iopad (
            .OE(N__6846),
            .DIN(N__6845),
            .DOUT(N__6844),
            .PACKAGEPIN(MA[3]));
    defparam MA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_3_preio (
            .PADOEN(N__6846),
            .PADOUT(N__6845),
            .PADIN(N__6844),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5639),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__6837),
            .DIN(N__6836),
            .DOUT(N__6835),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__6837),
            .PADOUT(N__6836),
            .PADIN(N__6835),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__6828),
            .DIN(N__6827),
            .DOUT(N__6826),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__6828),
            .PADOUT(N__6827),
            .PADIN(N__6826),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_27_iopad (
            .OE(N__6819),
            .DIN(N__6818),
            .DOUT(N__6817),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__6819),
            .PADOUT(N__6818),
            .PADIN(N__6817),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_6_iopad (
            .OE(N__6810),
            .DIN(N__6809),
            .DOUT(N__6808),
            .PACKAGEPIN(MA[6]));
    defparam MA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_6_preio (
            .PADOEN(N__6810),
            .PADOUT(N__6809),
            .PADIN(N__6808),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2939),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__6801),
            .DIN(N__6800),
            .DOUT(N__6799),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__6801),
            .PADOUT(N__6800),
            .PADIN(N__6799),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__6792),
            .DIN(N__6791),
            .DOUT(N__6790),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__6792),
            .PADOUT(N__6791),
            .PADIN(N__6790),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__6783),
            .DIN(N__6782),
            .DOUT(N__6781),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__6783),
            .PADOUT(N__6782),
            .PADIN(N__6781),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__6774),
            .DIN(N__6773),
            .DOUT(N__6772),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__6774),
            .PADOUT(N__6773),
            .PADIN(N__6772),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2852),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__6765),
            .DIN(N__6764),
            .DOUT(N__6763),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__6765),
            .PADOUT(N__6764),
            .PADIN(N__6763),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__6756),
            .DIN(N__6755),
            .DOUT(N__6754),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__6756),
            .PADOUT(N__6755),
            .PADIN(N__6754),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3380),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_11_iopad (
            .OE(N__6747),
            .DIN(N__6746),
            .DOUT(N__6745),
            .PACKAGEPIN(MA[11]));
    defparam MA_obuf_11_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_11_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_11_preio (
            .PADOEN(N__6747),
            .PADOUT(N__6746),
            .PADIN(N__6745),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5321),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TAn_obuft_iopad (
            .OE(N__6738),
            .DIN(N__6737),
            .DOUT(N__6736),
            .PACKAGEPIN(TAn));
    defparam TAn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TAn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TAn_obuft_preio (
            .PADOEN(N__6738),
            .PADOUT(N__6737),
            .PADIN(N__6736),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5672),
            .DIN0(),
            .DOUT0(N__3773),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__6729),
            .DIN(N__6728),
            .DOUT(N__6727),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__6729),
            .PADOUT(N__6728),
            .PADIN(N__6727),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_5_iopad (
            .OE(N__6720),
            .DIN(N__6719),
            .DOUT(N__6718),
            .PACKAGEPIN(MA[5]));
    defparam MA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_5_preio (
            .PADOEN(N__6720),
            .PADOUT(N__6719),
            .PADIN(N__6718),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5282),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__6711),
            .DIN(N__6710),
            .DOUT(N__6709),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__6711),
            .PADOUT(N__6710),
            .PADIN(N__6709),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__6702),
            .DIN(N__6701),
            .DOUT(N__6700),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__6702),
            .PADOUT(N__6701),
            .PADIN(N__6700),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam LBENn_obuf_iopad.PULLUP=1'b1;
    IO_PAD LBENn_obuf_iopad (
            .OE(N__6693),
            .DIN(N__6692),
            .DOUT(N__6691),
            .PACKAGEPIN(LBENn));
    defparam LBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LBENn_obuf_preio (
            .PADOEN(N__6693),
            .PADOUT(N__6692),
            .PADIN(N__6691),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5194),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_25_iopad (
            .OE(N__6684),
            .DIN(N__6683),
            .DOUT(N__6682),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__6684),
            .PADOUT(N__6683),
            .PADIN(N__6682),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CS1n_obuf_iopad (
            .OE(N__6675),
            .DIN(N__6674),
            .DOUT(N__6673),
            .PACKAGEPIN(CS1n));
    defparam CS1n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CS1n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CS1n_obuf_preio (
            .PADOEN(N__6675),
            .PADOUT(N__6674),
            .PADIN(N__6673),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3614),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__6666),
            .DIN(N__6665),
            .DOUT(N__6664),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__6666),
            .PADOUT(N__6665),
            .PADIN(N__6664),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_28_iopad (
            .OE(N__6657),
            .DIN(N__6656),
            .DOUT(N__6655),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__6657),
            .PADOUT(N__6656),
            .PADIN(N__6655),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_30_iopad (
            .OE(N__6648),
            .DIN(N__6647),
            .DOUT(N__6646),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__6648),
            .PADOUT(N__6647),
            .PADIN(N__6646),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__6639),
            .DIN(N__6638),
            .DOUT(N__6637),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__6639),
            .PADOUT(N__6638),
            .PADIN(N__6637),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__6630),
            .DIN(N__6629),
            .DOUT(N__6628),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__6630),
            .PADOUT(N__6629),
            .PADIN(N__6628),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2861),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_0_iopad (
            .OE(N__6621),
            .DIN(N__6620),
            .DOUT(N__6619),
            .PACKAGEPIN(MA[0]));
    defparam MA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_0_preio (
            .PADOEN(N__6621),
            .PADOUT(N__6620),
            .PADIN(N__6619),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5564),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__6612),
            .DIN(N__6611),
            .DOUT(N__6610),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__6612),
            .PADOUT(N__6611),
            .PADIN(N__6610),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__6603),
            .DIN(N__6602),
            .DOUT(N__6601),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__6603),
            .PADOUT(N__6602),
            .PADIN(N__6601),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__6594),
            .DIN(N__6593),
            .DOUT(N__6592),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__6594),
            .PADOUT(N__6593),
            .PADIN(N__6592),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CS0n_obuf_iopad (
            .OE(N__6585),
            .DIN(N__6584),
            .DOUT(N__6583),
            .PACKAGEPIN(CS0n));
    defparam CS0n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CS0n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CS0n_obuf_preio (
            .PADOEN(N__6585),
            .PADOUT(N__6584),
            .PADIN(N__6583),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2882),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_26_iopad (
            .OE(N__6576),
            .DIN(N__6575),
            .DOUT(N__6574),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__6576),
            .PADOUT(N__6575),
            .PADIN(N__6574),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__6567),
            .DIN(N__6566),
            .DOUT(N__6565),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__6567),
            .PADOUT(N__6566),
            .PADIN(N__6565),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5258),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__6558),
            .DIN(N__6557),
            .DOUT(N__6556),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__6558),
            .PADOUT(N__6557),
            .PADIN(N__6556),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_ibuf_gb_io_iopad (
            .OE(N__6549),
            .DIN(N__6548),
            .DOUT(N__6547),
            .PACKAGEPIN(CLK40));
    defparam CLK40_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_ibuf_gb_io_preio (
            .PADOEN(N__6549),
            .PADOUT(N__6548),
            .PADIN(N__6547),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1554 (
            .O(N__6530),
            .I(N__6527));
    LocalMux I__1553 (
            .O(N__6527),
            .I(N__6524));
    Span4Mux_s3_v I__1552 (
            .O(N__6524),
            .I(N__6521));
    Odrv4 I__1551 (
            .O(N__6521),
            .I(A_c_6));
    CascadeMux I__1550 (
            .O(N__6518),
            .I(N__6515));
    InMux I__1549 (
            .O(N__6515),
            .I(N__6512));
    LocalMux I__1548 (
            .O(N__6512),
            .I(N__6509));
    IoSpan4Mux I__1547 (
            .O(N__6509),
            .I(N__6506));
    Odrv4 I__1546 (
            .O(N__6506),
            .I(A_c_14));
    InMux I__1545 (
            .O(N__6503),
            .I(N__6492));
    InMux I__1544 (
            .O(N__6502),
            .I(N__6486));
    InMux I__1543 (
            .O(N__6501),
            .I(N__6482));
    InMux I__1542 (
            .O(N__6500),
            .I(N__6479));
    InMux I__1541 (
            .O(N__6499),
            .I(N__6476));
    InMux I__1540 (
            .O(N__6498),
            .I(N__6469));
    InMux I__1539 (
            .O(N__6497),
            .I(N__6469));
    InMux I__1538 (
            .O(N__6496),
            .I(N__6466));
    InMux I__1537 (
            .O(N__6495),
            .I(N__6463));
    LocalMux I__1536 (
            .O(N__6492),
            .I(N__6459));
    InMux I__1535 (
            .O(N__6491),
            .I(N__6454));
    InMux I__1534 (
            .O(N__6490),
            .I(N__6454));
    InMux I__1533 (
            .O(N__6489),
            .I(N__6451));
    LocalMux I__1532 (
            .O(N__6486),
            .I(N__6447));
    InMux I__1531 (
            .O(N__6485),
            .I(N__6444));
    LocalMux I__1530 (
            .O(N__6482),
            .I(N__6437));
    LocalMux I__1529 (
            .O(N__6479),
            .I(N__6437));
    LocalMux I__1528 (
            .O(N__6476),
            .I(N__6437));
    InMux I__1527 (
            .O(N__6475),
            .I(N__6432));
    InMux I__1526 (
            .O(N__6474),
            .I(N__6432));
    LocalMux I__1525 (
            .O(N__6469),
            .I(N__6427));
    LocalMux I__1524 (
            .O(N__6466),
            .I(N__6427));
    LocalMux I__1523 (
            .O(N__6463),
            .I(N__6422));
    InMux I__1522 (
            .O(N__6462),
            .I(N__6419));
    Span4Mux_v I__1521 (
            .O(N__6459),
            .I(N__6412));
    LocalMux I__1520 (
            .O(N__6454),
            .I(N__6412));
    LocalMux I__1519 (
            .O(N__6451),
            .I(N__6412));
    InMux I__1518 (
            .O(N__6450),
            .I(N__6409));
    Span4Mux_h I__1517 (
            .O(N__6447),
            .I(N__6400));
    LocalMux I__1516 (
            .O(N__6444),
            .I(N__6400));
    Span4Mux_v I__1515 (
            .O(N__6437),
            .I(N__6400));
    LocalMux I__1514 (
            .O(N__6432),
            .I(N__6400));
    Span12Mux_s8_v I__1513 (
            .O(N__6427),
            .I(N__6397));
    InMux I__1512 (
            .O(N__6426),
            .I(N__6394));
    InMux I__1511 (
            .O(N__6425),
            .I(N__6391));
    Span12Mux_s6_h I__1510 (
            .O(N__6422),
            .I(N__6386));
    LocalMux I__1509 (
            .O(N__6419),
            .I(N__6386));
    Span4Mux_v I__1508 (
            .O(N__6412),
            .I(N__6379));
    LocalMux I__1507 (
            .O(N__6409),
            .I(N__6379));
    Span4Mux_v I__1506 (
            .O(N__6400),
            .I(N__6379));
    Odrv12 I__1505 (
            .O(N__6397),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1504 (
            .O(N__6394),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1503 (
            .O(N__6391),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_2 ));
    Odrv12 I__1502 (
            .O(N__6386),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1501 (
            .O(N__6379),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_2 ));
    IoInMux I__1500 (
            .O(N__6368),
            .I(N__6365));
    LocalMux I__1499 (
            .O(N__6365),
            .I(N__6362));
    Span4Mux_s1_v I__1498 (
            .O(N__6362),
            .I(N__6359));
    Span4Mux_h I__1497 (
            .O(N__6359),
            .I(N__6356));
    Odrv4 I__1496 (
            .O(N__6356),
            .I(MA_c_4));
    InMux I__1495 (
            .O(N__6353),
            .I(N__6350));
    LocalMux I__1494 (
            .O(N__6350),
            .I(\U400_SDRAM.MA_5_iv_0_1 ));
    InMux I__1493 (
            .O(N__6347),
            .I(N__6344));
    LocalMux I__1492 (
            .O(N__6344),
            .I(N__6341));
    Odrv4 I__1491 (
            .O(N__6341),
            .I(A_c_11));
    InMux I__1490 (
            .O(N__6338),
            .I(N__6328));
    InMux I__1489 (
            .O(N__6337),
            .I(N__6325));
    InMux I__1488 (
            .O(N__6336),
            .I(N__6316));
    InMux I__1487 (
            .O(N__6335),
            .I(N__6316));
    InMux I__1486 (
            .O(N__6334),
            .I(N__6316));
    InMux I__1485 (
            .O(N__6333),
            .I(N__6316));
    InMux I__1484 (
            .O(N__6332),
            .I(N__6311));
    InMux I__1483 (
            .O(N__6331),
            .I(N__6311));
    LocalMux I__1482 (
            .O(N__6328),
            .I(N__6307));
    LocalMux I__1481 (
            .O(N__6325),
            .I(N__6304));
    LocalMux I__1480 (
            .O(N__6316),
            .I(N__6301));
    LocalMux I__1479 (
            .O(N__6311),
            .I(N__6298));
    InMux I__1478 (
            .O(N__6310),
            .I(N__6295));
    Span4Mux_h I__1477 (
            .O(N__6307),
            .I(N__6290));
    Span4Mux_s2_v I__1476 (
            .O(N__6304),
            .I(N__6290));
    Span4Mux_s2_v I__1475 (
            .O(N__6301),
            .I(N__6287));
    Odrv12 I__1474 (
            .O(N__6298),
            .I(\U400_SDRAM.MA19 ));
    LocalMux I__1473 (
            .O(N__6295),
            .I(\U400_SDRAM.MA19 ));
    Odrv4 I__1472 (
            .O(N__6290),
            .I(\U400_SDRAM.MA19 ));
    Odrv4 I__1471 (
            .O(N__6287),
            .I(\U400_SDRAM.MA19 ));
    IoInMux I__1470 (
            .O(N__6278),
            .I(N__6275));
    LocalMux I__1469 (
            .O(N__6275),
            .I(N__6272));
    Odrv4 I__1468 (
            .O(N__6272),
            .I(MA_c_1));
    CEMux I__1467 (
            .O(N__6269),
            .I(N__6262));
    CEMux I__1466 (
            .O(N__6268),
            .I(N__6259));
    CEMux I__1465 (
            .O(N__6267),
            .I(N__6255));
    CEMux I__1464 (
            .O(N__6266),
            .I(N__6251));
    CEMux I__1463 (
            .O(N__6265),
            .I(N__6248));
    LocalMux I__1462 (
            .O(N__6262),
            .I(N__6245));
    LocalMux I__1461 (
            .O(N__6259),
            .I(N__6242));
    CEMux I__1460 (
            .O(N__6258),
            .I(N__6238));
    LocalMux I__1459 (
            .O(N__6255),
            .I(N__6234));
    CEMux I__1458 (
            .O(N__6254),
            .I(N__6231));
    LocalMux I__1457 (
            .O(N__6251),
            .I(N__6228));
    LocalMux I__1456 (
            .O(N__6248),
            .I(N__6225));
    Span4Mux_v I__1455 (
            .O(N__6245),
            .I(N__6220));
    Span4Mux_h I__1454 (
            .O(N__6242),
            .I(N__6220));
    CEMux I__1453 (
            .O(N__6241),
            .I(N__6217));
    LocalMux I__1452 (
            .O(N__6238),
            .I(N__6214));
    CEMux I__1451 (
            .O(N__6237),
            .I(N__6211));
    Span4Mux_h I__1450 (
            .O(N__6234),
            .I(N__6206));
    LocalMux I__1449 (
            .O(N__6231),
            .I(N__6206));
    Odrv4 I__1448 (
            .O(N__6228),
            .I(\U400_SDRAM.un1_MA20_0_i_0 ));
    Odrv4 I__1447 (
            .O(N__6225),
            .I(\U400_SDRAM.un1_MA20_0_i_0 ));
    Odrv4 I__1446 (
            .O(N__6220),
            .I(\U400_SDRAM.un1_MA20_0_i_0 ));
    LocalMux I__1445 (
            .O(N__6217),
            .I(\U400_SDRAM.un1_MA20_0_i_0 ));
    Odrv12 I__1444 (
            .O(N__6214),
            .I(\U400_SDRAM.un1_MA20_0_i_0 ));
    LocalMux I__1443 (
            .O(N__6211),
            .I(\U400_SDRAM.un1_MA20_0_i_0 ));
    Odrv4 I__1442 (
            .O(N__6206),
            .I(\U400_SDRAM.un1_MA20_0_i_0 ));
    CascadeMux I__1441 (
            .O(N__6191),
            .I(N__6188));
    InMux I__1440 (
            .O(N__6188),
            .I(N__6184));
    InMux I__1439 (
            .O(N__6187),
            .I(N__6181));
    LocalMux I__1438 (
            .O(N__6184),
            .I(N__6174));
    LocalMux I__1437 (
            .O(N__6181),
            .I(N__6166));
    SRMux I__1436 (
            .O(N__6180),
            .I(N__6116));
    SRMux I__1435 (
            .O(N__6179),
            .I(N__6116));
    SRMux I__1434 (
            .O(N__6178),
            .I(N__6116));
    SRMux I__1433 (
            .O(N__6177),
            .I(N__6116));
    Glb2LocalMux I__1432 (
            .O(N__6174),
            .I(N__6116));
    SRMux I__1431 (
            .O(N__6173),
            .I(N__6116));
    SRMux I__1430 (
            .O(N__6172),
            .I(N__6116));
    SRMux I__1429 (
            .O(N__6171),
            .I(N__6116));
    SRMux I__1428 (
            .O(N__6170),
            .I(N__6116));
    SRMux I__1427 (
            .O(N__6169),
            .I(N__6116));
    Glb2LocalMux I__1426 (
            .O(N__6166),
            .I(N__6116));
    SRMux I__1425 (
            .O(N__6165),
            .I(N__6116));
    SRMux I__1424 (
            .O(N__6164),
            .I(N__6116));
    SRMux I__1423 (
            .O(N__6163),
            .I(N__6116));
    SRMux I__1422 (
            .O(N__6162),
            .I(N__6116));
    SRMux I__1421 (
            .O(N__6161),
            .I(N__6116));
    SRMux I__1420 (
            .O(N__6160),
            .I(N__6116));
    SRMux I__1419 (
            .O(N__6159),
            .I(N__6116));
    SRMux I__1418 (
            .O(N__6158),
            .I(N__6116));
    SRMux I__1417 (
            .O(N__6157),
            .I(N__6116));
    GlobalMux I__1416 (
            .O(N__6116),
            .I(N__6113));
    gio2CtrlBuf I__1415 (
            .O(N__6113),
            .I(RESETn_c_i_g));
    CascadeMux I__1414 (
            .O(N__6110),
            .I(N__6107));
    InMux I__1413 (
            .O(N__6107),
            .I(N__6104));
    LocalMux I__1412 (
            .O(N__6104),
            .I(N__6101));
    Span4Mux_v I__1411 (
            .O(N__6101),
            .I(N__6098));
    Span4Mux_v I__1410 (
            .O(N__6098),
            .I(N__6095));
    Span4Mux_v I__1409 (
            .O(N__6095),
            .I(N__6092));
    Sp12to4 I__1408 (
            .O(N__6092),
            .I(N__6089));
    Odrv12 I__1407 (
            .O(N__6089),
            .I(A_c_20));
    IoInMux I__1406 (
            .O(N__6086),
            .I(N__6083));
    LocalMux I__1405 (
            .O(N__6083),
            .I(N__6080));
    Odrv12 I__1404 (
            .O(N__6080),
            .I(MA_c_10));
    InMux I__1403 (
            .O(N__6077),
            .I(N__6071));
    InMux I__1402 (
            .O(N__6076),
            .I(N__6064));
    InMux I__1401 (
            .O(N__6075),
            .I(N__6059));
    InMux I__1400 (
            .O(N__6074),
            .I(N__6056));
    LocalMux I__1399 (
            .O(N__6071),
            .I(N__6053));
    InMux I__1398 (
            .O(N__6070),
            .I(N__6050));
    InMux I__1397 (
            .O(N__6069),
            .I(N__6047));
    InMux I__1396 (
            .O(N__6068),
            .I(N__6044));
    InMux I__1395 (
            .O(N__6067),
            .I(N__6041));
    LocalMux I__1394 (
            .O(N__6064),
            .I(N__6037));
    InMux I__1393 (
            .O(N__6063),
            .I(N__6032));
    InMux I__1392 (
            .O(N__6062),
            .I(N__6032));
    LocalMux I__1391 (
            .O(N__6059),
            .I(N__6022));
    LocalMux I__1390 (
            .O(N__6056),
            .I(N__6022));
    Span4Mux_h I__1389 (
            .O(N__6053),
            .I(N__6022));
    LocalMux I__1388 (
            .O(N__6050),
            .I(N__6022));
    LocalMux I__1387 (
            .O(N__6047),
            .I(N__6017));
    LocalMux I__1386 (
            .O(N__6044),
            .I(N__6017));
    LocalMux I__1385 (
            .O(N__6041),
            .I(N__6014));
    InMux I__1384 (
            .O(N__6040),
            .I(N__6011));
    Span4Mux_v I__1383 (
            .O(N__6037),
            .I(N__6006));
    LocalMux I__1382 (
            .O(N__6032),
            .I(N__6006));
    InMux I__1381 (
            .O(N__6031),
            .I(N__6003));
    Span4Mux_v I__1380 (
            .O(N__6022),
            .I(N__6000));
    Span4Mux_v I__1379 (
            .O(N__6017),
            .I(N__5991));
    Span4Mux_h I__1378 (
            .O(N__6014),
            .I(N__5991));
    LocalMux I__1377 (
            .O(N__6011),
            .I(N__5991));
    Span4Mux_v I__1376 (
            .O(N__6006),
            .I(N__5991));
    LocalMux I__1375 (
            .O(N__6003),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1374 (
            .O(N__6000),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1373 (
            .O(N__5991),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_1 ));
    CascadeMux I__1372 (
            .O(N__5984),
            .I(N__5981));
    InMux I__1371 (
            .O(N__5981),
            .I(N__5978));
    LocalMux I__1370 (
            .O(N__5978),
            .I(N__5975));
    Span4Mux_h I__1369 (
            .O(N__5975),
            .I(N__5972));
    Odrv4 I__1368 (
            .O(N__5972),
            .I(A_c_3));
    CascadeMux I__1367 (
            .O(N__5969),
            .I(N__5964));
    InMux I__1366 (
            .O(N__5968),
            .I(N__5961));
    InMux I__1365 (
            .O(N__5967),
            .I(N__5951));
    InMux I__1364 (
            .O(N__5964),
            .I(N__5948));
    LocalMux I__1363 (
            .O(N__5961),
            .I(N__5945));
    InMux I__1362 (
            .O(N__5960),
            .I(N__5942));
    InMux I__1361 (
            .O(N__5959),
            .I(N__5939));
    InMux I__1360 (
            .O(N__5958),
            .I(N__5936));
    InMux I__1359 (
            .O(N__5957),
            .I(N__5933));
    InMux I__1358 (
            .O(N__5956),
            .I(N__5930));
    InMux I__1357 (
            .O(N__5955),
            .I(N__5925));
    InMux I__1356 (
            .O(N__5954),
            .I(N__5925));
    LocalMux I__1355 (
            .O(N__5951),
            .I(N__5921));
    LocalMux I__1354 (
            .O(N__5948),
            .I(N__5918));
    Span4Mux_h I__1353 (
            .O(N__5945),
            .I(N__5913));
    LocalMux I__1352 (
            .O(N__5942),
            .I(N__5913));
    LocalMux I__1351 (
            .O(N__5939),
            .I(N__5906));
    LocalMux I__1350 (
            .O(N__5936),
            .I(N__5906));
    LocalMux I__1349 (
            .O(N__5933),
            .I(N__5906));
    LocalMux I__1348 (
            .O(N__5930),
            .I(N__5901));
    LocalMux I__1347 (
            .O(N__5925),
            .I(N__5901));
    InMux I__1346 (
            .O(N__5924),
            .I(N__5898));
    Span4Mux_h I__1345 (
            .O(N__5921),
            .I(N__5895));
    Span4Mux_h I__1344 (
            .O(N__5918),
            .I(N__5890));
    Span4Mux_v I__1343 (
            .O(N__5913),
            .I(N__5890));
    Span4Mux_v I__1342 (
            .O(N__5906),
            .I(N__5885));
    Span4Mux_v I__1341 (
            .O(N__5901),
            .I(N__5885));
    LocalMux I__1340 (
            .O(N__5898),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1339 (
            .O(N__5895),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1338 (
            .O(N__5890),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1337 (
            .O(N__5885),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_0 ));
    IoInMux I__1336 (
            .O(N__5876),
            .I(N__5873));
    LocalMux I__1335 (
            .O(N__5873),
            .I(N__5870));
    Odrv4 I__1334 (
            .O(N__5870),
            .I(N_63));
    InMux I__1333 (
            .O(N__5867),
            .I(N__5861));
    InMux I__1332 (
            .O(N__5866),
            .I(N__5861));
    LocalMux I__1331 (
            .O(N__5861),
            .I(N__5858));
    Span4Mux_v I__1330 (
            .O(N__5858),
            .I(N__5854));
    InMux I__1329 (
            .O(N__5857),
            .I(N__5850));
    Span4Mux_v I__1328 (
            .O(N__5854),
            .I(N__5847));
    InMux I__1327 (
            .O(N__5853),
            .I(N__5844));
    LocalMux I__1326 (
            .O(N__5850),
            .I(N__5841));
    Span4Mux_v I__1325 (
            .O(N__5847),
            .I(N__5838));
    LocalMux I__1324 (
            .O(N__5844),
            .I(N__5833));
    Sp12to4 I__1323 (
            .O(N__5841),
            .I(N__5833));
    Sp12to4 I__1322 (
            .O(N__5838),
            .I(N__5828));
    Span12Mux_v I__1321 (
            .O(N__5833),
            .I(N__5828));
    Odrv12 I__1320 (
            .O(N__5828),
            .I(A_c_1));
    CascadeMux I__1319 (
            .O(N__5825),
            .I(N__5819));
    InMux I__1318 (
            .O(N__5824),
            .I(N__5816));
    InMux I__1317 (
            .O(N__5823),
            .I(N__5813));
    InMux I__1316 (
            .O(N__5822),
            .I(N__5808));
    InMux I__1315 (
            .O(N__5819),
            .I(N__5805));
    LocalMux I__1314 (
            .O(N__5816),
            .I(N__5800));
    LocalMux I__1313 (
            .O(N__5813),
            .I(N__5800));
    InMux I__1312 (
            .O(N__5812),
            .I(N__5795));
    InMux I__1311 (
            .O(N__5811),
            .I(N__5795));
    LocalMux I__1310 (
            .O(N__5808),
            .I(N__5790));
    LocalMux I__1309 (
            .O(N__5805),
            .I(N__5790));
    Span4Mux_v I__1308 (
            .O(N__5800),
            .I(N__5787));
    LocalMux I__1307 (
            .O(N__5795),
            .I(N__5784));
    Span4Mux_v I__1306 (
            .O(N__5790),
            .I(N__5781));
    Span4Mux_h I__1305 (
            .O(N__5787),
            .I(N__5776));
    Span4Mux_v I__1304 (
            .O(N__5784),
            .I(N__5776));
    Odrv4 I__1303 (
            .O(N__5781),
            .I(SIZ_c_1));
    Odrv4 I__1302 (
            .O(N__5776),
            .I(SIZ_c_1));
    CascadeMux I__1301 (
            .O(N__5771),
            .I(N__5767));
    InMux I__1300 (
            .O(N__5770),
            .I(N__5762));
    InMux I__1299 (
            .O(N__5767),
            .I(N__5762));
    LocalMux I__1298 (
            .O(N__5762),
            .I(\U400_BYTE_ENABLE.N_168 ));
    InMux I__1297 (
            .O(N__5759),
            .I(N__5752));
    CascadeMux I__1296 (
            .O(N__5758),
            .I(N__5749));
    InMux I__1295 (
            .O(N__5757),
            .I(N__5745));
    InMux I__1294 (
            .O(N__5756),
            .I(N__5742));
    InMux I__1293 (
            .O(N__5755),
            .I(N__5739));
    LocalMux I__1292 (
            .O(N__5752),
            .I(N__5736));
    InMux I__1291 (
            .O(N__5749),
            .I(N__5731));
    InMux I__1290 (
            .O(N__5748),
            .I(N__5731));
    LocalMux I__1289 (
            .O(N__5745),
            .I(N__5728));
    LocalMux I__1288 (
            .O(N__5742),
            .I(N__5725));
    LocalMux I__1287 (
            .O(N__5739),
            .I(N__5718));
    Span4Mux_v I__1286 (
            .O(N__5736),
            .I(N__5718));
    LocalMux I__1285 (
            .O(N__5731),
            .I(N__5718));
    Span4Mux_v I__1284 (
            .O(N__5728),
            .I(N__5715));
    Span4Mux_v I__1283 (
            .O(N__5725),
            .I(N__5712));
    Span4Mux_h I__1282 (
            .O(N__5718),
            .I(N__5709));
    Span4Mux_h I__1281 (
            .O(N__5715),
            .I(N__5704));
    Span4Mux_h I__1280 (
            .O(N__5712),
            .I(N__5704));
    Span4Mux_v I__1279 (
            .O(N__5709),
            .I(N__5701));
    Odrv4 I__1278 (
            .O(N__5704),
            .I(SIZ_c_0));
    Odrv4 I__1277 (
            .O(N__5701),
            .I(SIZ_c_0));
    IoInMux I__1276 (
            .O(N__5696),
            .I(N__5693));
    LocalMux I__1275 (
            .O(N__5693),
            .I(N__5690));
    Span4Mux_s2_v I__1274 (
            .O(N__5690),
            .I(N__5687));
    Odrv4 I__1273 (
            .O(N__5687),
            .I(un1_LLBEn_i_0_0));
    InMux I__1272 (
            .O(N__5684),
            .I(N__5681));
    LocalMux I__1271 (
            .O(N__5681),
            .I(N__5678));
    Span4Mux_v I__1270 (
            .O(N__5678),
            .I(N__5675));
    Odrv4 I__1269 (
            .O(N__5675),
            .I(TA_EN_i_ess));
    IoInMux I__1268 (
            .O(N__5672),
            .I(N__5669));
    LocalMux I__1267 (
            .O(N__5669),
            .I(N__5666));
    Odrv4 I__1266 (
            .O(N__5666),
            .I(N_526_i));
    InMux I__1265 (
            .O(N__5663),
            .I(N__5660));
    LocalMux I__1264 (
            .O(N__5660),
            .I(N__5657));
    Odrv4 I__1263 (
            .O(N__5657),
            .I(A_c_5));
    CascadeMux I__1262 (
            .O(N__5654),
            .I(N__5651));
    InMux I__1261 (
            .O(N__5651),
            .I(N__5648));
    LocalMux I__1260 (
            .O(N__5648),
            .I(N__5645));
    Span4Mux_v I__1259 (
            .O(N__5645),
            .I(N__5642));
    Odrv4 I__1258 (
            .O(N__5642),
            .I(A_c_13));
    IoInMux I__1257 (
            .O(N__5639),
            .I(N__5636));
    LocalMux I__1256 (
            .O(N__5636),
            .I(N__5633));
    IoSpan4Mux I__1255 (
            .O(N__5633),
            .I(N__5630));
    Span4Mux_s3_h I__1254 (
            .O(N__5630),
            .I(N__5627));
    Span4Mux_h I__1253 (
            .O(N__5627),
            .I(N__5624));
    Odrv4 I__1252 (
            .O(N__5624),
            .I(MA_c_3));
    InMux I__1251 (
            .O(N__5621),
            .I(N__5618));
    LocalMux I__1250 (
            .O(N__5618),
            .I(N__5615));
    Span4Mux_v I__1249 (
            .O(N__5615),
            .I(N__5612));
    Odrv4 I__1248 (
            .O(N__5612),
            .I(A_c_4));
    CascadeMux I__1247 (
            .O(N__5609),
            .I(N__5606));
    InMux I__1246 (
            .O(N__5606),
            .I(N__5603));
    LocalMux I__1245 (
            .O(N__5603),
            .I(N__5600));
    Odrv4 I__1244 (
            .O(N__5600),
            .I(A_c_12));
    IoInMux I__1243 (
            .O(N__5597),
            .I(N__5594));
    LocalMux I__1242 (
            .O(N__5594),
            .I(N__5591));
    Odrv4 I__1241 (
            .O(N__5591),
            .I(MA_c_2));
    InMux I__1240 (
            .O(N__5588),
            .I(N__5585));
    LocalMux I__1239 (
            .O(N__5585),
            .I(N__5582));
    Span4Mux_h I__1238 (
            .O(N__5582),
            .I(N__5579));
    Odrv4 I__1237 (
            .O(N__5579),
            .I(A_c_2));
    CascadeMux I__1236 (
            .O(N__5576),
            .I(N__5573));
    InMux I__1235 (
            .O(N__5573),
            .I(N__5570));
    LocalMux I__1234 (
            .O(N__5570),
            .I(N__5567));
    Odrv4 I__1233 (
            .O(N__5567),
            .I(A_c_10));
    IoInMux I__1232 (
            .O(N__5564),
            .I(N__5561));
    LocalMux I__1231 (
            .O(N__5561),
            .I(N__5558));
    Span4Mux_s1_v I__1230 (
            .O(N__5558),
            .I(N__5555));
    Odrv4 I__1229 (
            .O(N__5555),
            .I(MA_c_0));
    InMux I__1228 (
            .O(N__5552),
            .I(N__5539));
    InMux I__1227 (
            .O(N__5551),
            .I(N__5539));
    InMux I__1226 (
            .O(N__5550),
            .I(N__5534));
    InMux I__1225 (
            .O(N__5549),
            .I(N__5534));
    CascadeMux I__1224 (
            .O(N__5548),
            .I(N__5530));
    CascadeMux I__1223 (
            .O(N__5547),
            .I(N__5524));
    CascadeMux I__1222 (
            .O(N__5546),
            .I(N__5517));
    CascadeMux I__1221 (
            .O(N__5545),
            .I(N__5513));
    CascadeMux I__1220 (
            .O(N__5544),
            .I(N__5510));
    LocalMux I__1219 (
            .O(N__5539),
            .I(N__5505));
    LocalMux I__1218 (
            .O(N__5534),
            .I(N__5505));
    InMux I__1217 (
            .O(N__5533),
            .I(N__5500));
    InMux I__1216 (
            .O(N__5530),
            .I(N__5500));
    InMux I__1215 (
            .O(N__5529),
            .I(N__5497));
    InMux I__1214 (
            .O(N__5528),
            .I(N__5494));
    InMux I__1213 (
            .O(N__5527),
            .I(N__5491));
    InMux I__1212 (
            .O(N__5524),
            .I(N__5484));
    InMux I__1211 (
            .O(N__5523),
            .I(N__5484));
    InMux I__1210 (
            .O(N__5522),
            .I(N__5484));
    InMux I__1209 (
            .O(N__5521),
            .I(N__5477));
    InMux I__1208 (
            .O(N__5520),
            .I(N__5477));
    InMux I__1207 (
            .O(N__5517),
            .I(N__5477));
    InMux I__1206 (
            .O(N__5516),
            .I(N__5474));
    InMux I__1205 (
            .O(N__5513),
            .I(N__5471));
    InMux I__1204 (
            .O(N__5510),
            .I(N__5468));
    Span4Mux_h I__1203 (
            .O(N__5505),
            .I(N__5465));
    LocalMux I__1202 (
            .O(N__5500),
            .I(N__5458));
    LocalMux I__1201 (
            .O(N__5497),
            .I(N__5458));
    LocalMux I__1200 (
            .O(N__5494),
            .I(N__5458));
    LocalMux I__1199 (
            .O(N__5491),
            .I(N__5449));
    LocalMux I__1198 (
            .O(N__5484),
            .I(N__5449));
    LocalMux I__1197 (
            .O(N__5477),
            .I(N__5449));
    LocalMux I__1196 (
            .O(N__5474),
            .I(N__5446));
    LocalMux I__1195 (
            .O(N__5471),
            .I(N__5441));
    LocalMux I__1194 (
            .O(N__5468),
            .I(N__5441));
    Span4Mux_v I__1193 (
            .O(N__5465),
            .I(N__5436));
    Span4Mux_v I__1192 (
            .O(N__5458),
            .I(N__5436));
    InMux I__1191 (
            .O(N__5457),
            .I(N__5431));
    InMux I__1190 (
            .O(N__5456),
            .I(N__5431));
    Span4Mux_v I__1189 (
            .O(N__5449),
            .I(N__5428));
    Span4Mux_v I__1188 (
            .O(N__5446),
            .I(N__5423));
    Span4Mux_h I__1187 (
            .O(N__5441),
            .I(N__5423));
    Odrv4 I__1186 (
            .O(N__5436),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1185 (
            .O(N__5431),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1184 (
            .O(N__5428),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1183 (
            .O(N__5423),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    InMux I__1182 (
            .O(N__5414),
            .I(N__5411));
    LocalMux I__1181 (
            .O(N__5411),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_0_0 ));
    CascadeMux I__1180 (
            .O(N__5408),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_1_0_cascade_ ));
    InMux I__1179 (
            .O(N__5405),
            .I(N__5402));
    LocalMux I__1178 (
            .O(N__5402),
            .I(N__5399));
    Span4Mux_v I__1177 (
            .O(N__5399),
            .I(N__5388));
    InMux I__1176 (
            .O(N__5398),
            .I(N__5383));
    InMux I__1175 (
            .O(N__5397),
            .I(N__5383));
    InMux I__1174 (
            .O(N__5396),
            .I(N__5380));
    InMux I__1173 (
            .O(N__5395),
            .I(N__5377));
    InMux I__1172 (
            .O(N__5394),
            .I(N__5370));
    InMux I__1171 (
            .O(N__5393),
            .I(N__5370));
    InMux I__1170 (
            .O(N__5392),
            .I(N__5370));
    InMux I__1169 (
            .O(N__5391),
            .I(N__5367));
    Odrv4 I__1168 (
            .O(N__5388),
            .I(\U400_SDRAM.N_114 ));
    LocalMux I__1167 (
            .O(N__5383),
            .I(\U400_SDRAM.N_114 ));
    LocalMux I__1166 (
            .O(N__5380),
            .I(\U400_SDRAM.N_114 ));
    LocalMux I__1165 (
            .O(N__5377),
            .I(\U400_SDRAM.N_114 ));
    LocalMux I__1164 (
            .O(N__5370),
            .I(\U400_SDRAM.N_114 ));
    LocalMux I__1163 (
            .O(N__5367),
            .I(\U400_SDRAM.N_114 ));
    CEMux I__1162 (
            .O(N__5354),
            .I(N__5351));
    LocalMux I__1161 (
            .O(N__5351),
            .I(N__5346));
    InMux I__1160 (
            .O(N__5350),
            .I(N__5341));
    InMux I__1159 (
            .O(N__5349),
            .I(N__5341));
    Odrv12 I__1158 (
            .O(N__5346),
            .I(\U400_SDRAM.N_71 ));
    LocalMux I__1157 (
            .O(N__5341),
            .I(\U400_SDRAM.N_71 ));
    CascadeMux I__1156 (
            .O(N__5336),
            .I(N__5333));
    InMux I__1155 (
            .O(N__5333),
            .I(N__5330));
    LocalMux I__1154 (
            .O(N__5330),
            .I(N__5327));
    Span12Mux_s7_v I__1153 (
            .O(N__5327),
            .I(N__5324));
    Odrv12 I__1152 (
            .O(N__5324),
            .I(A_c_25));
    IoInMux I__1151 (
            .O(N__5321),
            .I(N__5318));
    LocalMux I__1150 (
            .O(N__5318),
            .I(N__5315));
    Odrv12 I__1149 (
            .O(N__5315),
            .I(MA_c_11));
    CascadeMux I__1148 (
            .O(N__5312),
            .I(N__5309));
    InMux I__1147 (
            .O(N__5309),
            .I(N__5306));
    LocalMux I__1146 (
            .O(N__5306),
            .I(N__5303));
    Odrv12 I__1145 (
            .O(N__5303),
            .I(A_c_7));
    InMux I__1144 (
            .O(N__5300),
            .I(N__5297));
    LocalMux I__1143 (
            .O(N__5297),
            .I(N__5294));
    IoSpan4Mux I__1142 (
            .O(N__5294),
            .I(N__5291));
    Odrv4 I__1141 (
            .O(N__5291),
            .I(A_c_15));
    InMux I__1140 (
            .O(N__5288),
            .I(N__5285));
    LocalMux I__1139 (
            .O(N__5285),
            .I(\U400_SDRAM.MA_5_iv_0_5 ));
    IoInMux I__1138 (
            .O(N__5282),
            .I(N__5279));
    LocalMux I__1137 (
            .O(N__5279),
            .I(N__5276));
    Span4Mux_s2_v I__1136 (
            .O(N__5276),
            .I(N__5273));
    Span4Mux_h I__1135 (
            .O(N__5273),
            .I(N__5270));
    Odrv4 I__1134 (
            .O(N__5270),
            .I(MA_c_5));
    InMux I__1133 (
            .O(N__5267),
            .I(N__5264));
    LocalMux I__1132 (
            .O(N__5264),
            .I(\U400_BYTE_ENABLE.N_101_i ));
    CascadeMux I__1131 (
            .O(N__5261),
            .I(\U400_BYTE_ENABLE.N_101_i_cascade_ ));
    IoInMux I__1130 (
            .O(N__5258),
            .I(N__5255));
    LocalMux I__1129 (
            .O(N__5255),
            .I(N__5252));
    Span4Mux_s3_v I__1128 (
            .O(N__5252),
            .I(N__5249));
    Odrv4 I__1127 (
            .O(N__5249),
            .I(un1_LMBEn_i_0_0));
    InMux I__1126 (
            .O(N__5246),
            .I(N__5242));
    InMux I__1125 (
            .O(N__5245),
            .I(N__5239));
    LocalMux I__1124 (
            .O(N__5242),
            .I(N__5235));
    LocalMux I__1123 (
            .O(N__5239),
            .I(N__5232));
    InMux I__1122 (
            .O(N__5238),
            .I(N__5229));
    Span4Mux_v I__1121 (
            .O(N__5235),
            .I(N__5226));
    Span4Mux_v I__1120 (
            .O(N__5232),
            .I(N__5223));
    LocalMux I__1119 (
            .O(N__5229),
            .I(N__5220));
    Span4Mux_v I__1118 (
            .O(N__5226),
            .I(N__5217));
    Sp12to4 I__1117 (
            .O(N__5223),
            .I(N__5214));
    Span4Mux_h I__1116 (
            .O(N__5220),
            .I(N__5211));
    Span4Mux_v I__1115 (
            .O(N__5217),
            .I(N__5208));
    Span12Mux_s6_h I__1114 (
            .O(N__5214),
            .I(N__5203));
    Sp12to4 I__1113 (
            .O(N__5211),
            .I(N__5203));
    Sp12to4 I__1112 (
            .O(N__5208),
            .I(N__5198));
    Span12Mux_v I__1111 (
            .O(N__5203),
            .I(N__5198));
    Odrv12 I__1110 (
            .O(N__5198),
            .I(A_c_0));
    CascadeMux I__1109 (
            .O(N__5195),
            .I(N__5190));
    IoInMux I__1108 (
            .O(N__5194),
            .I(N__5187));
    InMux I__1107 (
            .O(N__5193),
            .I(N__5184));
    InMux I__1106 (
            .O(N__5190),
            .I(N__5180));
    LocalMux I__1105 (
            .O(N__5187),
            .I(N__5177));
    LocalMux I__1104 (
            .O(N__5184),
            .I(N__5174));
    InMux I__1103 (
            .O(N__5183),
            .I(N__5171));
    LocalMux I__1102 (
            .O(N__5180),
            .I(N__5168));
    Odrv12 I__1101 (
            .O(N__5177),
            .I(RAM_SPACE_i_o3_0_o2dup));
    Odrv4 I__1100 (
            .O(N__5174),
            .I(RAM_SPACE_i_o3_0_o2dup));
    LocalMux I__1099 (
            .O(N__5171),
            .I(RAM_SPACE_i_o3_0_o2dup));
    Odrv4 I__1098 (
            .O(N__5168),
            .I(RAM_SPACE_i_o3_0_o2dup));
    InMux I__1097 (
            .O(N__5159),
            .I(N__5156));
    LocalMux I__1096 (
            .O(N__5156),
            .I(\U400_SDRAM.un1_SDRAM_COUNTER52_2_0_i_1 ));
    CascadeMux I__1095 (
            .O(N__5153),
            .I(\U400_SDRAM.N_195_cascade_ ));
    InMux I__1094 (
            .O(N__5150),
            .I(N__5147));
    LocalMux I__1093 (
            .O(N__5147),
            .I(\U400_SDRAM.N_94 ));
    CascadeMux I__1092 (
            .O(N__5144),
            .I(N__5140));
    InMux I__1091 (
            .O(N__5143),
            .I(N__5137));
    InMux I__1090 (
            .O(N__5140),
            .I(N__5134));
    LocalMux I__1089 (
            .O(N__5137),
            .I(N__5131));
    LocalMux I__1088 (
            .O(N__5134),
            .I(N__5128));
    Span4Mux_v I__1087 (
            .O(N__5131),
            .I(N__5123));
    Span4Mux_v I__1086 (
            .O(N__5128),
            .I(N__5123));
    Odrv4 I__1085 (
            .O(N__5123),
            .I(U400_ADDRESS_DECODE_RAM_SPACE_i_o3_0_o2_1));
    InMux I__1084 (
            .O(N__5120),
            .I(N__5117));
    LocalMux I__1083 (
            .O(N__5117),
            .I(N__5113));
    InMux I__1082 (
            .O(N__5116),
            .I(N__5110));
    Span4Mux_h I__1081 (
            .O(N__5113),
            .I(N__5107));
    LocalMux I__1080 (
            .O(N__5110),
            .I(N__5104));
    Span4Mux_h I__1079 (
            .O(N__5107),
            .I(N__5101));
    Span12Mux_s10_h I__1078 (
            .O(N__5104),
            .I(N__5098));
    Span4Mux_v I__1077 (
            .O(N__5101),
            .I(N__5095));
    Odrv12 I__1076 (
            .O(N__5098),
            .I(A_c_31));
    Odrv4 I__1075 (
            .O(N__5095),
            .I(A_c_31));
    CascadeMux I__1074 (
            .O(N__5090),
            .I(N__5087));
    InMux I__1073 (
            .O(N__5087),
            .I(N__5084));
    LocalMux I__1072 (
            .O(N__5084),
            .I(N__5080));
    InMux I__1071 (
            .O(N__5083),
            .I(N__5077));
    Span4Mux_v I__1070 (
            .O(N__5080),
            .I(N__5072));
    LocalMux I__1069 (
            .O(N__5077),
            .I(N__5072));
    Span4Mux_v I__1068 (
            .O(N__5072),
            .I(N__5069));
    Sp12to4 I__1067 (
            .O(N__5069),
            .I(N__5066));
    Odrv12 I__1066 (
            .O(N__5066),
            .I(U400_ADDRESS_DECODE_RAM_SPACE_i_o3_0_o2_2));
    InMux I__1065 (
            .O(N__5063),
            .I(N__5060));
    LocalMux I__1064 (
            .O(N__5060),
            .I(N__5057));
    Odrv12 I__1063 (
            .O(N__5057),
            .I(TSn_c));
    InMux I__1062 (
            .O(N__5054),
            .I(N__5051));
    LocalMux I__1061 (
            .O(N__5051),
            .I(\U400_SDRAM.N_225 ));
    CascadeMux I__1060 (
            .O(N__5048),
            .I(N__5040));
    InMux I__1059 (
            .O(N__5047),
            .I(N__5036));
    InMux I__1058 (
            .O(N__5046),
            .I(N__5031));
    InMux I__1057 (
            .O(N__5045),
            .I(N__5031));
    InMux I__1056 (
            .O(N__5044),
            .I(N__5028));
    InMux I__1055 (
            .O(N__5043),
            .I(N__5025));
    InMux I__1054 (
            .O(N__5040),
            .I(N__5022));
    InMux I__1053 (
            .O(N__5039),
            .I(N__5019));
    LocalMux I__1052 (
            .O(N__5036),
            .I(N__5016));
    LocalMux I__1051 (
            .O(N__5031),
            .I(\U400_SDRAM.N_236 ));
    LocalMux I__1050 (
            .O(N__5028),
            .I(\U400_SDRAM.N_236 ));
    LocalMux I__1049 (
            .O(N__5025),
            .I(\U400_SDRAM.N_236 ));
    LocalMux I__1048 (
            .O(N__5022),
            .I(\U400_SDRAM.N_236 ));
    LocalMux I__1047 (
            .O(N__5019),
            .I(\U400_SDRAM.N_236 ));
    Odrv4 I__1046 (
            .O(N__5016),
            .I(\U400_SDRAM.N_236 ));
    InMux I__1045 (
            .O(N__5003),
            .I(N__4990));
    InMux I__1044 (
            .O(N__5002),
            .I(N__4990));
    InMux I__1043 (
            .O(N__5001),
            .I(N__4987));
    InMux I__1042 (
            .O(N__5000),
            .I(N__4984));
    InMux I__1041 (
            .O(N__4999),
            .I(N__4975));
    InMux I__1040 (
            .O(N__4998),
            .I(N__4975));
    InMux I__1039 (
            .O(N__4997),
            .I(N__4975));
    InMux I__1038 (
            .O(N__4996),
            .I(N__4975));
    InMux I__1037 (
            .O(N__4995),
            .I(N__4972));
    LocalMux I__1036 (
            .O(N__4990),
            .I(\U400_SDRAM.RAM_CYCLE_STARTZ0 ));
    LocalMux I__1035 (
            .O(N__4987),
            .I(\U400_SDRAM.RAM_CYCLE_STARTZ0 ));
    LocalMux I__1034 (
            .O(N__4984),
            .I(\U400_SDRAM.RAM_CYCLE_STARTZ0 ));
    LocalMux I__1033 (
            .O(N__4975),
            .I(\U400_SDRAM.RAM_CYCLE_STARTZ0 ));
    LocalMux I__1032 (
            .O(N__4972),
            .I(\U400_SDRAM.RAM_CYCLE_STARTZ0 ));
    InMux I__1031 (
            .O(N__4961),
            .I(N__4958));
    LocalMux I__1030 (
            .O(N__4958),
            .I(\U400_SDRAM.N_228 ));
    CascadeMux I__1029 (
            .O(N__4955),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_a2_2_0_1_cascade_ ));
    CascadeMux I__1028 (
            .O(N__4952),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_1_1_cascade_ ));
    CascadeMux I__1027 (
            .O(N__4949),
            .I(N__4943));
    InMux I__1026 (
            .O(N__4948),
            .I(N__4937));
    InMux I__1025 (
            .O(N__4947),
            .I(N__4932));
    InMux I__1024 (
            .O(N__4946),
            .I(N__4932));
    InMux I__1023 (
            .O(N__4943),
            .I(N__4927));
    InMux I__1022 (
            .O(N__4942),
            .I(N__4920));
    InMux I__1021 (
            .O(N__4941),
            .I(N__4920));
    InMux I__1020 (
            .O(N__4940),
            .I(N__4917));
    LocalMux I__1019 (
            .O(N__4937),
            .I(N__4914));
    LocalMux I__1018 (
            .O(N__4932),
            .I(N__4911));
    InMux I__1017 (
            .O(N__4931),
            .I(N__4902));
    InMux I__1016 (
            .O(N__4930),
            .I(N__4902));
    LocalMux I__1015 (
            .O(N__4927),
            .I(N__4895));
    InMux I__1014 (
            .O(N__4926),
            .I(N__4892));
    InMux I__1013 (
            .O(N__4925),
            .I(N__4889));
    LocalMux I__1012 (
            .O(N__4920),
            .I(N__4884));
    LocalMux I__1011 (
            .O(N__4917),
            .I(N__4884));
    Span4Mux_h I__1010 (
            .O(N__4914),
            .I(N__4881));
    Span4Mux_v I__1009 (
            .O(N__4911),
            .I(N__4878));
    InMux I__1008 (
            .O(N__4910),
            .I(N__4871));
    InMux I__1007 (
            .O(N__4909),
            .I(N__4871));
    InMux I__1006 (
            .O(N__4908),
            .I(N__4871));
    InMux I__1005 (
            .O(N__4907),
            .I(N__4868));
    LocalMux I__1004 (
            .O(N__4902),
            .I(N__4865));
    InMux I__1003 (
            .O(N__4901),
            .I(N__4862));
    InMux I__1002 (
            .O(N__4900),
            .I(N__4857));
    InMux I__1001 (
            .O(N__4899),
            .I(N__4857));
    InMux I__1000 (
            .O(N__4898),
            .I(N__4854));
    Span4Mux_v I__999 (
            .O(N__4895),
            .I(N__4845));
    LocalMux I__998 (
            .O(N__4892),
            .I(N__4845));
    LocalMux I__997 (
            .O(N__4889),
            .I(N__4845));
    Span4Mux_h I__996 (
            .O(N__4884),
            .I(N__4845));
    Odrv4 I__995 (
            .O(N__4881),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__994 (
            .O(N__4878),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__993 (
            .O(N__4871),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__992 (
            .O(N__4868),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv12 I__991 (
            .O(N__4865),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__990 (
            .O(N__4862),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__989 (
            .O(N__4857),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__988 (
            .O(N__4854),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__987 (
            .O(N__4845),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    InMux I__986 (
            .O(N__4826),
            .I(N__4823));
    LocalMux I__985 (
            .O(N__4823),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_2_1 ));
    InMux I__984 (
            .O(N__4820),
            .I(N__4814));
    InMux I__983 (
            .O(N__4819),
            .I(N__4810));
    InMux I__982 (
            .O(N__4818),
            .I(N__4803));
    InMux I__981 (
            .O(N__4817),
            .I(N__4800));
    LocalMux I__980 (
            .O(N__4814),
            .I(N__4791));
    CascadeMux I__979 (
            .O(N__4813),
            .I(N__4786));
    LocalMux I__978 (
            .O(N__4810),
            .I(N__4782));
    InMux I__977 (
            .O(N__4809),
            .I(N__4775));
    InMux I__976 (
            .O(N__4808),
            .I(N__4775));
    InMux I__975 (
            .O(N__4807),
            .I(N__4775));
    InMux I__974 (
            .O(N__4806),
            .I(N__4770));
    LocalMux I__973 (
            .O(N__4803),
            .I(N__4765));
    LocalMux I__972 (
            .O(N__4800),
            .I(N__4765));
    InMux I__971 (
            .O(N__4799),
            .I(N__4760));
    InMux I__970 (
            .O(N__4798),
            .I(N__4760));
    InMux I__969 (
            .O(N__4797),
            .I(N__4757));
    InMux I__968 (
            .O(N__4796),
            .I(N__4754));
    InMux I__967 (
            .O(N__4795),
            .I(N__4751));
    InMux I__966 (
            .O(N__4794),
            .I(N__4748));
    Span4Mux_h I__965 (
            .O(N__4791),
            .I(N__4745));
    InMux I__964 (
            .O(N__4790),
            .I(N__4742));
    InMux I__963 (
            .O(N__4789),
            .I(N__4739));
    InMux I__962 (
            .O(N__4786),
            .I(N__4734));
    InMux I__961 (
            .O(N__4785),
            .I(N__4734));
    Span4Mux_v I__960 (
            .O(N__4782),
            .I(N__4731));
    LocalMux I__959 (
            .O(N__4775),
            .I(N__4728));
    InMux I__958 (
            .O(N__4774),
            .I(N__4725));
    InMux I__957 (
            .O(N__4773),
            .I(N__4722));
    LocalMux I__956 (
            .O(N__4770),
            .I(N__4717));
    Span4Mux_h I__955 (
            .O(N__4765),
            .I(N__4717));
    LocalMux I__954 (
            .O(N__4760),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__953 (
            .O(N__4757),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__952 (
            .O(N__4754),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__951 (
            .O(N__4751),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__950 (
            .O(N__4748),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__949 (
            .O(N__4745),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__948 (
            .O(N__4742),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__947 (
            .O(N__4739),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__946 (
            .O(N__4734),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__945 (
            .O(N__4731),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv12 I__944 (
            .O(N__4728),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__943 (
            .O(N__4725),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__942 (
            .O(N__4722),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__941 (
            .O(N__4717),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    CascadeMux I__940 (
            .O(N__4688),
            .I(N__4684));
    CascadeMux I__939 (
            .O(N__4687),
            .I(N__4681));
    InMux I__938 (
            .O(N__4684),
            .I(N__4675));
    InMux I__937 (
            .O(N__4681),
            .I(N__4672));
    InMux I__936 (
            .O(N__4680),
            .I(N__4668));
    CascadeMux I__935 (
            .O(N__4679),
            .I(N__4665));
    CascadeMux I__934 (
            .O(N__4678),
            .I(N__4660));
    LocalMux I__933 (
            .O(N__4675),
            .I(N__4656));
    LocalMux I__932 (
            .O(N__4672),
            .I(N__4653));
    InMux I__931 (
            .O(N__4671),
            .I(N__4650));
    LocalMux I__930 (
            .O(N__4668),
            .I(N__4647));
    InMux I__929 (
            .O(N__4665),
            .I(N__4640));
    InMux I__928 (
            .O(N__4664),
            .I(N__4640));
    InMux I__927 (
            .O(N__4663),
            .I(N__4640));
    InMux I__926 (
            .O(N__4660),
            .I(N__4635));
    InMux I__925 (
            .O(N__4659),
            .I(N__4635));
    Span4Mux_v I__924 (
            .O(N__4656),
            .I(N__4630));
    Span4Mux_v I__923 (
            .O(N__4653),
            .I(N__4630));
    LocalMux I__922 (
            .O(N__4650),
            .I(\U400_SDRAM.WRITE_CYCLEZ0 ));
    Odrv4 I__921 (
            .O(N__4647),
            .I(\U400_SDRAM.WRITE_CYCLEZ0 ));
    LocalMux I__920 (
            .O(N__4640),
            .I(\U400_SDRAM.WRITE_CYCLEZ0 ));
    LocalMux I__919 (
            .O(N__4635),
            .I(\U400_SDRAM.WRITE_CYCLEZ0 ));
    Odrv4 I__918 (
            .O(N__4630),
            .I(\U400_SDRAM.WRITE_CYCLEZ0 ));
    CascadeMux I__917 (
            .O(N__4619),
            .I(N__4612));
    InMux I__916 (
            .O(N__4618),
            .I(N__4605));
    InMux I__915 (
            .O(N__4617),
            .I(N__4602));
    CascadeMux I__914 (
            .O(N__4616),
            .I(N__4599));
    CascadeMux I__913 (
            .O(N__4615),
            .I(N__4593));
    InMux I__912 (
            .O(N__4612),
            .I(N__4580));
    InMux I__911 (
            .O(N__4611),
            .I(N__4580));
    InMux I__910 (
            .O(N__4610),
            .I(N__4580));
    InMux I__909 (
            .O(N__4609),
            .I(N__4575));
    InMux I__908 (
            .O(N__4608),
            .I(N__4575));
    LocalMux I__907 (
            .O(N__4605),
            .I(N__4569));
    LocalMux I__906 (
            .O(N__4602),
            .I(N__4566));
    InMux I__905 (
            .O(N__4599),
            .I(N__4561));
    InMux I__904 (
            .O(N__4598),
            .I(N__4561));
    CascadeMux I__903 (
            .O(N__4597),
            .I(N__4558));
    InMux I__902 (
            .O(N__4596),
            .I(N__4555));
    InMux I__901 (
            .O(N__4593),
            .I(N__4550));
    InMux I__900 (
            .O(N__4592),
            .I(N__4550));
    InMux I__899 (
            .O(N__4591),
            .I(N__4547));
    InMux I__898 (
            .O(N__4590),
            .I(N__4540));
    InMux I__897 (
            .O(N__4589),
            .I(N__4540));
    InMux I__896 (
            .O(N__4588),
            .I(N__4540));
    InMux I__895 (
            .O(N__4587),
            .I(N__4537));
    LocalMux I__894 (
            .O(N__4580),
            .I(N__4532));
    LocalMux I__893 (
            .O(N__4575),
            .I(N__4532));
    InMux I__892 (
            .O(N__4574),
            .I(N__4529));
    InMux I__891 (
            .O(N__4573),
            .I(N__4524));
    InMux I__890 (
            .O(N__4572),
            .I(N__4524));
    Span4Mux_v I__889 (
            .O(N__4569),
            .I(N__4517));
    Span4Mux_v I__888 (
            .O(N__4566),
            .I(N__4517));
    LocalMux I__887 (
            .O(N__4561),
            .I(N__4517));
    InMux I__886 (
            .O(N__4558),
            .I(N__4514));
    LocalMux I__885 (
            .O(N__4555),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__884 (
            .O(N__4550),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__883 (
            .O(N__4547),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__882 (
            .O(N__4540),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__881 (
            .O(N__4537),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__880 (
            .O(N__4532),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__879 (
            .O(N__4529),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__878 (
            .O(N__4524),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__877 (
            .O(N__4517),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__876 (
            .O(N__4514),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    InMux I__875 (
            .O(N__4493),
            .I(N__4485));
    InMux I__874 (
            .O(N__4492),
            .I(N__4482));
    InMux I__873 (
            .O(N__4491),
            .I(N__4479));
    InMux I__872 (
            .O(N__4490),
            .I(N__4474));
    InMux I__871 (
            .O(N__4489),
            .I(N__4474));
    InMux I__870 (
            .O(N__4488),
            .I(N__4470));
    LocalMux I__869 (
            .O(N__4485),
            .I(N__4463));
    LocalMux I__868 (
            .O(N__4482),
            .I(N__4463));
    LocalMux I__867 (
            .O(N__4479),
            .I(N__4456));
    LocalMux I__866 (
            .O(N__4474),
            .I(N__4456));
    InMux I__865 (
            .O(N__4473),
            .I(N__4453));
    LocalMux I__864 (
            .O(N__4470),
            .I(N__4450));
    InMux I__863 (
            .O(N__4469),
            .I(N__4445));
    InMux I__862 (
            .O(N__4468),
            .I(N__4445));
    Span4Mux_v I__861 (
            .O(N__4463),
            .I(N__4438));
    InMux I__860 (
            .O(N__4462),
            .I(N__4435));
    InMux I__859 (
            .O(N__4461),
            .I(N__4432));
    Span4Mux_h I__858 (
            .O(N__4456),
            .I(N__4429));
    LocalMux I__857 (
            .O(N__4453),
            .I(N__4426));
    Span4Mux_v I__856 (
            .O(N__4450),
            .I(N__4421));
    LocalMux I__855 (
            .O(N__4445),
            .I(N__4421));
    InMux I__854 (
            .O(N__4444),
            .I(N__4414));
    InMux I__853 (
            .O(N__4443),
            .I(N__4414));
    InMux I__852 (
            .O(N__4442),
            .I(N__4414));
    InMux I__851 (
            .O(N__4441),
            .I(N__4411));
    Odrv4 I__850 (
            .O(N__4438),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__849 (
            .O(N__4435),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__848 (
            .O(N__4432),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__847 (
            .O(N__4429),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__846 (
            .O(N__4426),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__845 (
            .O(N__4421),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__844 (
            .O(N__4414),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__843 (
            .O(N__4411),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__842 (
            .O(N__4394),
            .I(N__4390));
    InMux I__841 (
            .O(N__4393),
            .I(N__4387));
    LocalMux I__840 (
            .O(N__4390),
            .I(N__4382));
    LocalMux I__839 (
            .O(N__4387),
            .I(N__4382));
    Span4Mux_h I__838 (
            .O(N__4382),
            .I(N__4377));
    InMux I__837 (
            .O(N__4381),
            .I(N__4374));
    InMux I__836 (
            .O(N__4380),
            .I(N__4371));
    Odrv4 I__835 (
            .O(N__4377),
            .I(\U400_SDRAM.N_256 ));
    LocalMux I__834 (
            .O(N__4374),
            .I(\U400_SDRAM.N_256 ));
    LocalMux I__833 (
            .O(N__4371),
            .I(\U400_SDRAM.N_256 ));
    CascadeMux I__832 (
            .O(N__4364),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_a2_0_1_0_cascade_ ));
    InMux I__831 (
            .O(N__4361),
            .I(N__4358));
    LocalMux I__830 (
            .O(N__4358),
            .I(N__4353));
    InMux I__829 (
            .O(N__4357),
            .I(N__4350));
    InMux I__828 (
            .O(N__4356),
            .I(N__4346));
    Span4Mux_v I__827 (
            .O(N__4353),
            .I(N__4341));
    LocalMux I__826 (
            .O(N__4350),
            .I(N__4341));
    InMux I__825 (
            .O(N__4349),
            .I(N__4338));
    LocalMux I__824 (
            .O(N__4346),
            .I(N__4328));
    Span4Mux_h I__823 (
            .O(N__4341),
            .I(N__4325));
    LocalMux I__822 (
            .O(N__4338),
            .I(N__4322));
    InMux I__821 (
            .O(N__4337),
            .I(N__4317));
    InMux I__820 (
            .O(N__4336),
            .I(N__4317));
    InMux I__819 (
            .O(N__4335),
            .I(N__4308));
    InMux I__818 (
            .O(N__4334),
            .I(N__4308));
    InMux I__817 (
            .O(N__4333),
            .I(N__4308));
    InMux I__816 (
            .O(N__4332),
            .I(N__4308));
    InMux I__815 (
            .O(N__4331),
            .I(N__4305));
    Odrv4 I__814 (
            .O(N__4328),
            .I(\U400_SDRAM.N_97 ));
    Odrv4 I__813 (
            .O(N__4325),
            .I(\U400_SDRAM.N_97 ));
    Odrv4 I__812 (
            .O(N__4322),
            .I(\U400_SDRAM.N_97 ));
    LocalMux I__811 (
            .O(N__4317),
            .I(\U400_SDRAM.N_97 ));
    LocalMux I__810 (
            .O(N__4308),
            .I(\U400_SDRAM.N_97 ));
    LocalMux I__809 (
            .O(N__4305),
            .I(\U400_SDRAM.N_97 ));
    CascadeMux I__808 (
            .O(N__4292),
            .I(\U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0_cascade_ ));
    CascadeMux I__807 (
            .O(N__4289),
            .I(N__4285));
    InMux I__806 (
            .O(N__4288),
            .I(N__4281));
    InMux I__805 (
            .O(N__4285),
            .I(N__4273));
    InMux I__804 (
            .O(N__4284),
            .I(N__4273));
    LocalMux I__803 (
            .O(N__4281),
            .I(N__4270));
    InMux I__802 (
            .O(N__4280),
            .I(N__4263));
    InMux I__801 (
            .O(N__4279),
            .I(N__4263));
    InMux I__800 (
            .O(N__4278),
            .I(N__4263));
    LocalMux I__799 (
            .O(N__4273),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_2 ));
    Odrv4 I__798 (
            .O(N__4270),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_2 ));
    LocalMux I__797 (
            .O(N__4263),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_2 ));
    CascadeMux I__796 (
            .O(N__4256),
            .I(N__4250));
    CascadeMux I__795 (
            .O(N__4255),
            .I(N__4246));
    CascadeMux I__794 (
            .O(N__4254),
            .I(N__4243));
    InMux I__793 (
            .O(N__4253),
            .I(N__4240));
    InMux I__792 (
            .O(N__4250),
            .I(N__4237));
    InMux I__791 (
            .O(N__4249),
            .I(N__4230));
    InMux I__790 (
            .O(N__4246),
            .I(N__4230));
    InMux I__789 (
            .O(N__4243),
            .I(N__4230));
    LocalMux I__788 (
            .O(N__4240),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_3 ));
    LocalMux I__787 (
            .O(N__4237),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_3 ));
    LocalMux I__786 (
            .O(N__4230),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_3 ));
    CascadeMux I__785 (
            .O(N__4223),
            .I(N__4219));
    CascadeMux I__784 (
            .O(N__4222),
            .I(N__4214));
    InMux I__783 (
            .O(N__4219),
            .I(N__4207));
    InMux I__782 (
            .O(N__4218),
            .I(N__4207));
    InMux I__781 (
            .O(N__4217),
            .I(N__4204));
    InMux I__780 (
            .O(N__4214),
            .I(N__4197));
    InMux I__779 (
            .O(N__4213),
            .I(N__4197));
    InMux I__778 (
            .O(N__4212),
            .I(N__4197));
    LocalMux I__777 (
            .O(N__4207),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_1 ));
    LocalMux I__776 (
            .O(N__4204),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_1 ));
    LocalMux I__775 (
            .O(N__4197),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_1 ));
    InMux I__774 (
            .O(N__4190),
            .I(N__4186));
    InMux I__773 (
            .O(N__4189),
            .I(N__4183));
    LocalMux I__772 (
            .O(N__4186),
            .I(\U400_SDRAM.CO1 ));
    LocalMux I__771 (
            .O(N__4183),
            .I(\U400_SDRAM.CO1 ));
    CascadeMux I__770 (
            .O(N__4178),
            .I(N__4174));
    InMux I__769 (
            .O(N__4177),
            .I(N__4168));
    InMux I__768 (
            .O(N__4174),
            .I(N__4163));
    InMux I__767 (
            .O(N__4173),
            .I(N__4163));
    InMux I__766 (
            .O(N__4172),
            .I(N__4158));
    InMux I__765 (
            .O(N__4171),
            .I(N__4158));
    LocalMux I__764 (
            .O(N__4168),
            .I(\U400_SDRAM.TA_COUNTER23 ));
    LocalMux I__763 (
            .O(N__4163),
            .I(\U400_SDRAM.TA_COUNTER23 ));
    LocalMux I__762 (
            .O(N__4158),
            .I(\U400_SDRAM.TA_COUNTER23 ));
    InMux I__761 (
            .O(N__4151),
            .I(N__4143));
    InMux I__760 (
            .O(N__4150),
            .I(N__4138));
    InMux I__759 (
            .O(N__4149),
            .I(N__4138));
    InMux I__758 (
            .O(N__4148),
            .I(N__4135));
    InMux I__757 (
            .O(N__4147),
            .I(N__4130));
    InMux I__756 (
            .O(N__4146),
            .I(N__4130));
    LocalMux I__755 (
            .O(N__4143),
            .I(\U400_SDRAM.TACKZ0 ));
    LocalMux I__754 (
            .O(N__4138),
            .I(\U400_SDRAM.TACKZ0 ));
    LocalMux I__753 (
            .O(N__4135),
            .I(\U400_SDRAM.TACKZ0 ));
    LocalMux I__752 (
            .O(N__4130),
            .I(\U400_SDRAM.TACKZ0 ));
    CascadeMux I__751 (
            .O(N__4121),
            .I(\U400_SDRAM.TA_COUNTER_7_f1_0_0_cascade_ ));
    InMux I__750 (
            .O(N__4118),
            .I(N__4112));
    InMux I__749 (
            .O(N__4117),
            .I(N__4112));
    LocalMux I__748 (
            .O(N__4112),
            .I(\U400_SDRAM.TA_COUNTER_0_sqmuxa ));
    InMux I__747 (
            .O(N__4109),
            .I(N__4095));
    InMux I__746 (
            .O(N__4108),
            .I(N__4095));
    InMux I__745 (
            .O(N__4107),
            .I(N__4095));
    InMux I__744 (
            .O(N__4106),
            .I(N__4092));
    InMux I__743 (
            .O(N__4105),
            .I(N__4083));
    InMux I__742 (
            .O(N__4104),
            .I(N__4083));
    InMux I__741 (
            .O(N__4103),
            .I(N__4083));
    InMux I__740 (
            .O(N__4102),
            .I(N__4083));
    LocalMux I__739 (
            .O(N__4095),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_0 ));
    LocalMux I__738 (
            .O(N__4092),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_0 ));
    LocalMux I__737 (
            .O(N__4083),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_0 ));
    ClkMux I__736 (
            .O(N__4076),
            .I(N__3995));
    ClkMux I__735 (
            .O(N__4075),
            .I(N__3995));
    ClkMux I__734 (
            .O(N__4074),
            .I(N__3995));
    ClkMux I__733 (
            .O(N__4073),
            .I(N__3995));
    ClkMux I__732 (
            .O(N__4072),
            .I(N__3995));
    ClkMux I__731 (
            .O(N__4071),
            .I(N__3995));
    ClkMux I__730 (
            .O(N__4070),
            .I(N__3995));
    ClkMux I__729 (
            .O(N__4069),
            .I(N__3995));
    ClkMux I__728 (
            .O(N__4068),
            .I(N__3995));
    ClkMux I__727 (
            .O(N__4067),
            .I(N__3995));
    ClkMux I__726 (
            .O(N__4066),
            .I(N__3995));
    ClkMux I__725 (
            .O(N__4065),
            .I(N__3995));
    ClkMux I__724 (
            .O(N__4064),
            .I(N__3995));
    ClkMux I__723 (
            .O(N__4063),
            .I(N__3995));
    ClkMux I__722 (
            .O(N__4062),
            .I(N__3995));
    ClkMux I__721 (
            .O(N__4061),
            .I(N__3995));
    ClkMux I__720 (
            .O(N__4060),
            .I(N__3995));
    ClkMux I__719 (
            .O(N__4059),
            .I(N__3995));
    ClkMux I__718 (
            .O(N__4058),
            .I(N__3995));
    ClkMux I__717 (
            .O(N__4057),
            .I(N__3995));
    ClkMux I__716 (
            .O(N__4056),
            .I(N__3995));
    ClkMux I__715 (
            .O(N__4055),
            .I(N__3995));
    ClkMux I__714 (
            .O(N__4054),
            .I(N__3995));
    ClkMux I__713 (
            .O(N__4053),
            .I(N__3995));
    ClkMux I__712 (
            .O(N__4052),
            .I(N__3995));
    ClkMux I__711 (
            .O(N__4051),
            .I(N__3995));
    ClkMux I__710 (
            .O(N__4050),
            .I(N__3995));
    GlobalMux I__709 (
            .O(N__3995),
            .I(N__3992));
    gio2CtrlBuf I__708 (
            .O(N__3992),
            .I(CLK40_c_g));
    InMux I__707 (
            .O(N__3989),
            .I(N__3986));
    LocalMux I__706 (
            .O(N__3986),
            .I(\U400_SDRAM.N_189 ));
    InMux I__705 (
            .O(N__3983),
            .I(N__3977));
    InMux I__704 (
            .O(N__3982),
            .I(N__3974));
    CascadeMux I__703 (
            .O(N__3981),
            .I(N__3971));
    InMux I__702 (
            .O(N__3980),
            .I(N__3962));
    LocalMux I__701 (
            .O(N__3977),
            .I(N__3959));
    LocalMux I__700 (
            .O(N__3974),
            .I(N__3956));
    InMux I__699 (
            .O(N__3971),
            .I(N__3953));
    InMux I__698 (
            .O(N__3970),
            .I(N__3943));
    InMux I__697 (
            .O(N__3969),
            .I(N__3943));
    InMux I__696 (
            .O(N__3968),
            .I(N__3943));
    InMux I__695 (
            .O(N__3967),
            .I(N__3943));
    CascadeMux I__694 (
            .O(N__3966),
            .I(N__3937));
    CascadeMux I__693 (
            .O(N__3965),
            .I(N__3933));
    LocalMux I__692 (
            .O(N__3962),
            .I(N__3927));
    Span4Mux_v I__691 (
            .O(N__3959),
            .I(N__3920));
    Span4Mux_v I__690 (
            .O(N__3956),
            .I(N__3920));
    LocalMux I__689 (
            .O(N__3953),
            .I(N__3920));
    InMux I__688 (
            .O(N__3952),
            .I(N__3917));
    LocalMux I__687 (
            .O(N__3943),
            .I(N__3914));
    InMux I__686 (
            .O(N__3942),
            .I(N__3911));
    InMux I__685 (
            .O(N__3941),
            .I(N__3908));
    InMux I__684 (
            .O(N__3940),
            .I(N__3903));
    InMux I__683 (
            .O(N__3937),
            .I(N__3903));
    InMux I__682 (
            .O(N__3936),
            .I(N__3896));
    InMux I__681 (
            .O(N__3933),
            .I(N__3896));
    InMux I__680 (
            .O(N__3932),
            .I(N__3896));
    InMux I__679 (
            .O(N__3931),
            .I(N__3893));
    InMux I__678 (
            .O(N__3930),
            .I(N__3890));
    Span4Mux_v I__677 (
            .O(N__3927),
            .I(N__3887));
    Span4Mux_h I__676 (
            .O(N__3920),
            .I(N__3882));
    LocalMux I__675 (
            .O(N__3917),
            .I(N__3882));
    Span4Mux_v I__674 (
            .O(N__3914),
            .I(N__3877));
    LocalMux I__673 (
            .O(N__3911),
            .I(N__3877));
    LocalMux I__672 (
            .O(N__3908),
            .I(N__3870));
    LocalMux I__671 (
            .O(N__3903),
            .I(N__3870));
    LocalMux I__670 (
            .O(N__3896),
            .I(N__3870));
    LocalMux I__669 (
            .O(N__3893),
            .I(N__3865));
    LocalMux I__668 (
            .O(N__3890),
            .I(N__3865));
    Span4Mux_h I__667 (
            .O(N__3887),
            .I(N__3860));
    Span4Mux_v I__666 (
            .O(N__3882),
            .I(N__3860));
    Span4Mux_v I__665 (
            .O(N__3877),
            .I(N__3857));
    Span4Mux_v I__664 (
            .O(N__3870),
            .I(N__3854));
    Span12Mux_s8_v I__663 (
            .O(N__3865),
            .I(N__3851));
    Span4Mux_h I__662 (
            .O(N__3860),
            .I(N__3848));
    Span4Mux_h I__661 (
            .O(N__3857),
            .I(N__3845));
    Span4Mux_h I__660 (
            .O(N__3854),
            .I(N__3842));
    Odrv12 I__659 (
            .O(N__3851),
            .I(RESETn_c));
    Odrv4 I__658 (
            .O(N__3848),
            .I(RESETn_c));
    Odrv4 I__657 (
            .O(N__3845),
            .I(RESETn_c));
    Odrv4 I__656 (
            .O(N__3842),
            .I(RESETn_c));
    InMux I__655 (
            .O(N__3833),
            .I(N__3830));
    LocalMux I__654 (
            .O(N__3830),
            .I(N__3826));
    InMux I__653 (
            .O(N__3829),
            .I(N__3823));
    Odrv4 I__652 (
            .O(N__3826),
            .I(\U400_SDRAM.un1_REFRESH_COUNTERlto7_5 ));
    LocalMux I__651 (
            .O(N__3823),
            .I(\U400_SDRAM.un1_REFRESH_COUNTERlto7_5 ));
    InMux I__650 (
            .O(N__3818),
            .I(N__3815));
    LocalMux I__649 (
            .O(N__3815),
            .I(N__3811));
    InMux I__648 (
            .O(N__3814),
            .I(N__3808));
    Odrv4 I__647 (
            .O(N__3811),
            .I(\U400_SDRAM.un1_REFRESH_COUNTERlto7_4 ));
    LocalMux I__646 (
            .O(N__3808),
            .I(\U400_SDRAM.un1_REFRESH_COUNTERlto7_4 ));
    CascadeMux I__645 (
            .O(N__3803),
            .I(N__3800));
    InMux I__644 (
            .O(N__3800),
            .I(N__3796));
    InMux I__643 (
            .O(N__3799),
            .I(N__3793));
    LocalMux I__642 (
            .O(N__3796),
            .I(N__3789));
    LocalMux I__641 (
            .O(N__3793),
            .I(N__3786));
    InMux I__640 (
            .O(N__3792),
            .I(N__3783));
    Span4Mux_h I__639 (
            .O(N__3789),
            .I(N__3778));
    Span4Mux_h I__638 (
            .O(N__3786),
            .I(N__3778));
    LocalMux I__637 (
            .O(N__3783),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_8 ));
    Odrv4 I__636 (
            .O(N__3778),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_8 ));
    IoInMux I__635 (
            .O(N__3773),
            .I(N__3770));
    LocalMux I__634 (
            .O(N__3770),
            .I(N__3766));
    CascadeMux I__633 (
            .O(N__3769),
            .I(N__3763));
    Span12Mux_s5_h I__632 (
            .O(N__3766),
            .I(N__3760));
    InMux I__631 (
            .O(N__3763),
            .I(N__3757));
    Odrv12 I__630 (
            .O(N__3760),
            .I(TA_OUT));
    LocalMux I__629 (
            .O(N__3757),
            .I(TA_OUT));
    IoInMux I__628 (
            .O(N__3752),
            .I(N__3749));
    LocalMux I__627 (
            .O(N__3749),
            .I(N__3746));
    Odrv4 I__626 (
            .O(N__3746),
            .I(N_66));
    CascadeMux I__625 (
            .O(N__3743),
            .I(N__3740));
    InMux I__624 (
            .O(N__3740),
            .I(N__3735));
    InMux I__623 (
            .O(N__3739),
            .I(N__3732));
    InMux I__622 (
            .O(N__3738),
            .I(N__3729));
    LocalMux I__621 (
            .O(N__3735),
            .I(\U400_SDRAM.BURSTZ0 ));
    LocalMux I__620 (
            .O(N__3732),
            .I(\U400_SDRAM.BURSTZ0 ));
    LocalMux I__619 (
            .O(N__3729),
            .I(\U400_SDRAM.BURSTZ0 ));
    InMux I__618 (
            .O(N__3722),
            .I(N__3719));
    LocalMux I__617 (
            .O(N__3719),
            .I(\U400_SDRAM.TA_EN11_m ));
    CascadeMux I__616 (
            .O(N__3716),
            .I(\U400_SDRAM.un1_TA_COUNTER26_0_cascade_ ));
    InMux I__615 (
            .O(N__3713),
            .I(N__3710));
    LocalMux I__614 (
            .O(N__3710),
            .I(\U400_SDRAM.un1_TA_COUNTER26_2_0 ));
    InMux I__613 (
            .O(N__3707),
            .I(N__3703));
    InMux I__612 (
            .O(N__3706),
            .I(N__3700));
    LocalMux I__611 (
            .O(N__3703),
            .I(\U400_SDRAM.TA_COUNTER27 ));
    LocalMux I__610 (
            .O(N__3700),
            .I(\U400_SDRAM.TA_COUNTER27 ));
    InMux I__609 (
            .O(N__3695),
            .I(N__3692));
    LocalMux I__608 (
            .O(N__3692),
            .I(\U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0 ));
    InMux I__607 (
            .O(N__3689),
            .I(N__3686));
    LocalMux I__606 (
            .O(N__3686),
            .I(N__3683));
    Odrv4 I__605 (
            .O(N__3683),
            .I(\U400_SDRAM.N_207 ));
    CascadeMux I__604 (
            .O(N__3680),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_5_1_cascade_ ));
    CascadeMux I__603 (
            .O(N__3677),
            .I(N__3674));
    InMux I__602 (
            .O(N__3674),
            .I(N__3671));
    LocalMux I__601 (
            .O(N__3671),
            .I(\U400_SDRAM.N_250 ));
    CascadeMux I__600 (
            .O(N__3668),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_0_31_i_i_i_2_cascade_ ));
    CascadeMux I__599 (
            .O(N__3665),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_0_31_i_i_i_3_cascade_ ));
    InMux I__598 (
            .O(N__3662),
            .I(N__3658));
    InMux I__597 (
            .O(N__3661),
            .I(N__3655));
    LocalMux I__596 (
            .O(N__3658),
            .I(\U400_SDRAM.N_261 ));
    LocalMux I__595 (
            .O(N__3655),
            .I(\U400_SDRAM.N_261 ));
    InMux I__594 (
            .O(N__3650),
            .I(N__3644));
    InMux I__593 (
            .O(N__3649),
            .I(N__3644));
    LocalMux I__592 (
            .O(N__3644),
            .I(\U400_SDRAM.N_140 ));
    InMux I__591 (
            .O(N__3641),
            .I(N__3638));
    LocalMux I__590 (
            .O(N__3638),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_4_1 ));
    CascadeMux I__589 (
            .O(N__3635),
            .I(N__3632));
    InMux I__588 (
            .O(N__3632),
            .I(N__3628));
    InMux I__587 (
            .O(N__3631),
            .I(N__3625));
    LocalMux I__586 (
            .O(N__3628),
            .I(N__3622));
    LocalMux I__585 (
            .O(N__3625),
            .I(N__3619));
    Odrv4 I__584 (
            .O(N__3622),
            .I(\U400_SDRAM.CS1_ENZ0 ));
    Odrv4 I__583 (
            .O(N__3619),
            .I(\U400_SDRAM.CS1_ENZ0 ));
    IoInMux I__582 (
            .O(N__3614),
            .I(N__3611));
    LocalMux I__581 (
            .O(N__3611),
            .I(N__3608));
    Odrv12 I__580 (
            .O(N__3608),
            .I(CS1n_c));
    CascadeMux I__579 (
            .O(N__3605),
            .I(N__3602));
    InMux I__578 (
            .O(N__3602),
            .I(N__3599));
    LocalMux I__577 (
            .O(N__3599),
            .I(N__3596));
    Span4Mux_v I__576 (
            .O(N__3596),
            .I(N__3593));
    Span4Mux_v I__575 (
            .O(N__3593),
            .I(N__3590));
    IoSpan4Mux I__574 (
            .O(N__3590),
            .I(N__3587));
    Odrv4 I__573 (
            .O(N__3587),
            .I(A_c_26));
    IoInMux I__572 (
            .O(N__3584),
            .I(N__3581));
    LocalMux I__571 (
            .O(N__3581),
            .I(N__3578));
    Odrv12 I__570 (
            .O(N__3578),
            .I(MA_c_12));
    CascadeMux I__569 (
            .O(N__3575),
            .I(\U400_SDRAM.N_236_cascade_ ));
    InMux I__568 (
            .O(N__3572),
            .I(N__3563));
    InMux I__567 (
            .O(N__3571),
            .I(N__3563));
    InMux I__566 (
            .O(N__3570),
            .I(N__3563));
    LocalMux I__565 (
            .O(N__3563),
            .I(\U400_SDRAM.N_23_i ));
    CascadeMux I__564 (
            .O(N__3560),
            .I(\U400_SDRAM.N_23_i_cascade_ ));
    InMux I__563 (
            .O(N__3557),
            .I(N__3554));
    LocalMux I__562 (
            .O(N__3554),
            .I(\U400_SDRAM.N_242 ));
    InMux I__561 (
            .O(N__3551),
            .I(N__3545));
    InMux I__560 (
            .O(N__3550),
            .I(N__3545));
    LocalMux I__559 (
            .O(N__3545),
            .I(\U400_SDRAM.N_139 ));
    InMux I__558 (
            .O(N__3542),
            .I(N__3539));
    LocalMux I__557 (
            .O(N__3539),
            .I(N__3536));
    Span4Mux_h I__556 (
            .O(N__3536),
            .I(N__3533));
    Odrv4 I__555 (
            .O(N__3533),
            .I(\U400_SDRAM.SDRAM_COUNTER_s_1 ));
    CascadeMux I__554 (
            .O(N__3530),
            .I(N__3527));
    InMux I__553 (
            .O(N__3527),
            .I(N__3524));
    LocalMux I__552 (
            .O(N__3524),
            .I(\U400_SDRAM.N_198 ));
    InMux I__551 (
            .O(N__3521),
            .I(N__3515));
    InMux I__550 (
            .O(N__3520),
            .I(N__3515));
    LocalMux I__549 (
            .O(N__3515),
            .I(\U400_SDRAM.N_259 ));
    CascadeMux I__548 (
            .O(N__3512),
            .I(N__3508));
    InMux I__547 (
            .O(N__3511),
            .I(N__3503));
    InMux I__546 (
            .O(N__3508),
            .I(N__3503));
    LocalMux I__545 (
            .O(N__3503),
            .I(\U400_SDRAM.N_118 ));
    CascadeMux I__544 (
            .O(N__3500),
            .I(N__3493));
    InMux I__543 (
            .O(N__3499),
            .I(N__3487));
    InMux I__542 (
            .O(N__3498),
            .I(N__3480));
    InMux I__541 (
            .O(N__3497),
            .I(N__3480));
    InMux I__540 (
            .O(N__3496),
            .I(N__3480));
    InMux I__539 (
            .O(N__3493),
            .I(N__3475));
    InMux I__538 (
            .O(N__3492),
            .I(N__3475));
    InMux I__537 (
            .O(N__3491),
            .I(N__3470));
    InMux I__536 (
            .O(N__3490),
            .I(N__3470));
    LocalMux I__535 (
            .O(N__3487),
            .I(N__3467));
    LocalMux I__534 (
            .O(N__3480),
            .I(\U400_SDRAM.N_39 ));
    LocalMux I__533 (
            .O(N__3475),
            .I(\U400_SDRAM.N_39 ));
    LocalMux I__532 (
            .O(N__3470),
            .I(\U400_SDRAM.N_39 ));
    Odrv4 I__531 (
            .O(N__3467),
            .I(\U400_SDRAM.N_39 ));
    InMux I__530 (
            .O(N__3458),
            .I(N__3455));
    LocalMux I__529 (
            .O(N__3455),
            .I(N__3452));
    Span4Mux_h I__528 (
            .O(N__3452),
            .I(N__3449));
    Odrv4 I__527 (
            .O(N__3449),
            .I(\U400_SDRAM.SDRAM_COUNTER_s_3 ));
    CEMux I__526 (
            .O(N__3446),
            .I(N__3441));
    CEMux I__525 (
            .O(N__3445),
            .I(N__3438));
    CEMux I__524 (
            .O(N__3444),
            .I(N__3435));
    LocalMux I__523 (
            .O(N__3441),
            .I(\U400_SDRAM.N_219_i ));
    LocalMux I__522 (
            .O(N__3438),
            .I(\U400_SDRAM.N_219_i ));
    LocalMux I__521 (
            .O(N__3435),
            .I(\U400_SDRAM.N_219_i ));
    InMux I__520 (
            .O(N__3428),
            .I(N__3425));
    LocalMux I__519 (
            .O(N__3425),
            .I(N__3422));
    Span4Mux_h I__518 (
            .O(N__3422),
            .I(N__3416));
    InMux I__517 (
            .O(N__3421),
            .I(N__3413));
    InMux I__516 (
            .O(N__3420),
            .I(N__3410));
    InMux I__515 (
            .O(N__3419),
            .I(N__3407));
    Odrv4 I__514 (
            .O(N__3416),
            .I(\U400_SDRAM.N_239 ));
    LocalMux I__513 (
            .O(N__3413),
            .I(\U400_SDRAM.N_239 ));
    LocalMux I__512 (
            .O(N__3410),
            .I(\U400_SDRAM.N_239 ));
    LocalMux I__511 (
            .O(N__3407),
            .I(\U400_SDRAM.N_239 ));
    CascadeMux I__510 (
            .O(N__3398),
            .I(N__3395));
    InMux I__509 (
            .O(N__3395),
            .I(N__3392));
    LocalMux I__508 (
            .O(N__3392),
            .I(N__3389));
    Span4Mux_v I__507 (
            .O(N__3389),
            .I(N__3386));
    Sp12to4 I__506 (
            .O(N__3386),
            .I(N__3383));
    Odrv12 I__505 (
            .O(N__3383),
            .I(A_c_21));
    IoInMux I__504 (
            .O(N__3380),
            .I(N__3377));
    LocalMux I__503 (
            .O(N__3377),
            .I(N__3374));
    IoSpan4Mux I__502 (
            .O(N__3374),
            .I(N__3371));
    Span4Mux_s3_h I__501 (
            .O(N__3371),
            .I(N__3368));
    Span4Mux_v I__500 (
            .O(N__3368),
            .I(N__3364));
    InMux I__499 (
            .O(N__3367),
            .I(N__3361));
    Odrv4 I__498 (
            .O(N__3364),
            .I(BANK0_c));
    LocalMux I__497 (
            .O(N__3361),
            .I(BANK0_c));
    CascadeMux I__496 (
            .O(N__3356),
            .I(N__3353));
    InMux I__495 (
            .O(N__3353),
            .I(N__3350));
    LocalMux I__494 (
            .O(N__3350),
            .I(N__3347));
    Span12Mux_s9_h I__493 (
            .O(N__3347),
            .I(N__3344));
    Odrv12 I__492 (
            .O(N__3344),
            .I(A_c_22));
    InMux I__491 (
            .O(N__3341),
            .I(N__3337));
    InMux I__490 (
            .O(N__3340),
            .I(N__3334));
    LocalMux I__489 (
            .O(N__3337),
            .I(\U400_SDRAM.N_240 ));
    LocalMux I__488 (
            .O(N__3334),
            .I(\U400_SDRAM.N_240 ));
    IoInMux I__487 (
            .O(N__3329),
            .I(N__3326));
    LocalMux I__486 (
            .O(N__3326),
            .I(N__3323));
    IoSpan4Mux I__485 (
            .O(N__3323),
            .I(N__3320));
    IoSpan4Mux I__484 (
            .O(N__3320),
            .I(N__3317));
    Span4Mux_s3_h I__483 (
            .O(N__3317),
            .I(N__3313));
    InMux I__482 (
            .O(N__3316),
            .I(N__3310));
    Odrv4 I__481 (
            .O(N__3313),
            .I(BANK1_c));
    LocalMux I__480 (
            .O(N__3310),
            .I(BANK1_c));
    InMux I__479 (
            .O(N__3305),
            .I(N__3302));
    LocalMux I__478 (
            .O(N__3302),
            .I(N__3299));
    Span12Mux_v I__477 (
            .O(N__3299),
            .I(N__3296));
    Odrv12 I__476 (
            .O(N__3296),
            .I(RnW_c));
    InMux I__475 (
            .O(N__3293),
            .I(N__3290));
    LocalMux I__474 (
            .O(N__3290),
            .I(\U400_SDRAM.N_82 ));
    InMux I__473 (
            .O(N__3287),
            .I(N__3284));
    LocalMux I__472 (
            .O(N__3284),
            .I(\U400_SDRAM.N_34 ));
    CascadeMux I__471 (
            .O(N__3281),
            .I(\U400_SDRAM.N_118_cascade_ ));
    InMux I__470 (
            .O(N__3278),
            .I(N__3275));
    LocalMux I__469 (
            .O(N__3275),
            .I(\U400_SDRAM.N_215 ));
    InMux I__468 (
            .O(N__3272),
            .I(N__3268));
    InMux I__467 (
            .O(N__3271),
            .I(N__3265));
    LocalMux I__466 (
            .O(N__3268),
            .I(\U400_SDRAM.RAM_CYCLEZ0 ));
    LocalMux I__465 (
            .O(N__3265),
            .I(\U400_SDRAM.RAM_CYCLEZ0 ));
    InMux I__464 (
            .O(N__3260),
            .I(N__3251));
    InMux I__463 (
            .O(N__3259),
            .I(N__3251));
    InMux I__462 (
            .O(N__3258),
            .I(N__3251));
    LocalMux I__461 (
            .O(N__3251),
            .I(\U400_SDRAM.SDRAM_CONFIGURED_RNI5POA3Z0Z_0 ));
    CascadeMux I__460 (
            .O(N__3248),
            .I(\U400_SDRAM.N_230_cascade_ ));
    CascadeMux I__459 (
            .O(N__3245),
            .I(N__3242));
    InMux I__458 (
            .O(N__3242),
            .I(N__3239));
    LocalMux I__457 (
            .O(N__3239),
            .I(N__3236));
    Sp12to4 I__456 (
            .O(N__3236),
            .I(N__3233));
    Span12Mux_s10_v I__455 (
            .O(N__3233),
            .I(N__3230));
    Odrv12 I__454 (
            .O(N__3230),
            .I(A_c_19));
    IoInMux I__453 (
            .O(N__3227),
            .I(N__3224));
    LocalMux I__452 (
            .O(N__3224),
            .I(N__3221));
    Odrv12 I__451 (
            .O(N__3221),
            .I(MA_c_9));
    InMux I__450 (
            .O(N__3218),
            .I(N__3215));
    LocalMux I__449 (
            .O(N__3215),
            .I(A_c_30));
    InMux I__448 (
            .O(N__3212),
            .I(N__3209));
    LocalMux I__447 (
            .O(N__3209),
            .I(N__3206));
    Span12Mux_s10_h I__446 (
            .O(N__3206),
            .I(N__3203));
    Odrv12 I__445 (
            .O(N__3203),
            .I(A_c_29));
    CascadeMux I__444 (
            .O(N__3200),
            .I(\U400_SDRAM.TA_COUNTER_0_sqmuxa_cascade_ ));
    InMux I__443 (
            .O(N__3197),
            .I(N__3194));
    LocalMux I__442 (
            .O(N__3194),
            .I(\U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en ));
    CEMux I__441 (
            .O(N__3191),
            .I(N__3188));
    LocalMux I__440 (
            .O(N__3188),
            .I(\U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en_0 ));
    CascadeMux I__439 (
            .O(N__3185),
            .I(\U400_SDRAM.CS0_EN_0_cascade_ ));
    InMux I__438 (
            .O(N__3182),
            .I(N__3178));
    InMux I__437 (
            .O(N__3181),
            .I(N__3175));
    LocalMux I__436 (
            .O(N__3178),
            .I(\U400_SDRAM.CS0_ENZ0 ));
    LocalMux I__435 (
            .O(N__3175),
            .I(\U400_SDRAM.CS0_ENZ0 ));
    CascadeMux I__434 (
            .O(N__3170),
            .I(N__3166));
    CascadeMux I__433 (
            .O(N__3169),
            .I(N__3163));
    InMux I__432 (
            .O(N__3166),
            .I(N__3158));
    InMux I__431 (
            .O(N__3163),
            .I(N__3158));
    LocalMux I__430 (
            .O(N__3158),
            .I(N__3155));
    Span4Mux_v I__429 (
            .O(N__3155),
            .I(N__3152));
    Odrv4 I__428 (
            .O(N__3152),
            .I(A_c_23));
    CascadeMux I__427 (
            .O(N__3149),
            .I(\U400_SDRAM.CS1_EN_0_cascade_ ));
    CascadeMux I__426 (
            .O(N__3146),
            .I(\U400_SDRAM.N_114_cascade_ ));
    InMux I__425 (
            .O(N__3143),
            .I(N__3140));
    LocalMux I__424 (
            .O(N__3140),
            .I(\U400_SDRAM.N_220 ));
    InMux I__423 (
            .O(N__3137),
            .I(N__3134));
    LocalMux I__422 (
            .O(N__3134),
            .I(\U400_SDRAM.N_258 ));
    InMux I__421 (
            .O(N__3131),
            .I(N__3128));
    LocalMux I__420 (
            .O(N__3128),
            .I(\U400_SDRAM.un1_SDRAM_COUNTER52_4_i_0_1 ));
    CascadeMux I__419 (
            .O(N__3125),
            .I(\U400_SDRAM.N_258_cascade_ ));
    InMux I__418 (
            .O(N__3122),
            .I(N__3119));
    LocalMux I__417 (
            .O(N__3119),
            .I(N__3116));
    Span4Mux_h I__416 (
            .O(N__3116),
            .I(N__3113));
    Odrv4 I__415 (
            .O(N__3113),
            .I(\U400_SDRAM.un1_SDRAM_COUNTER52_4_i_0_0 ));
    CascadeMux I__414 (
            .O(N__3110),
            .I(\U400_SDRAM.N_240_cascade_ ));
    InMux I__413 (
            .O(N__3107),
            .I(N__3103));
    InMux I__412 (
            .O(N__3106),
            .I(N__3100));
    LocalMux I__411 (
            .O(N__3103),
            .I(N__3097));
    LocalMux I__410 (
            .O(N__3100),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_3 ));
    Odrv4 I__409 (
            .O(N__3097),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__408 (
            .O(N__3092),
            .I(N__3088));
    InMux I__407 (
            .O(N__3091),
            .I(N__3085));
    LocalMux I__406 (
            .O(N__3088),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_2 ));
    LocalMux I__405 (
            .O(N__3085),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_2 ));
    CascadeMux I__404 (
            .O(N__3080),
            .I(N__3076));
    InMux I__403 (
            .O(N__3079),
            .I(N__3073));
    InMux I__402 (
            .O(N__3076),
            .I(N__3070));
    LocalMux I__401 (
            .O(N__3073),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__400 (
            .O(N__3070),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__399 (
            .O(N__3065),
            .I(N__3060));
    InMux I__398 (
            .O(N__3064),
            .I(N__3055));
    InMux I__397 (
            .O(N__3063),
            .I(N__3055));
    LocalMux I__396 (
            .O(N__3060),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_1 ));
    LocalMux I__395 (
            .O(N__3055),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_1 ));
    InMux I__394 (
            .O(N__3050),
            .I(N__3046));
    InMux I__393 (
            .O(N__3049),
            .I(N__3043));
    LocalMux I__392 (
            .O(N__3046),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__391 (
            .O(N__3043),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__390 (
            .O(N__3038),
            .I(N__3034));
    InMux I__389 (
            .O(N__3037),
            .I(N__3031));
    LocalMux I__388 (
            .O(N__3034),
            .I(N__3028));
    LocalMux I__387 (
            .O(N__3031),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_6 ));
    Odrv4 I__386 (
            .O(N__3028),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_6 ));
    CascadeMux I__385 (
            .O(N__3023),
            .I(N__3019));
    InMux I__384 (
            .O(N__3022),
            .I(N__3016));
    InMux I__383 (
            .O(N__3019),
            .I(N__3013));
    LocalMux I__382 (
            .O(N__3016),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_7 ));
    LocalMux I__381 (
            .O(N__3013),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_7 ));
    CascadeMux I__380 (
            .O(N__3008),
            .I(N__3004));
    CascadeMux I__379 (
            .O(N__3007),
            .I(N__3001));
    InMux I__378 (
            .O(N__3004),
            .I(N__2996));
    InMux I__377 (
            .O(N__3001),
            .I(N__2989));
    InMux I__376 (
            .O(N__3000),
            .I(N__2989));
    InMux I__375 (
            .O(N__2999),
            .I(N__2989));
    LocalMux I__374 (
            .O(N__2996),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_0 ));
    LocalMux I__373 (
            .O(N__2989),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_0 ));
    SRMux I__372 (
            .O(N__2984),
            .I(N__2981));
    LocalMux I__371 (
            .O(N__2981),
            .I(N__2977));
    SRMux I__370 (
            .O(N__2980),
            .I(N__2974));
    Span4Mux_h I__369 (
            .O(N__2977),
            .I(N__2971));
    LocalMux I__368 (
            .O(N__2974),
            .I(\U400_SDRAM.SDRAM_CONFIGURED_RNIJKCAZ0Z2 ));
    Odrv4 I__367 (
            .O(N__2971),
            .I(\U400_SDRAM.SDRAM_CONFIGURED_RNIJKCAZ0Z2 ));
    InMux I__366 (
            .O(N__2966),
            .I(N__2963));
    LocalMux I__365 (
            .O(N__2963),
            .I(N__2960));
    Odrv12 I__364 (
            .O(N__2960),
            .I(A_c_8));
    CascadeMux I__363 (
            .O(N__2957),
            .I(N__2954));
    InMux I__362 (
            .O(N__2954),
            .I(N__2951));
    LocalMux I__361 (
            .O(N__2951),
            .I(N__2948));
    Span4Mux_v I__360 (
            .O(N__2948),
            .I(N__2945));
    Span4Mux_v I__359 (
            .O(N__2945),
            .I(N__2942));
    Odrv4 I__358 (
            .O(N__2942),
            .I(A_c_16));
    IoInMux I__357 (
            .O(N__2939),
            .I(N__2936));
    LocalMux I__356 (
            .O(N__2936),
            .I(N__2933));
    Odrv4 I__355 (
            .O(N__2933),
            .I(MA_c_6));
    InMux I__354 (
            .O(N__2930),
            .I(N__2927));
    LocalMux I__353 (
            .O(N__2927),
            .I(\U400_SDRAM.N_216 ));
    InMux I__352 (
            .O(N__2924),
            .I(N__2921));
    LocalMux I__351 (
            .O(N__2921),
            .I(N__2917));
    InMux I__350 (
            .O(N__2920),
            .I(N__2914));
    Odrv4 I__349 (
            .O(N__2917),
            .I(\U400_SDRAM.N_187 ));
    LocalMux I__348 (
            .O(N__2914),
            .I(\U400_SDRAM.N_187 ));
    InMux I__347 (
            .O(N__2909),
            .I(N__2906));
    LocalMux I__346 (
            .O(N__2906),
            .I(N__2903));
    Odrv4 I__345 (
            .O(N__2903),
            .I(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_2_0 ));
    CascadeMux I__344 (
            .O(N__2900),
            .I(N__2897));
    InMux I__343 (
            .O(N__2897),
            .I(N__2894));
    LocalMux I__342 (
            .O(N__2894),
            .I(\U400_SDRAM.SDRAM_COUNTER_s_0 ));
    InMux I__341 (
            .O(N__2891),
            .I(N__2888));
    LocalMux I__340 (
            .O(N__2888),
            .I(\U400_SDRAM.TACK_7_iv_i_i_2 ));
    CascadeMux I__339 (
            .O(N__2885),
            .I(\U400_SDRAM.TACK_7_iv_i_i_1_0_cascade_ ));
    IoInMux I__338 (
            .O(N__2882),
            .I(N__2879));
    LocalMux I__337 (
            .O(N__2879),
            .I(N__2876));
    Span4Mux_s3_h I__336 (
            .O(N__2876),
            .I(N__2873));
    Odrv4 I__335 (
            .O(N__2873),
            .I(CS0n_c));
    IoInMux I__334 (
            .O(N__2870),
            .I(N__2867));
    LocalMux I__333 (
            .O(N__2867),
            .I(N__2864));
    Odrv12 I__332 (
            .O(N__2864),
            .I(CASn_c));
    IoInMux I__331 (
            .O(N__2861),
            .I(N__2858));
    LocalMux I__330 (
            .O(N__2858),
            .I(N__2855));
    Odrv12 I__329 (
            .O(N__2855),
            .I(WEn_c));
    IoInMux I__328 (
            .O(N__2852),
            .I(N__2849));
    LocalMux I__327 (
            .O(N__2849),
            .I(N__2846));
    Odrv12 I__326 (
            .O(N__2846),
            .I(RASn_c));
    InMux I__325 (
            .O(N__2843),
            .I(N__2840));
    LocalMux I__324 (
            .O(N__2840),
            .I(N__2837));
    Span4Mux_h I__323 (
            .O(N__2837),
            .I(N__2834));
    Sp12to4 I__322 (
            .O(N__2834),
            .I(N__2831));
    Span12Mux_v I__321 (
            .O(N__2831),
            .I(N__2828));
    Odrv12 I__320 (
            .O(N__2828),
            .I(A_c_24));
    CascadeMux I__319 (
            .O(N__2825),
            .I(N__2822));
    InMux I__318 (
            .O(N__2822),
            .I(N__2819));
    LocalMux I__317 (
            .O(N__2819),
            .I(N__2816));
    Span12Mux_s10_v I__316 (
            .O(N__2816),
            .I(N__2813));
    Odrv12 I__315 (
            .O(N__2813),
            .I(A_c_18));
    IoInMux I__314 (
            .O(N__2810),
            .I(N__2807));
    LocalMux I__313 (
            .O(N__2807),
            .I(N__2804));
    Span4Mux_s1_v I__312 (
            .O(N__2804),
            .I(N__2801));
    Odrv4 I__311 (
            .O(N__2801),
            .I(MA_c_8));
    InMux I__310 (
            .O(N__2798),
            .I(N__2795));
    LocalMux I__309 (
            .O(N__2795),
            .I(N__2792));
    Odrv12 I__308 (
            .O(N__2792),
            .I(A_c_9));
    CascadeMux I__307 (
            .O(N__2789),
            .I(N__2786));
    InMux I__306 (
            .O(N__2786),
            .I(N__2783));
    LocalMux I__305 (
            .O(N__2783),
            .I(N__2780));
    Span4Mux_v I__304 (
            .O(N__2780),
            .I(N__2777));
    Odrv4 I__303 (
            .O(N__2777),
            .I(A_c_17));
    IoInMux I__302 (
            .O(N__2774),
            .I(N__2771));
    LocalMux I__301 (
            .O(N__2771),
            .I(N__2768));
    Span4Mux_s1_v I__300 (
            .O(N__2768),
            .I(N__2765));
    Odrv4 I__299 (
            .O(N__2765),
            .I(MA_c_7));
    InMux I__298 (
            .O(N__2762),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_4 ));
    InMux I__297 (
            .O(N__2759),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_5 ));
    InMux I__296 (
            .O(N__2756),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_6 ));
    InMux I__295 (
            .O(N__2753),
            .I(N__2750));
    LocalMux I__294 (
            .O(N__2750),
            .I(N__2747));
    Odrv4 I__293 (
            .O(N__2747),
            .I(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_0_0 ));
    CascadeMux I__292 (
            .O(N__2744),
            .I(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_a2_1_0_cascade_ ));
    InMux I__291 (
            .O(N__2741),
            .I(N__2737));
    InMux I__290 (
            .O(N__2740),
            .I(N__2734));
    LocalMux I__289 (
            .O(N__2737),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__288 (
            .O(N__2734),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__287 (
            .O(N__2729),
            .I(N__2725));
    InMux I__286 (
            .O(N__2728),
            .I(N__2722));
    LocalMux I__285 (
            .O(N__2725),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__284 (
            .O(N__2722),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__283 (
            .O(N__2717),
            .I(N__2713));
    InMux I__282 (
            .O(N__2716),
            .I(N__2710));
    InMux I__281 (
            .O(N__2713),
            .I(N__2707));
    LocalMux I__280 (
            .O(N__2710),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__279 (
            .O(N__2707),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_7 ));
    InMux I__278 (
            .O(N__2702),
            .I(N__2698));
    InMux I__277 (
            .O(N__2701),
            .I(N__2695));
    LocalMux I__276 (
            .O(N__2698),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__275 (
            .O(N__2695),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_4 ));
    CascadeMux I__274 (
            .O(N__2690),
            .I(\U400_SDRAM.N_97_cascade_ ));
    CascadeMux I__273 (
            .O(N__2687),
            .I(\U400_SDRAM.N_256_cascade_ ));
    InMux I__272 (
            .O(N__2684),
            .I(N__2681));
    LocalMux I__271 (
            .O(N__2681),
            .I(N__2677));
    InMux I__270 (
            .O(N__2680),
            .I(N__2674));
    Odrv4 I__269 (
            .O(N__2677),
            .I(\U400_SDRAM.SDRAM_CMD_3_sqmuxa ));
    LocalMux I__268 (
            .O(N__2674),
            .I(\U400_SDRAM.SDRAM_CMD_3_sqmuxa ));
    InMux I__267 (
            .O(N__2669),
            .I(\U400_SDRAM.un2_REFRESH_COUNTER_cry_4 ));
    InMux I__266 (
            .O(N__2666),
            .I(\U400_SDRAM.un2_REFRESH_COUNTER_cry_5 ));
    InMux I__265 (
            .O(N__2663),
            .I(\U400_SDRAM.un2_REFRESH_COUNTER_cry_6 ));
    InMux I__264 (
            .O(N__2660),
            .I(\U400_SDRAM.un2_REFRESH_COUNTER_cry_7 ));
    InMux I__263 (
            .O(N__2657),
            .I(bfn_4_6_0_));
    InMux I__262 (
            .O(N__2654),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_0 ));
    InMux I__261 (
            .O(N__2651),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_1 ));
    InMux I__260 (
            .O(N__2648),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_2 ));
    InMux I__259 (
            .O(N__2645),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_3 ));
    IoInMux I__258 (
            .O(N__2642),
            .I(N__2639));
    LocalMux I__257 (
            .O(N__2639),
            .I(RESETn_c_i));
    IoInMux I__256 (
            .O(N__2636),
            .I(N__2633));
    LocalMux I__255 (
            .O(N__2633),
            .I(CONSTANT_ONE_NET));
    InMux I__254 (
            .O(N__2630),
            .I(N__2627));
    LocalMux I__253 (
            .O(N__2627),
            .I(N__2624));
    Odrv12 I__252 (
            .O(N__2624),
            .I(A_c_27));
    InMux I__251 (
            .O(N__2621),
            .I(N__2618));
    LocalMux I__250 (
            .O(N__2618),
            .I(N__2615));
    Odrv4 I__249 (
            .O(N__2615),
            .I(A_c_28));
    CascadeMux I__248 (
            .O(N__2612),
            .I(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_a2_1_0_0_cascade_ ));
    InMux I__247 (
            .O(N__2609),
            .I(\U400_SDRAM.un2_REFRESH_COUNTER_cry_1 ));
    InMux I__246 (
            .O(N__2606),
            .I(\U400_SDRAM.un2_REFRESH_COUNTER_cry_2 ));
    InMux I__245 (
            .O(N__2603),
            .I(\U400_SDRAM.un2_REFRESH_COUNTER_cry_3 ));
    IoInMux I__244 (
            .O(N__2600),
            .I(N__2597));
    LocalMux I__243 (
            .O(N__2597),
            .I(N__2594));
    IoSpan4Mux I__242 (
            .O(N__2594),
            .I(N__2591));
    IoSpan4Mux I__241 (
            .O(N__2591),
            .I(N__2588));
    Span4Mux_s2_h I__240 (
            .O(N__2588),
            .I(N__2585));
    Sp12to4 I__239 (
            .O(N__2585),
            .I(N__2582));
    Odrv12 I__238 (
            .O(N__2582),
            .I(CLK40_ibuf_gb_io_gb_input));
    INV \INVU400_SDRAM.MA_nesr_2C  (
            .O(\INVU400_SDRAM.MA_nesr_2C_net ),
            .I(N__4076));
    INV \INVU400_SDRAM.MA_nesr_3C  (
            .O(\INVU400_SDRAM.MA_nesr_3C_net ),
            .I(N__4075));
    INV \INVU400_SDRAM.MA_nesr_10C  (
            .O(\INVU400_SDRAM.MA_nesr_10C_net ),
            .I(N__4072));
    INV \INVU400_SDRAM.MA_nesr_5C  (
            .O(\INVU400_SDRAM.MA_nesr_5C_net ),
            .I(N__4073));
    INV \INVU400_SDRAM.MA_nesr_11C  (
            .O(\INVU400_SDRAM.MA_nesr_11C_net ),
            .I(N__4069));
    INV \INVU400_SDRAM.SDRAM_CMD_ne_0C  (
            .O(\INVU400_SDRAM.SDRAM_CMD_ne_0C_net ),
            .I(N__4062));
    INV \INVU400_SDRAM.MA_nesr_12C  (
            .O(\INVU400_SDRAM.MA_nesr_12C_net ),
            .I(N__4066));
    INV \INVU400_SDRAM.CS1nC  (
            .O(\INVU400_SDRAM.CS1nC_net ),
            .I(N__4053));
    INV \INVU400_SDRAM.SDRAM_CMD_1C  (
            .O(\INVU400_SDRAM.SDRAM_CMD_1C_net ),
            .I(N__4057));
    INV \INVU400_SDRAM.SDRAM_COUNTER_1C  (
            .O(\INVU400_SDRAM.SDRAM_COUNTER_1C_net ),
            .I(N__4061));
    INV \INVU400_SDRAM.BANK0C  (
            .O(\INVU400_SDRAM.BANK0C_net ),
            .I(N__4068));
    INV \INVU400_SDRAM.MA_nesr_9C  (
            .O(\INVU400_SDRAM.MA_nesr_9C_net ),
            .I(N__4059));
    INV \INVU400_SDRAM.CS0_ENC  (
            .O(\INVU400_SDRAM.CS0_ENC_net ),
            .I(N__4056));
    INV \INVU400_SDRAM.REFRESH_COUNTER_1C  (
            .O(\INVU400_SDRAM.REFRESH_COUNTER_1C_net ),
            .I(N__4060));
    INV \INVU400_SDRAM.SDRAM_COUNTER_0C  (
            .O(\INVU400_SDRAM.SDRAM_COUNTER_0C_net ),
            .I(N__4065));
    INV \INVU400_SDRAM.MA_nesr_6C  (
            .O(\INVU400_SDRAM.MA_nesr_6C_net ),
            .I(N__4063));
    INV \INVU400_SDRAM.MA_nesr_8C  (
            .O(\INVU400_SDRAM.MA_nesr_8C_net ),
            .I(N__4054));
    INV \INVU400_SDRAM.RASnC  (
            .O(\INVU400_SDRAM.RASnC_net ),
            .I(N__4051));
    INV \INVU400_SDRAM.CASnC  (
            .O(\INVU400_SDRAM.CASnC_net ),
            .I(N__4050));
    INV \INVU400_SDRAM.CS0nC  (
            .O(\INVU400_SDRAM.CS0nC_net ),
            .I(N__4052));
    INV \INVU400_SDRAM.SDRAM_COUNTER_2C  (
            .O(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .I(N__4055));
    INV \INVU400_SDRAM.REFRESH_COUNTER_2C  (
            .O(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .I(N__4058));
    INV \INVU400_SDRAM.SDRAM_CONFIGUREDC  (
            .O(\INVU400_SDRAM.SDRAM_CONFIGUREDC_net ),
            .I(N__4064));
    defparam IN_MUX_bfv_4_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_5_0_));
    defparam IN_MUX_bfv_4_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_6_0_));
    ICE_GB CLK40_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__2600),
            .GLOBALBUFFEROUTPUT(CLK40_c_g));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__2642),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_1_8_6.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_1_8_6.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_1_8_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_1_8_6 (
            .in0(N__3980),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_1_14_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_1_14_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_1_14_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_1_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_0_o2_2_LC_4_2_5 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_0_o2_2_LC_4_2_5 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_0_o2_2_LC_4_2_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_0_o2_2_LC_4_2_5  (
            .in0(N__2630),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2621),
            .lcout(U400_ADDRESS_DECODE_RAM_SPACE_i_o3_0_o2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_LC_4_4_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_LC_4_4_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_LC_4_4_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_LC_4_4_1  (
            .in0(_gnd_net_),
            .in1(N__5457),
            .in2(_gnd_net_),
            .in3(N__2684),
            .lcout(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_CONFIGUREDC_net ),
            .ce(),
            .sr(N__6163));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_5_0_LC_4_4_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_5_0_LC_4_4_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_5_0_LC_4_4_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_5_0_LC_4_4_4  (
            .in0(N__4817),
            .in1(N__4617),
            .in2(_gnd_net_),
            .in3(N__4898),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_a2_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_3_0_LC_4_4_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_3_0_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_3_0_LC_4_4_5 .LUT_INIT=16'b0101010111010101;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_3_0_LC_4_4_5  (
            .in0(N__3931),
            .in1(N__5456),
            .in2(N__2612),
            .in3(N__4349),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.un2_REFRESH_COUNTER_cry_1_c_LC_4_5_0 .C_ON=1'b1;
    defparam \U400_SDRAM.un2_REFRESH_COUNTER_cry_1_c_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.un2_REFRESH_COUNTER_cry_1_c_LC_4_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U400_SDRAM.un2_REFRESH_COUNTER_cry_1_c_LC_4_5_0  (
            .in0(_gnd_net_),
            .in1(N__3065),
            .in2(N__3008),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_5_0_),
            .carryout(\U400_SDRAM.un2_REFRESH_COUNTER_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_2_LC_4_5_1 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_2_LC_4_5_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_2_LC_4_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_2_LC_4_5_1  (
            .in0(_gnd_net_),
            .in1(N__3092),
            .in2(_gnd_net_),
            .in3(N__2609),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U400_SDRAM.un2_REFRESH_COUNTER_cry_1 ),
            .carryout(\U400_SDRAM.un2_REFRESH_COUNTER_cry_2 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__2984));
    defparam \U400_SDRAM.REFRESH_COUNTER_3_LC_4_5_2 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_3_LC_4_5_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_3_LC_4_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_3_LC_4_5_2  (
            .in0(_gnd_net_),
            .in1(N__3106),
            .in2(_gnd_net_),
            .in3(N__2606),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U400_SDRAM.un2_REFRESH_COUNTER_cry_2 ),
            .carryout(\U400_SDRAM.un2_REFRESH_COUNTER_cry_3 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__2984));
    defparam \U400_SDRAM.REFRESH_COUNTER_4_LC_4_5_3 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_4_LC_4_5_3 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_4_LC_4_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_4_LC_4_5_3  (
            .in0(_gnd_net_),
            .in1(N__3079),
            .in2(_gnd_net_),
            .in3(N__2603),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U400_SDRAM.un2_REFRESH_COUNTER_cry_3 ),
            .carryout(\U400_SDRAM.un2_REFRESH_COUNTER_cry_4 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__2984));
    defparam \U400_SDRAM.REFRESH_COUNTER_5_LC_4_5_4 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_5_LC_4_5_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_5_LC_4_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_5_LC_4_5_4  (
            .in0(_gnd_net_),
            .in1(N__3050),
            .in2(_gnd_net_),
            .in3(N__2669),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U400_SDRAM.un2_REFRESH_COUNTER_cry_4 ),
            .carryout(\U400_SDRAM.un2_REFRESH_COUNTER_cry_5 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__2984));
    defparam \U400_SDRAM.REFRESH_COUNTER_6_LC_4_5_5 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_6_LC_4_5_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_6_LC_4_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_6_LC_4_5_5  (
            .in0(_gnd_net_),
            .in1(N__3037),
            .in2(_gnd_net_),
            .in3(N__2666),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U400_SDRAM.un2_REFRESH_COUNTER_cry_5 ),
            .carryout(\U400_SDRAM.un2_REFRESH_COUNTER_cry_6 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__2984));
    defparam \U400_SDRAM.REFRESH_COUNTER_7_LC_4_5_6 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_7_LC_4_5_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_7_LC_4_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_7_LC_4_5_6  (
            .in0(_gnd_net_),
            .in1(N__3022),
            .in2(_gnd_net_),
            .in3(N__2663),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(\U400_SDRAM.un2_REFRESH_COUNTER_cry_6 ),
            .carryout(\U400_SDRAM.un2_REFRESH_COUNTER_cry_7 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__2984));
    defparam \U400_SDRAM.REFRESH_COUNTER_8_LC_4_5_7 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_8_LC_4_5_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_8_LC_4_5_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_8_LC_4_5_7  (
            .in0(_gnd_net_),
            .in1(N__3792),
            .in2(_gnd_net_),
            .in3(N__2660),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__2984));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_2_0_LC_4_6_0 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_2_0_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_2_0_LC_4_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_2_0_LC_4_6_0  (
            .in0(_gnd_net_),
            .in1(N__4907),
            .in2(_gnd_net_),
            .in3(N__2657),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(bfn_4_6_0_),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_4_6_1 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_4_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_4_6_1  (
            .in0(_gnd_net_),
            .in1(N__4819),
            .in2(_gnd_net_),
            .in3(N__2654),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_s_1 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_2_LC_4_6_2 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_2_LC_4_6_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_2_LC_4_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_2_LC_4_6_2  (
            .in0(N__3496),
            .in1(N__4462),
            .in2(_gnd_net_),
            .in3(N__2651),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_2 ),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__3444),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_4_6_3 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_4_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_4_6_3  (
            .in0(_gnd_net_),
            .in1(N__4618),
            .in2(_gnd_net_),
            .in3(N__2648),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_s_3 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_4_LC_4_6_4 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_4_LC_4_6_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_4_LC_4_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_4_LC_4_6_4  (
            .in0(N__3497),
            .in1(N__2702),
            .in2(_gnd_net_),
            .in3(N__2645),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_4 ),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__3444),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_5_LC_4_6_5 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_5_LC_4_6_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_5_LC_4_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_5_LC_4_6_5  (
            .in0(N__3490),
            .in1(N__2729),
            .in2(_gnd_net_),
            .in3(N__2762),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_5 ),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__3444),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_6_LC_4_6_6 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_6_LC_4_6_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_6_LC_4_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_6_LC_4_6_6  (
            .in0(N__3498),
            .in1(N__2741),
            .in2(_gnd_net_),
            .in3(N__2759),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_6 ),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__3444),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_7_LC_4_6_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_7_LC_4_6_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_7_LC_4_6_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_7_LC_4_6_7  (
            .in0(N__3491),
            .in1(N__2716),
            .in2(_gnd_net_),
            .in3(N__2756),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__3444),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_4_0_LC_4_7_0 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_4_0_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_4_0_LC_4_7_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_4_0_LC_4_7_0  (
            .in0(N__5516),
            .in1(N__2924),
            .in2(_gnd_net_),
            .in3(N__4444),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_a2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_1_0_LC_4_7_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_1_0_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_1_0_LC_4_7_1 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_1_0_LC_4_7_1  (
            .in0(N__2753),
            .in1(N__3420),
            .in2(N__2744),
            .in3(N__2680),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_4_7_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_4_7_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_4_7_2  (
            .in0(N__2740),
            .in1(N__2728),
            .in2(N__2717),
            .in3(N__2701),
            .lcout(\U400_SDRAM.N_97 ),
            .ltout(\U400_SDRAM.N_97_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_0_2_LC_4_7_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_0_2_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_0_2_LC_4_7_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_0_2_LC_4_7_3  (
            .in0(N__4442),
            .in1(N__4598),
            .in2(N__2690),
            .in3(N__4926),
            .lcout(\U400_SDRAM.N_256 ),
            .ltout(\U400_SDRAM.N_256_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNITAGQ1_LC_4_7_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNITAGQ1_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNITAGQ1_LC_4_7_4 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNITAGQ1_LC_4_7_4  (
            .in0(_gnd_net_),
            .in1(N__5523),
            .in2(N__2687),
            .in3(N__4808),
            .lcout(\U400_SDRAM.SDRAM_CMD_3_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIJKCA2_LC_4_7_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIJKCA2_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIJKCA2_LC_4_7_5 .LUT_INIT=16'b0011001110110011;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNIJKCA2_LC_4_7_5  (
            .in0(N__4809),
            .in1(N__3930),
            .in2(N__5547),
            .in3(N__5396),
            .lcout(\U400_SDRAM.SDRAM_CONFIGURED_RNIJKCAZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_2_LC_4_7_6 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_2_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_2_LC_4_7_6 .LUT_INIT=16'b1111101110111011;
    LogicCell40 \U400_SDRAM.TACK_RNO_2_LC_4_7_6  (
            .in0(N__4337),
            .in1(N__5522),
            .in2(N__4616),
            .in3(N__4443),
            .lcout(\U400_SDRAM.un1_SDRAM_COUNTER52_4_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIE9F21_1_LC_4_7_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIE9F21_1_LC_4_7_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIE9F21_1_LC_4_7_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIE9F21_1_LC_4_7_7  (
            .in0(N__4807),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4336),
            .lcout(\U400_SDRAM.N_239 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.CS0n_LC_4_8_0 .C_ON=1'b0;
    defparam \U400_SDRAM.CS0n_LC_4_8_0 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.CS0n_LC_4_8_0 .LUT_INIT=16'b1000000011111111;
    LogicCell40 \U400_SDRAM.CS0n_LC_4_8_0  (
            .in0(N__6450),
            .in1(N__6067),
            .in2(N__5969),
            .in3(N__3182),
            .lcout(CS0n_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS0nC_net ),
            .ce(),
            .sr(N__6157));
    defparam \U400_SDRAM.CASn_LC_4_9_3 .C_ON=1'b0;
    defparam \U400_SDRAM.CASn_LC_4_9_3 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.CASn_LC_4_9_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U400_SDRAM.CASn_LC_4_9_3  (
            .in0(N__6069),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CASnC_net ),
            .ce(),
            .sr(N__6158));
    defparam \U400_SDRAM.WEn_LC_4_9_6 .C_ON=1'b0;
    defparam \U400_SDRAM.WEn_LC_4_9_6 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.WEn_LC_4_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U400_SDRAM.WEn_LC_4_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5967),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CASnC_net ),
            .ce(),
            .sr(N__6158));
    defparam \U400_SDRAM.RASn_LC_4_10_0 .C_ON=1'b0;
    defparam \U400_SDRAM.RASn_LC_4_10_0 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.RASn_LC_4_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U400_SDRAM.RASn_LC_4_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6489),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.RASnC_net ),
            .ce(),
            .sr(N__6159));
    defparam \U400_SDRAM.MA_nesr_8_LC_4_12_2 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_8_LC_4_12_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_8_LC_4_12_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U400_SDRAM.MA_nesr_8_LC_4_12_2  (
            .in0(N__6491),
            .in1(N__2843),
            .in2(N__2825),
            .in3(N__6332),
            .lcout(MA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_8C_net ),
            .ce(N__6268),
            .sr(N__6162));
    defparam \U400_SDRAM.MA_nesr_7_LC_4_12_4 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_7_LC_4_12_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_7_LC_4_12_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U400_SDRAM.MA_nesr_7_LC_4_12_4  (
            .in0(N__6490),
            .in1(N__2798),
            .in2(N__2789),
            .in3(N__6331),
            .lcout(MA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_8C_net ),
            .ce(N__6268),
            .sr(N__6162));
    defparam \U400_SDRAM.MA_nesr_6_LC_4_14_3 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_6_LC_4_14_3 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_6_LC_4_14_3 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U400_SDRAM.MA_nesr_6_LC_4_14_3  (
            .in0(N__2966),
            .in1(N__6503),
            .in2(N__2957),
            .in3(N__6338),
            .lcout(MA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_6C_net ),
            .ce(N__6269),
            .sr(N__6169));
    defparam \U400_SDRAM.TACK_RNO_3_LC_5_4_0 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_3_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_3_LC_5_4_0 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \U400_SDRAM.TACK_RNO_3_LC_5_4_0  (
            .in0(N__2930),
            .in1(N__2920),
            .in2(_gnd_net_),
            .in3(N__4488),
            .lcout(\U400_SDRAM.un1_SDRAM_COUNTER52_4_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_EN_i_ess_RNO_0_LC_5_4_2 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_EN_i_ess_RNO_0_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_EN_i_ess_RNO_0_LC_5_4_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U400_SDRAM.TA_EN_i_ess_RNO_0_LC_5_4_2  (
            .in0(N__6187),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3197),
            .lcout(\U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_6_LC_5_4_3 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_6_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_6_LC_5_4_3 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \U400_SDRAM.TACK_RNO_6_LC_5_4_3  (
            .in0(N__4818),
            .in1(N__4900),
            .in2(N__4678),
            .in3(N__4609),
            .lcout(\U400_SDRAM.N_216 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.WRITE_CYCLE_RNI07LH_LC_5_4_7 .C_ON=1'b0;
    defparam \U400_SDRAM.WRITE_CYCLE_RNI07LH_LC_5_4_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.WRITE_CYCLE_RNI07LH_LC_5_4_7 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \U400_SDRAM.WRITE_CYCLE_RNI07LH_LC_5_4_7  (
            .in0(N__4659),
            .in1(N__4899),
            .in2(_gnd_net_),
            .in3(N__4608),
            .lcout(\U400_SDRAM.N_187 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_0_LC_5_5_0 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_0_LC_5_5_0 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_0_LC_5_5_0 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_0_LC_5_5_0  (
            .in0(N__3278),
            .in1(N__2909),
            .in2(N__2900),
            .in3(N__3499),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_0C_net ),
            .ce(N__3445),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_5_LC_5_5_1 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_5_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_5_LC_5_5_1 .LUT_INIT=16'b1111010110100010;
    LogicCell40 \U400_SDRAM.TACK_RNO_5_LC_5_5_1  (
            .in0(N__4908),
            .in1(N__4664),
            .in2(N__4619),
            .in3(N__4461),
            .lcout(\U400_SDRAM.TACK_7_iv_i_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_4_LC_5_5_2 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_4_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_4_LC_5_5_2 .LUT_INIT=16'b0110010101001110;
    LogicCell40 \U400_SDRAM.TACK_RNO_4_LC_5_5_2  (
            .in0(N__4820),
            .in1(N__4611),
            .in2(N__4679),
            .in3(N__4909),
            .lcout(),
            .ltout(\U400_SDRAM.TACK_7_iv_i_i_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_1_LC_5_5_3 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_1_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_1_LC_5_5_3 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U400_SDRAM.TACK_RNO_1_LC_5_5_3  (
            .in0(N__2891),
            .in1(N__3137),
            .in2(N__2885),
            .in3(N__4356),
            .lcout(\U400_SDRAM.N_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.WRITE_CYCLE_RNI18LH_LC_5_5_4 .C_ON=1'b0;
    defparam \U400_SDRAM.WRITE_CYCLE_RNI18LH_LC_5_5_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.WRITE_CYCLE_RNI18LH_LC_5_5_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U400_SDRAM.WRITE_CYCLE_RNI18LH_LC_5_5_4  (
            .in0(N__4663),
            .in1(N__4806),
            .in2(_gnd_net_),
            .in3(N__4610),
            .lcout(\U400_SDRAM.N_258 ),
            .ltout(\U400_SDRAM.N_258_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_0_LC_5_5_5 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_0_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_0_LC_5_5_5 .LUT_INIT=16'b1111111101110011;
    LogicCell40 \U400_SDRAM.TACK_RNO_0_LC_5_5_5  (
            .in0(N__4910),
            .in1(N__3131),
            .in2(N__3125),
            .in3(N__3122),
            .lcout(\U400_SDRAM.N_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNISAQQ4_1_LC_5_6_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNISAQQ4_1_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNISAQQ4_1_LC_5_6_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNISAQQ4_1_LC_5_6_1  (
            .in0(N__4795),
            .in1(N__5039),
            .in2(_gnd_net_),
            .in3(N__5395),
            .lcout(\U400_SDRAM.N_240 ),
            .ltout(\U400_SDRAM.N_240_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5_LC_5_6_2 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5_LC_5_6_2 .LUT_INIT=16'b1111111100111111;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5_LC_5_6_2  (
            .in0(_gnd_net_),
            .in1(N__3982),
            .in2(N__3110),
            .in3(N__5001),
            .lcout(\U400_SDRAM.N_219_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIMIPA1_1_LC_5_6_3 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIMIPA1_1_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIMIPA1_1_LC_5_6_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_RNIMIPA1_1_LC_5_6_3  (
            .in0(N__3107),
            .in1(N__3091),
            .in2(N__3080),
            .in3(N__3063),
            .lcout(\U400_SDRAM.un1_REFRESH_COUNTERlto7_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_1_LC_5_6_4 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_1_LC_5_6_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_1_LC_5_6_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_1_LC_5_6_4  (
            .in0(N__3064),
            .in1(_gnd_net_),
            .in2(N__3007),
            .in3(_gnd_net_),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_1C_net ),
            .ce(),
            .sr(N__2980));
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIUQPA1_5_LC_5_6_5 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIUQPA1_5_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIUQPA1_5_LC_5_6_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_RNIUQPA1_5_LC_5_6_5  (
            .in0(N__3049),
            .in1(N__3038),
            .in2(N__3023),
            .in3(N__2999),
            .lcout(\U400_SDRAM.un1_REFRESH_COUNTERlto7_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_0_LC_5_6_6 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_0_LC_5_6_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_0_LC_5_6_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_0_LC_5_6_6  (
            .in0(N__3000),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_1C_net ),
            .ce(),
            .sr(N__2980));
    defparam \U400_SDRAM.CS0_EN_RNO_0_LC_5_7_1 .C_ON=1'b0;
    defparam \U400_SDRAM.CS0_EN_RNO_0_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.CS0_EN_RNO_0_LC_5_7_1 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \U400_SDRAM.CS0_EN_RNO_0_LC_5_7_1  (
            .in0(N__3181),
            .in1(N__3259),
            .in2(N__3169),
            .in3(N__3550),
            .lcout(),
            .ltout(\U400_SDRAM.CS0_EN_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.CS0_EN_LC_5_7_2 .C_ON=1'b0;
    defparam \U400_SDRAM.CS0_EN_LC_5_7_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.CS0_EN_LC_5_7_2 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \U400_SDRAM.CS0_EN_LC_5_7_2  (
            .in0(N__4798),
            .in1(N__5045),
            .in2(N__3185),
            .in3(N__5397),
            .lcout(\U400_SDRAM.CS0_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS0_ENC_net ),
            .ce(),
            .sr(N__6160));
    defparam \U400_SDRAM.CS1_EN_RNO_0_LC_5_7_3 .C_ON=1'b0;
    defparam \U400_SDRAM.CS1_EN_RNO_0_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.CS1_EN_RNO_0_LC_5_7_3 .LUT_INIT=16'b0010001000101110;
    LogicCell40 \U400_SDRAM.CS1_EN_RNO_0_LC_5_7_3  (
            .in0(N__3631),
            .in1(N__3260),
            .in2(N__3170),
            .in3(N__3551),
            .lcout(),
            .ltout(\U400_SDRAM.CS1_EN_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.CS1_EN_LC_5_7_4 .C_ON=1'b0;
    defparam \U400_SDRAM.CS1_EN_LC_5_7_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.CS1_EN_LC_5_7_4 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \U400_SDRAM.CS1_EN_LC_5_7_4  (
            .in0(N__4799),
            .in1(N__5046),
            .in2(N__3149),
            .in3(N__5398),
            .lcout(\U400_SDRAM.CS1_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS0_ENC_net ),
            .ce(),
            .sr(N__6160));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_2_LC_5_7_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_2_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_2_LC_5_7_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_2_LC_5_7_5  (
            .in0(N__4441),
            .in1(N__4925),
            .in2(N__4597),
            .in3(N__4331),
            .lcout(\U400_SDRAM.N_114 ),
            .ltout(\U400_SDRAM.N_114_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNI5POA3_LC_5_7_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNI5POA3_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNI5POA3_LC_5_7_6 .LUT_INIT=16'b0100110000001000;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNI5POA3_LC_5_7_6  (
            .in0(N__5527),
            .in1(N__4789),
            .in2(N__3146),
            .in3(N__4380),
            .lcout(\U400_SDRAM.N_242 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIVG1P5_2_LC_5_7_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIVG1P5_2_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIVG1P5_2_LC_5_7_7 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIVG1P5_2_LC_5_7_7  (
            .in0(N__3143),
            .in1(N__3941),
            .in2(_gnd_net_),
            .in3(N__3258),
            .lcout(\U400_SDRAM.N_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI4ECU1_2_LC_5_8_0 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI4ECU1_2_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI4ECU1_2_LC_5_8_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI4ECU1_2_LC_5_8_0  (
            .in0(N__4333),
            .in1(N__4468),
            .in2(N__3530),
            .in3(N__5520),
            .lcout(\U400_SDRAM.N_220 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIRRB91_0_LC_5_8_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIRRB91_0_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIRRB91_0_LC_5_8_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIRRB91_0_LC_5_8_1  (
            .in0(N__4930),
            .in1(N__4589),
            .in2(_gnd_net_),
            .in3(N__4335),
            .lcout(\U400_SDRAM.N_261 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI7D8G1_0_LC_5_8_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI7D8G1_0_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI7D8G1_0_LC_5_8_3 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI7D8G1_0_LC_5_8_3  (
            .in0(N__4931),
            .in1(N__4588),
            .in2(N__4813),
            .in3(N__4332),
            .lcout(\U400_SDRAM.N_140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_1_LC_5_8_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_1_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_1_LC_5_8_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_0_1_LC_5_8_4  (
            .in0(N__4590),
            .in1(N__3421),
            .in2(_gnd_net_),
            .in3(N__5047),
            .lcout(\U400_SDRAM.N_207 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNI5POA3_0_LC_5_8_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNI5POA3_0_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNI5POA3_0_LC_5_8_5 .LUT_INIT=16'b0011101100110001;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNI5POA3_0_LC_5_8_5  (
            .in0(N__4785),
            .in1(N__5391),
            .in2(N__5546),
            .in3(N__4381),
            .lcout(\U400_SDRAM.SDRAM_CONFIGURED_RNI5POA3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI36NC1_2_LC_5_8_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI36NC1_2_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI36NC1_2_LC_5_8_6 .LUT_INIT=16'b0000000011101111;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI36NC1_2_LC_5_8_6  (
            .in0(N__4334),
            .in1(N__4469),
            .in2(N__4949),
            .in3(N__5521),
            .lcout(),
            .ltout(\U400_SDRAM.N_230_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI2LE84_2_LC_5_8_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI2LE84_2_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI2LE84_2_LC_5_8_7 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI2LE84_2_LC_5_8_7  (
            .in0(N__3952),
            .in1(N__3661),
            .in2(N__3248),
            .in3(N__3419),
            .lcout(\U400_SDRAM.N_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_9_LC_5_12_6 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_9_LC_5_12_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_9_LC_5_12_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U400_SDRAM.MA_nesr_9_LC_5_12_6  (
            .in0(N__6502),
            .in1(N__6068),
            .in2(N__3245),
            .in3(N__5968),
            .lcout(MA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_9C_net ),
            .ce(N__6267),
            .sr(N__6164));
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_0_o2_1_LC_6_1_0 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_0_o2_1_LC_6_1_0 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_0_o2_1_LC_6_1_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_0_o2_1_LC_6_1_0  (
            .in0(N__3218),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3212),
            .lcout(U400_ADDRESS_DECODE_RAM_SPACE_i_o3_0_o2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.BURST_RNISKH51_LC_6_4_0 .C_ON=1'b0;
    defparam \U400_SDRAM.BURST_RNISKH51_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.BURST_RNISKH51_LC_6_4_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U400_SDRAM.BURST_RNISKH51_LC_6_4_0  (
            .in0(N__4217),
            .in1(N__4106),
            .in2(N__4256),
            .in3(N__3738),
            .lcout(\U400_SDRAM.TA_COUNTER_0_sqmuxa ),
            .ltout(\U400_SDRAM.TA_COUNTER_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_EN_i_ess_RNO_1_LC_6_4_1 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_EN_i_ess_RNO_1_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_EN_i_ess_RNO_1_LC_6_4_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \U400_SDRAM.TA_EN_i_ess_RNO_1_LC_6_4_1  (
            .in0(N__4171),
            .in1(N__3706),
            .in2(N__3200),
            .in3(N__4146),
            .lcout(\U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_EN_i_ess_LC_6_4_4 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_EN_i_ess_LC_6_4_4 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.TA_EN_i_ess_LC_6_4_4 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U400_SDRAM.TA_EN_i_ess_LC_6_4_4  (
            .in0(N__4147),
            .in1(N__3983),
            .in2(_gnd_net_),
            .in3(N__4172),
            .lcout(TA_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4070),
            .ce(N__3191),
            .sr(N__6171));
    defparam \U400_SDRAM.BANK0_LC_6_5_0 .C_ON=1'b0;
    defparam \U400_SDRAM.BANK0_LC_6_5_0 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.BANK0_LC_6_5_0 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \U400_SDRAM.BANK0_LC_6_5_0  (
            .in0(N__3367),
            .in1(N__3340),
            .in2(N__3398),
            .in3(N__5002),
            .lcout(BANK0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.BANK0C_net ),
            .ce(),
            .sr(N__6165));
    defparam \U400_SDRAM.BANK1_LC_6_5_1 .C_ON=1'b0;
    defparam \U400_SDRAM.BANK1_LC_6_5_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.BANK1_LC_6_5_1 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U400_SDRAM.BANK1_LC_6_5_1  (
            .in0(N__5003),
            .in1(N__3316),
            .in2(N__3356),
            .in3(N__3341),
            .lcout(BANK1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.BANK0C_net ),
            .ce(),
            .sr(N__6165));
    defparam \U400_SDRAM.RAM_CYCLE_LC_6_5_2 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_LC_6_5_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.RAM_CYCLE_LC_6_5_2 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_LC_6_5_2  (
            .in0(N__3272),
            .in1(N__3572),
            .in2(N__3981),
            .in3(N__5150),
            .lcout(\U400_SDRAM.RAM_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.BANK0C_net ),
            .ce(),
            .sr(N__6165));
    defparam \U400_SDRAM.WRITE_CYCLE_LC_6_5_3 .C_ON=1'b0;
    defparam \U400_SDRAM.WRITE_CYCLE_LC_6_5_3 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.WRITE_CYCLE_LC_6_5_3 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \U400_SDRAM.WRITE_CYCLE_LC_6_5_3  (
            .in0(N__3570),
            .in1(N__3305),
            .in2(_gnd_net_),
            .in3(N__4671),
            .lcout(\U400_SDRAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.BANK0C_net ),
            .ce(),
            .sr(N__6165));
    defparam \U400_SDRAM.TACK_LC_6_5_5 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_LC_6_5_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TACK_LC_6_5_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \U400_SDRAM.TACK_LC_6_5_5  (
            .in0(N__3293),
            .in1(N__3287),
            .in2(_gnd_net_),
            .in3(N__4151),
            .lcout(\U400_SDRAM.TACKZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.BANK0C_net ),
            .ce(),
            .sr(N__6165));
    defparam \U400_SDRAM.BURST_LC_6_5_6 .C_ON=1'b0;
    defparam \U400_SDRAM.BURST_LC_6_5_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.BURST_LC_6_5_6 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \U400_SDRAM.BURST_LC_6_5_6  (
            .in0(N__5757),
            .in1(N__3571),
            .in2(N__3743),
            .in3(N__5824),
            .lcout(\U400_SDRAM.BURSTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.BANK0C_net ),
            .ce(),
            .sr(N__6165));
    defparam \U400_SDRAM.BURST8_i_0_i_i_o2_LC_6_6_0 .C_ON=1'b0;
    defparam \U400_SDRAM.BURST8_i_0_i_i_o2_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.BURST8_i_0_i_i_o2_LC_6_6_0 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U400_SDRAM.BURST8_i_0_i_i_o2_LC_6_6_0  (
            .in0(N__5756),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5823),
            .lcout(\U400_SDRAM.N_118 ),
            .ltout(\U400_SDRAM.N_118_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_0_LC_6_6_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_0_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_0_LC_6_6_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_0_0_LC_6_6_1  (
            .in0(N__5394),
            .in1(N__5043),
            .in2(N__3281),
            .in3(N__4998),
            .lcout(\U400_SDRAM.N_215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_LC_6_6_2 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_LC_6_6_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.RAM_CYCLE_START_LC_6_6_2 .LUT_INIT=16'b1100000011100000;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_LC_6_6_2  (
            .in0(N__4999),
            .in1(N__5054),
            .in2(N__3966),
            .in3(N__3271),
            .lcout(\U400_SDRAM.RAM_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4067),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_RNO_3_LC_6_6_3 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_3_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_3_LC_6_6_3 .LUT_INIT=16'b1101110110101010;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_RNO_3_LC_6_6_3  (
            .in0(N__4774),
            .in1(N__4587),
            .in2(_gnd_net_),
            .in3(N__4901),
            .lcout(\U400_SDRAM.N_189 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_RNI8BL33_8_LC_6_6_4 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNI8BL33_8_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNI8BL33_8_LC_6_6_4 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_RNI8BL33_8_LC_6_6_4  (
            .in0(N__3799),
            .in1(N__3829),
            .in2(N__5544),
            .in3(N__3814),
            .lcout(\U400_SDRAM.N_236 ),
            .ltout(\U400_SDRAM.N_236_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_RNI58I35_LC_6_6_5 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNI58I35_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNI58I35_LC_6_6_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_RNI58I35_LC_6_6_5  (
            .in0(N__5393),
            .in1(N__4794),
            .in2(N__3575),
            .in3(N__4996),
            .lcout(\U400_SDRAM.N_23_i ),
            .ltout(\U400_SDRAM.N_23_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5_0_LC_6_6_6 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5_0_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5_0_LC_6_6_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5_0_LC_6_6_6  (
            .in0(N__3940),
            .in1(_gnd_net_),
            .in2(N__3560),
            .in3(_gnd_net_),
            .lcout(\U400_SDRAM.N_259 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIUFE78_LC_6_6_7 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIUFE78_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIUFE78_LC_6_6_7 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_RNIUFE78_LC_6_6_7  (
            .in0(N__5392),
            .in1(N__3557),
            .in2(N__5048),
            .in3(N__4997),
            .lcout(\U400_SDRAM.N_139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_1_LC_6_7_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_1_LC_6_7_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_1_LC_6_7_1 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_1_LC_6_7_1  (
            .in0(N__3542),
            .in1(N__3492),
            .in2(N__3512),
            .in3(N__3520),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_1C_net ),
            .ce(N__3446),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.WRITE_CYCLE_RNICOHO_LC_6_7_2 .C_ON=1'b0;
    defparam \U400_SDRAM.WRITE_CYCLE_RNICOHO_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.WRITE_CYCLE_RNICOHO_LC_6_7_2 .LUT_INIT=16'b0111011001100110;
    LogicCell40 \U400_SDRAM.WRITE_CYCLE_RNICOHO_LC_6_7_2  (
            .in0(N__4773),
            .in1(N__4574),
            .in2(N__4687),
            .in3(N__4940),
            .lcout(\U400_SDRAM.N_198 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_3_LC_6_7_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_3_LC_6_7_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_3_LC_6_7_4 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_3_LC_6_7_4  (
            .in0(N__3521),
            .in1(N__3511),
            .in2(N__3500),
            .in3(N__3458),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_1C_net ),
            .ce(N__3446),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_1_LC_6_8_0 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_1_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_1_LC_6_8_0 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_1_1_LC_6_8_0  (
            .in0(N__3428),
            .in1(N__4826),
            .in2(N__3677),
            .in3(N__3641),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_1_LC_6_8_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_1_LC_6_8_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_CMD_1_LC_6_8_1 .LUT_INIT=16'b1111110010101010;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_1_LC_6_8_1  (
            .in0(N__6040),
            .in1(N__3689),
            .in2(N__3680),
            .in3(N__5349),
            .lcout(\U400_SDRAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_CMD_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_1_LC_6_8_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_1_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_1_LC_6_8_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_2_1_LC_6_8_2  (
            .in0(N__5549),
            .in1(N__4592),
            .in2(_gnd_net_),
            .in3(N__4946),
            .lcout(\U400_SDRAM.N_250 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_2_LC_6_8_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_2_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_2_LC_6_8_3 .LUT_INIT=16'b0011100111101010;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_2_2_LC_6_8_3  (
            .in0(N__4947),
            .in1(N__5550),
            .in2(N__4615),
            .in3(N__4492),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_cnst_0_31_i_i_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_2_LC_6_8_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_2_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_2_LC_6_8_4 .LUT_INIT=16'b1111001111111011;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_1_2_LC_6_8_4  (
            .in0(N__3650),
            .in1(N__3932),
            .in2(N__3668),
            .in3(N__5552),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_cnst_0_31_i_i_i_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_2_LC_6_8_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_2_LC_6_8_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_CMD_2_LC_6_8_5 .LUT_INIT=16'b1110111011100010;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_2_LC_6_8_5  (
            .in0(N__6425),
            .in1(N__5350),
            .in2(N__3665),
            .in3(N__4961),
            .lcout(\U400_SDRAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_CMD_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_ne_RNO_0_0_LC_6_8_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_ne_RNO_0_0_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_ne_RNO_0_0_LC_6_8_6 .LUT_INIT=16'b0010101011111111;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_ne_RNO_0_0_LC_6_8_6  (
            .in0(N__3662),
            .in1(N__4796),
            .in2(N__4688),
            .in3(N__3936),
            .lcout(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_4_1_LC_6_8_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_4_1_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_4_1_LC_6_8_7 .LUT_INIT=16'b1111111101001111;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_4_1_LC_6_8_7  (
            .in0(N__5551),
            .in1(N__3649),
            .in2(N__3965),
            .in3(N__4393),
            .lcout(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.CS1n_LC_6_9_2 .C_ON=1'b0;
    defparam \U400_SDRAM.CS1n_LC_6_9_2 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.CS1n_LC_6_9_2 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \U400_SDRAM.CS1n_LC_6_9_2  (
            .in0(N__6426),
            .in1(N__6031),
            .in2(N__3635),
            .in3(N__5924),
            .lcout(CS1n_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS1nC_net ),
            .ce(),
            .sr(N__6161));
    defparam \U400_SDRAM.MA_nesr_12_LC_6_12_2 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_12_LC_6_12_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_12_LC_6_12_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U400_SDRAM.MA_nesr_12_LC_6_12_2  (
            .in0(N__6462),
            .in1(N__6074),
            .in2(N__3605),
            .in3(N__5960),
            .lcout(MA_c_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_12C_net ),
            .ce(N__6258),
            .sr(N__6170));
    defparam \U400_SDRAM.TA_OUT_LC_7_3_3 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_OUT_LC_7_3_3 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.TA_OUT_LC_7_3_3 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \U400_SDRAM.TA_OUT_LC_7_3_3  (
            .in0(N__4288),
            .in1(N__3713),
            .in2(N__3769),
            .in3(N__3722),
            .lcout(TA_OUT),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4074),
            .ce(),
            .sr(N__6173));
    defparam \U400_SDRAM.TA_COUNTER_RNIAJGG1_3_LC_7_4_1 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_RNIAJGG1_3_LC_7_4_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_COUNTER_RNIAJGG1_3_LC_7_4_1 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_RNIAJGG1_3_LC_7_4_1  (
            .in0(N__4279),
            .in1(N__4213),
            .in2(N__4255),
            .in3(N__4102),
            .lcout(\U400_SDRAM.TA_COUNTER27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_BYTE_ENABLE.un1_UUBEn_i_0_0_LC_7_4_2 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un1_UUBEn_i_0_0_LC_7_4_2 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un1_UUBEn_i_0_0_LC_7_4_2 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \U400_BYTE_ENABLE.un1_UUBEn_i_0_0_LC_7_4_2  (
            .in0(N__5857),
            .in1(N__5246),
            .in2(N__5195),
            .in3(N__5267),
            .lcout(N_66),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_RNIAJGG1_0_3_LC_7_4_3 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_RNIAJGG1_0_3_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_COUNTER_RNIAJGG1_0_3_LC_7_4_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U400_SDRAM.TA_COUNTER_RNIAJGG1_0_3_LC_7_4_3  (
            .in0(N__4278),
            .in1(N__4212),
            .in2(N__4254),
            .in3(N__4103),
            .lcout(\U400_SDRAM.TA_COUNTER23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_OUT_RNO_0_LC_7_4_4 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_OUT_RNO_0_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_OUT_RNO_0_LC_7_4_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U400_SDRAM.TA_OUT_RNO_0_LC_7_4_4  (
            .in0(N__4105),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3739),
            .lcout(\U400_SDRAM.TA_EN11_m ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_OUT_RNO_2_LC_7_4_6 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_OUT_RNO_2_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_OUT_RNO_2_LC_7_4_6 .LUT_INIT=16'b1110111011111100;
    LogicCell40 \U400_SDRAM.TA_OUT_RNO_2_LC_7_4_6  (
            .in0(N__4104),
            .in1(N__4249),
            .in2(N__4222),
            .in3(N__4280),
            .lcout(),
            .ltout(\U400_SDRAM.un1_TA_COUNTER26_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_OUT_RNO_1_LC_7_4_7 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_OUT_RNO_1_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_OUT_RNO_1_LC_7_4_7 .LUT_INIT=16'b0000111100000011;
    LogicCell40 \U400_SDRAM.TA_OUT_RNO_1_LC_7_4_7  (
            .in0(_gnd_net_),
            .in1(N__4177),
            .in2(N__3716),
            .in3(N__4148),
            .lcout(\U400_SDRAM.un1_TA_COUNTER26_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_1_LC_7_5_0 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_1_LC_7_5_0 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_1_LC_7_5_0 .LUT_INIT=16'b0100100000000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_1_LC_7_5_0  (
            .in0(N__4109),
            .in1(N__3968),
            .in2(N__4223),
            .in3(N__3695),
            .lcout(\U400_SDRAM.TA_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4071),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNI0LUG4_LC_7_5_1 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNI0LUG4_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNI0LUG4_LC_7_5_1 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \U400_SDRAM.TACK_RNI0LUG4_LC_7_5_1  (
            .in0(N__4149),
            .in1(N__3707),
            .in2(N__4178),
            .in3(N__4117),
            .lcout(\U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0 ),
            .ltout(\U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_2_LC_7_5_2 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_2_LC_7_5_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_2_LC_7_5_2 .LUT_INIT=16'b0110000000000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_2_LC_7_5_2  (
            .in0(N__4284),
            .in1(N__4189),
            .in2(N__4292),
            .in3(N__3969),
            .lcout(\U400_SDRAM.TA_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4071),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_3_LC_7_5_4 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_3_LC_7_5_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_3_LC_7_5_4 .LUT_INIT=16'b0100110010000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_3_LC_7_5_4  (
            .in0(N__4190),
            .in1(N__3970),
            .in2(N__4289),
            .in3(N__4253),
            .lcout(\U400_SDRAM.TA_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4071),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_RNIJ78O_1_LC_7_5_5 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_RNIJ78O_1_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_COUNTER_RNIJ78O_1_LC_7_5_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_RNIJ78O_1_LC_7_5_5  (
            .in0(_gnd_net_),
            .in1(N__4218),
            .in2(_gnd_net_),
            .in3(N__4107),
            .lcout(\U400_SDRAM.CO1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_RNO_0_0_LC_7_5_6 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_RNO_0_0_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_COUNTER_RNO_0_0_LC_7_5_6 .LUT_INIT=16'b0010001001100110;
    LogicCell40 \U400_SDRAM.TA_COUNTER_RNO_0_0_LC_7_5_6  (
            .in0(N__4108),
            .in1(N__4173),
            .in2(_gnd_net_),
            .in3(N__4150),
            .lcout(),
            .ltout(\U400_SDRAM.TA_COUNTER_7_f1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_0_LC_7_5_7 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_0_LC_7_5_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_0_LC_7_5_7 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \U400_SDRAM.TA_COUNTER_0_LC_7_5_7  (
            .in0(N__3967),
            .in1(_gnd_net_),
            .in2(N__4121),
            .in3(N__4118),
            .lcout(\U400_SDRAM.TA_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4071),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_RNO_2_LC_7_6_0 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_2_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_2_LC_7_6_0 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_RNO_2_LC_7_6_0  (
            .in0(N__3989),
            .in1(N__4473),
            .in2(N__5545),
            .in3(N__4357),
            .lcout(\U400_SDRAM.un1_SDRAM_COUNTER52_2_0_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_0_o2dup_LC_7_6_1 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_0_o2dup_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_0_o2dup_LC_7_6_1 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_0_o2dup_LC_7_6_1  (
            .in0(N__5083),
            .in1(N__5120),
            .in2(N__5144),
            .in3(N__3942),
            .lcout(RAM_SPACE_i_o3_0_o2dup),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_RNO_1_LC_7_6_6 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_1_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_1_LC_7_6_6 .LUT_INIT=16'b1111100011111111;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_RNO_1_LC_7_6_6  (
            .in0(N__3833),
            .in1(N__3818),
            .in2(N__3803),
            .in3(N__4995),
            .lcout(),
            .ltout(\U400_SDRAM.N_195_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_RNO_0_LC_7_6_7 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_0_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_0_LC_7_6_7 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_RNO_0_LC_7_6_7  (
            .in0(N__5159),
            .in1(N__4596),
            .in2(N__5153),
            .in3(N__4948),
            .lcout(\U400_SDRAM.N_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_RNO_0_LC_7_7_3 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNO_0_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNO_0_LC_7_7_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_RNO_0_LC_7_7_3  (
            .in0(N__5143),
            .in1(N__5116),
            .in2(N__5090),
            .in3(N__5063),
            .lcout(\U400_SDRAM.N_225 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_2_LC_7_7_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_2_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_2_LC_7_7_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_0_2_LC_7_7_4  (
            .in0(N__4491),
            .in1(N__5044),
            .in2(_gnd_net_),
            .in3(N__5000),
            .lcout(\U400_SDRAM.N_228 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_6_1_LC_7_7_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_6_1_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_6_1_LC_7_7_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_6_1_LC_7_7_5  (
            .in0(N__4790),
            .in1(N__4572),
            .in2(_gnd_net_),
            .in3(N__4941),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_a2_2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_5_1_LC_7_7_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_5_1_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_5_1_LC_7_7_6 .LUT_INIT=16'b0011001000110000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_5_1_LC_7_7_6  (
            .in0(N__4573),
            .in1(N__5528),
            .in2(N__4955),
            .in3(N__4489),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_3_1_LC_7_7_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_3_1_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_3_1_LC_7_7_7 .LUT_INIT=16'b1111000111111010;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_3_1_LC_7_7_7  (
            .in0(N__4490),
            .in1(N__5529),
            .in2(N__4952),
            .in3(N__4942),
            .lcout(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_ne_RNO_2_0_LC_7_8_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_ne_RNO_2_0_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_ne_RNO_2_0_LC_7_8_4 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_ne_RNO_2_0_LC_7_8_4  (
            .in0(N__4797),
            .in1(N__4680),
            .in2(N__5548),
            .in3(N__4591),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_a2_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_ne_RNO_1_0_LC_7_8_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_ne_RNO_1_0_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_ne_RNO_1_0_LC_7_8_5 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_ne_RNO_1_0_LC_7_8_5  (
            .in0(N__4493),
            .in1(N__4394),
            .in2(N__4364),
            .in3(N__4361),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_ne_0_LC_7_8_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_ne_0_LC_7_8_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_CMD_ne_0_LC_7_8_6 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_ne_0_LC_7_8_6  (
            .in0(N__5533),
            .in1(N__5414),
            .in2(N__5408),
            .in3(N__5405),
            .lcout(\U400_SDRAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_CMD_ne_0C_net ),
            .ce(N__5354),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_11_LC_7_12_5 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_11_LC_7_12_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_11_LC_7_12_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U400_SDRAM.MA_nesr_11_LC_7_12_5  (
            .in0(N__6485),
            .in1(N__6075),
            .in2(N__5336),
            .in3(N__5959),
            .lcout(MA_c_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_11C_net ),
            .ce(N__6254),
            .sr(N__6172));
    defparam \U400_SDRAM.MA_nesr_RNO_0_5_LC_7_14_7 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_RNO_0_5_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.MA_nesr_RNO_0_5_LC_7_14_7 .LUT_INIT=16'b0101111101001110;
    LogicCell40 \U400_SDRAM.MA_nesr_RNO_0_5_LC_7_14_7  (
            .in0(N__6499),
            .in1(N__6070),
            .in2(N__5312),
            .in3(N__5958),
            .lcout(\U400_SDRAM.MA_5_iv_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_5_LC_7_15_7 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_5_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_5_LC_7_15_7 .LUT_INIT=16'b1011101100110011;
    LogicCell40 \U400_SDRAM.MA_nesr_5_LC_7_15_7  (
            .in0(N__5300),
            .in1(N__5288),
            .in2(_gnd_net_),
            .in3(N__6337),
            .lcout(MA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_5C_net ),
            .ce(N__6265),
            .sr(N__6178));
    defparam \U400_BYTE_ENABLE.un1_UUBEn_i_0_0_x2_LC_8_4_4 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un1_UUBEn_i_0_0_x2_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un1_UUBEn_i_0_0_x2_LC_8_4_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U400_BYTE_ENABLE.un1_UUBEn_i_0_0_x2_LC_8_4_4  (
            .in0(_gnd_net_),
            .in1(N__5822),
            .in2(_gnd_net_),
            .in3(N__5755),
            .lcout(\U400_BYTE_ENABLE.N_101_i ),
            .ltout(\U400_BYTE_ENABLE.N_101_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_BYTE_ENABLE.un1_LMBEn_i_0_0_LC_8_4_5 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un1_LMBEn_i_0_0_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un1_LMBEn_i_0_0_LC_8_4_5 .LUT_INIT=16'b1111111111010000;
    LogicCell40 \U400_BYTE_ENABLE.un1_LMBEn_i_0_0_LC_8_4_5  (
            .in0(N__5853),
            .in1(N__5245),
            .in2(N__5261),
            .in3(N__5193),
            .lcout(un1_LMBEn_i_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_BYTE_ENABLE.un1_UMBEn_i_0_0_o2_LC_8_5_0 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un1_UMBEn_i_0_0_o2_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un1_UMBEn_i_0_0_o2_LC_8_5_0 .LUT_INIT=16'b1111111100000010;
    LogicCell40 \U400_BYTE_ENABLE.un1_UMBEn_i_0_0_o2_LC_8_5_0  (
            .in0(N__5759),
            .in1(N__5238),
            .in2(N__5825),
            .in3(N__5183),
            .lcout(\U400_BYTE_ENABLE.N_168 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_ne_RNIIMNC_0_LC_8_12_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_ne_RNIIMNC_0_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_ne_RNIIMNC_0_LC_8_12_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_ne_RNIIMNC_0_LC_8_12_1  (
            .in0(N__6474),
            .in1(N__6062),
            .in2(_gnd_net_),
            .in3(N__5954),
            .lcout(\U400_SDRAM.MA19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_ne_RNI80KS_0_LC_8_12_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_ne_RNI80KS_0_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_ne_RNI80KS_0_LC_8_12_3 .LUT_INIT=16'b1111011011110111;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_ne_RNI80KS_0_LC_8_12_3  (
            .in0(N__6475),
            .in1(N__6063),
            .in2(N__6191),
            .in3(N__5955),
            .lcout(\U400_SDRAM.un1_MA20_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_10_LC_8_13_3 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_10_LC_8_13_3 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_10_LC_8_13_3 .LUT_INIT=16'b0100000001000100;
    LogicCell40 \U400_SDRAM.MA_nesr_10_LC_8_13_3  (
            .in0(N__6501),
            .in1(N__6076),
            .in2(N__6110),
            .in3(N__5956),
            .lcout(MA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_10C_net ),
            .ce(N__6237),
            .sr(N__6177));
    defparam \U400_SDRAM.MA_nesr_RNO_0_1_LC_8_14_7 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_RNO_0_1_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.MA_nesr_RNO_0_1_LC_8_14_7 .LUT_INIT=16'b0101111101001110;
    LogicCell40 \U400_SDRAM.MA_nesr_RNO_0_1_LC_8_14_7  (
            .in0(N__6500),
            .in1(N__6077),
            .in2(N__5984),
            .in3(N__5957),
            .lcout(\U400_SDRAM.MA_5_iv_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_BYTE_ENABLE.un1_UMBEn_i_0_0_LC_9_4_0 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un1_UMBEn_i_0_0_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un1_UMBEn_i_0_0_LC_9_4_0 .LUT_INIT=16'b1111111101001000;
    LogicCell40 \U400_BYTE_ENABLE.un1_UMBEn_i_0_0_LC_9_4_0  (
            .in0(N__5812),
            .in1(N__5867),
            .in2(N__5758),
            .in3(N__5770),
            .lcout(N_63),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_BYTE_ENABLE.un1_LLBEn_i_0_0_LC_9_4_7 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un1_LLBEn_i_0_0_LC_9_4_7 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un1_LLBEn_i_0_0_LC_9_4_7 .LUT_INIT=16'b1111000111110100;
    LogicCell40 \U400_BYTE_ENABLE.un1_LLBEn_i_0_0_LC_9_4_7  (
            .in0(N__5866),
            .in1(N__5811),
            .in2(N__5771),
            .in3(N__5748),
            .lcout(un1_LLBEn_i_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TAn_obuft_RNO_LC_9_6_1.C_ON=1'b0;
    defparam TAn_obuft_RNO_LC_9_6_1.SEQ_MODE=4'b0000;
    defparam TAn_obuft_RNO_LC_9_6_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 TAn_obuft_RNO_LC_9_6_1 (
            .in0(N__5684),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_526_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_3_LC_9_13_7 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_3_LC_9_13_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_3_LC_9_13_7 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U400_SDRAM.MA_nesr_3_LC_9_13_7  (
            .in0(N__5663),
            .in1(N__6495),
            .in2(N__5654),
            .in3(N__6310),
            .lcout(MA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_3C_net ),
            .ce(N__6241),
            .sr(N__6179));
    defparam \U400_SDRAM.MA_nesr_2_LC_9_15_0 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_2_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_2_LC_9_15_0 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \U400_SDRAM.MA_nesr_2_LC_9_15_0  (
            .in0(N__6335),
            .in1(N__5621),
            .in2(N__5609),
            .in3(N__6497),
            .lcout(MA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_2C_net ),
            .ce(N__6266),
            .sr(N__6180));
    defparam \U400_SDRAM.MA_nesr_0_LC_9_15_3 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_0_LC_9_15_3 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_0_LC_9_15_3 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U400_SDRAM.MA_nesr_0_LC_9_15_3  (
            .in0(N__5588),
            .in1(N__6496),
            .in2(N__5576),
            .in3(N__6334),
            .lcout(MA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_2C_net ),
            .ce(N__6266),
            .sr(N__6180));
    defparam \U400_SDRAM.MA_nesr_4_LC_9_15_4 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_4_LC_9_15_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_4_LC_9_15_4 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \U400_SDRAM.MA_nesr_4_LC_9_15_4  (
            .in0(N__6336),
            .in1(N__6530),
            .in2(N__6518),
            .in3(N__6498),
            .lcout(MA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_2C_net ),
            .ce(N__6266),
            .sr(N__6180));
    defparam \U400_SDRAM.MA_nesr_1_LC_9_15_5 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_1_LC_9_15_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_1_LC_9_15_5 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \U400_SDRAM.MA_nesr_1_LC_9_15_5  (
            .in0(N__6353),
            .in1(N__6347),
            .in2(_gnd_net_),
            .in3(N__6333),
            .lcout(MA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_2C_net ),
            .ce(N__6266),
            .sr(N__6180));
endmodule // U400_TOP

module U110_BUFFERS (

    output IDELENn, IDEHRENn, IDEHWENn, IDELATCH

);

//ATA BUFFERS

assign IDELENn = 1;
assign IDEHRENn = 1;
assign IDEHWENn = 1;
assign IDELATCH = 0;


endmodule

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 16 2025 18:12:46

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    CMA,
    SIZ,
    DRA,
    A,
    RAMENn,
    TSn,
    LMBEn,
    DMA_LATCH_EN,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    UUBEn,
    LDSn,
    LATCH_CLK,
    CASUn,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    UMBEn,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    RAMSPACEn,
    WEn,
    REGENn,
    LLBEn,
    DBRn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    output [10:0] CMA;
    input [1:0] SIZ;
    input [9:0] DRA;
    input [20:0] A;
    output RAMENn;
    input TSn;
    output LMBEn;
    output DMA_LATCH_EN;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output UUBEn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    output UMBEn;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    output LLBEn;
    input DBRn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__11850;
    wire N__11849;
    wire N__11848;
    wire N__11841;
    wire N__11840;
    wire N__11839;
    wire N__11832;
    wire N__11831;
    wire N__11830;
    wire N__11823;
    wire N__11822;
    wire N__11821;
    wire N__11814;
    wire N__11813;
    wire N__11812;
    wire N__11805;
    wire N__11804;
    wire N__11803;
    wire N__11796;
    wire N__11795;
    wire N__11794;
    wire N__11787;
    wire N__11786;
    wire N__11785;
    wire N__11778;
    wire N__11777;
    wire N__11776;
    wire N__11769;
    wire N__11768;
    wire N__11767;
    wire N__11760;
    wire N__11759;
    wire N__11758;
    wire N__11751;
    wire N__11750;
    wire N__11749;
    wire N__11742;
    wire N__11741;
    wire N__11740;
    wire N__11733;
    wire N__11732;
    wire N__11731;
    wire N__11724;
    wire N__11723;
    wire N__11722;
    wire N__11715;
    wire N__11714;
    wire N__11713;
    wire N__11706;
    wire N__11705;
    wire N__11704;
    wire N__11697;
    wire N__11696;
    wire N__11695;
    wire N__11688;
    wire N__11687;
    wire N__11686;
    wire N__11679;
    wire N__11678;
    wire N__11677;
    wire N__11670;
    wire N__11669;
    wire N__11668;
    wire N__11661;
    wire N__11660;
    wire N__11659;
    wire N__11652;
    wire N__11651;
    wire N__11650;
    wire N__11643;
    wire N__11642;
    wire N__11641;
    wire N__11634;
    wire N__11633;
    wire N__11632;
    wire N__11625;
    wire N__11624;
    wire N__11623;
    wire N__11616;
    wire N__11615;
    wire N__11614;
    wire N__11607;
    wire N__11606;
    wire N__11605;
    wire N__11598;
    wire N__11597;
    wire N__11596;
    wire N__11589;
    wire N__11588;
    wire N__11587;
    wire N__11580;
    wire N__11579;
    wire N__11578;
    wire N__11571;
    wire N__11570;
    wire N__11569;
    wire N__11562;
    wire N__11561;
    wire N__11560;
    wire N__11553;
    wire N__11552;
    wire N__11551;
    wire N__11544;
    wire N__11543;
    wire N__11542;
    wire N__11535;
    wire N__11534;
    wire N__11533;
    wire N__11526;
    wire N__11525;
    wire N__11524;
    wire N__11517;
    wire N__11516;
    wire N__11515;
    wire N__11508;
    wire N__11507;
    wire N__11506;
    wire N__11499;
    wire N__11498;
    wire N__11497;
    wire N__11490;
    wire N__11489;
    wire N__11488;
    wire N__11481;
    wire N__11480;
    wire N__11479;
    wire N__11472;
    wire N__11471;
    wire N__11470;
    wire N__11463;
    wire N__11462;
    wire N__11461;
    wire N__11454;
    wire N__11453;
    wire N__11452;
    wire N__11445;
    wire N__11444;
    wire N__11443;
    wire N__11436;
    wire N__11435;
    wire N__11434;
    wire N__11427;
    wire N__11426;
    wire N__11425;
    wire N__11418;
    wire N__11417;
    wire N__11416;
    wire N__11409;
    wire N__11408;
    wire N__11407;
    wire N__11400;
    wire N__11399;
    wire N__11398;
    wire N__11391;
    wire N__11390;
    wire N__11389;
    wire N__11382;
    wire N__11381;
    wire N__11380;
    wire N__11373;
    wire N__11372;
    wire N__11371;
    wire N__11364;
    wire N__11363;
    wire N__11362;
    wire N__11355;
    wire N__11354;
    wire N__11353;
    wire N__11346;
    wire N__11345;
    wire N__11344;
    wire N__11337;
    wire N__11336;
    wire N__11335;
    wire N__11328;
    wire N__11327;
    wire N__11326;
    wire N__11319;
    wire N__11318;
    wire N__11317;
    wire N__11310;
    wire N__11309;
    wire N__11308;
    wire N__11301;
    wire N__11300;
    wire N__11299;
    wire N__11292;
    wire N__11291;
    wire N__11290;
    wire N__11283;
    wire N__11282;
    wire N__11281;
    wire N__11274;
    wire N__11273;
    wire N__11272;
    wire N__11265;
    wire N__11264;
    wire N__11263;
    wire N__11256;
    wire N__11255;
    wire N__11254;
    wire N__11247;
    wire N__11246;
    wire N__11245;
    wire N__11238;
    wire N__11237;
    wire N__11236;
    wire N__11229;
    wire N__11228;
    wire N__11227;
    wire N__11220;
    wire N__11219;
    wire N__11218;
    wire N__11211;
    wire N__11210;
    wire N__11209;
    wire N__11202;
    wire N__11201;
    wire N__11200;
    wire N__11193;
    wire N__11192;
    wire N__11191;
    wire N__11184;
    wire N__11183;
    wire N__11182;
    wire N__11175;
    wire N__11174;
    wire N__11173;
    wire N__11166;
    wire N__11165;
    wire N__11164;
    wire N__11157;
    wire N__11156;
    wire N__11155;
    wire N__11148;
    wire N__11147;
    wire N__11146;
    wire N__11139;
    wire N__11138;
    wire N__11137;
    wire N__11130;
    wire N__11129;
    wire N__11128;
    wire N__11121;
    wire N__11120;
    wire N__11119;
    wire N__11112;
    wire N__11111;
    wire N__11110;
    wire N__11103;
    wire N__11102;
    wire N__11101;
    wire N__11094;
    wire N__11093;
    wire N__11092;
    wire N__11085;
    wire N__11084;
    wire N__11083;
    wire N__11076;
    wire N__11075;
    wire N__11074;
    wire N__11067;
    wire N__11066;
    wire N__11065;
    wire N__11058;
    wire N__11057;
    wire N__11056;
    wire N__11049;
    wire N__11048;
    wire N__11047;
    wire N__11030;
    wire N__11029;
    wire N__11028;
    wire N__11027;
    wire N__11024;
    wire N__11021;
    wire N__11018;
    wire N__11015;
    wire N__11014;
    wire N__11013;
    wire N__11012;
    wire N__11009;
    wire N__11008;
    wire N__11007;
    wire N__11004;
    wire N__11003;
    wire N__11002;
    wire N__11001;
    wire N__11000;
    wire N__10999;
    wire N__10996;
    wire N__10995;
    wire N__10994;
    wire N__10993;
    wire N__10992;
    wire N__10991;
    wire N__10990;
    wire N__10989;
    wire N__10988;
    wire N__10987;
    wire N__10984;
    wire N__10983;
    wire N__10982;
    wire N__10981;
    wire N__10980;
    wire N__10979;
    wire N__10978;
    wire N__10977;
    wire N__10976;
    wire N__10975;
    wire N__10974;
    wire N__10973;
    wire N__10972;
    wire N__10901;
    wire N__10898;
    wire N__10895;
    wire N__10892;
    wire N__10889;
    wire N__10886;
    wire N__10883;
    wire N__10880;
    wire N__10879;
    wire N__10876;
    wire N__10873;
    wire N__10868;
    wire N__10865;
    wire N__10864;
    wire N__10861;
    wire N__10858;
    wire N__10857;
    wire N__10854;
    wire N__10851;
    wire N__10848;
    wire N__10841;
    wire N__10838;
    wire N__10837;
    wire N__10836;
    wire N__10833;
    wire N__10832;
    wire N__10829;
    wire N__10826;
    wire N__10823;
    wire N__10820;
    wire N__10817;
    wire N__10814;
    wire N__10809;
    wire N__10806;
    wire N__10803;
    wire N__10800;
    wire N__10797;
    wire N__10794;
    wire N__10791;
    wire N__10784;
    wire N__10783;
    wire N__10782;
    wire N__10779;
    wire N__10776;
    wire N__10775;
    wire N__10772;
    wire N__10767;
    wire N__10764;
    wire N__10763;
    wire N__10760;
    wire N__10755;
    wire N__10752;
    wire N__10749;
    wire N__10744;
    wire N__10741;
    wire N__10740;
    wire N__10737;
    wire N__10734;
    wire N__10731;
    wire N__10728;
    wire N__10723;
    wire N__10718;
    wire N__10715;
    wire N__10712;
    wire N__10709;
    wire N__10706;
    wire N__10703;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10693;
    wire N__10692;
    wire N__10691;
    wire N__10690;
    wire N__10687;
    wire N__10686;
    wire N__10683;
    wire N__10680;
    wire N__10679;
    wire N__10678;
    wire N__10675;
    wire N__10674;
    wire N__10673;
    wire N__10672;
    wire N__10671;
    wire N__10670;
    wire N__10667;
    wire N__10664;
    wire N__10661;
    wire N__10656;
    wire N__10655;
    wire N__10654;
    wire N__10651;
    wire N__10648;
    wire N__10647;
    wire N__10646;
    wire N__10645;
    wire N__10642;
    wire N__10641;
    wire N__10640;
    wire N__10639;
    wire N__10636;
    wire N__10635;
    wire N__10626;
    wire N__10617;
    wire N__10612;
    wire N__10607;
    wire N__10604;
    wire N__10599;
    wire N__10596;
    wire N__10591;
    wire N__10588;
    wire N__10585;
    wire N__10582;
    wire N__10575;
    wire N__10574;
    wire N__10573;
    wire N__10570;
    wire N__10567;
    wire N__10564;
    wire N__10555;
    wire N__10552;
    wire N__10549;
    wire N__10546;
    wire N__10543;
    wire N__10536;
    wire N__10533;
    wire N__10528;
    wire N__10517;
    wire N__10516;
    wire N__10513;
    wire N__10510;
    wire N__10505;
    wire N__10502;
    wire N__10499;
    wire N__10496;
    wire N__10493;
    wire N__10490;
    wire N__10487;
    wire N__10484;
    wire N__10481;
    wire N__10478;
    wire N__10475;
    wire N__10472;
    wire N__10469;
    wire N__10466;
    wire N__10463;
    wire N__10460;
    wire N__10457;
    wire N__10454;
    wire N__10451;
    wire N__10448;
    wire N__10445;
    wire N__10442;
    wire N__10439;
    wire N__10436;
    wire N__10433;
    wire N__10430;
    wire N__10427;
    wire N__10424;
    wire N__10423;
    wire N__10420;
    wire N__10417;
    wire N__10416;
    wire N__10413;
    wire N__10408;
    wire N__10407;
    wire N__10406;
    wire N__10405;
    wire N__10404;
    wire N__10403;
    wire N__10400;
    wire N__10397;
    wire N__10394;
    wire N__10385;
    wire N__10382;
    wire N__10377;
    wire N__10374;
    wire N__10371;
    wire N__10368;
    wire N__10365;
    wire N__10362;
    wire N__10357;
    wire N__10354;
    wire N__10349;
    wire N__10348;
    wire N__10347;
    wire N__10342;
    wire N__10339;
    wire N__10338;
    wire N__10337;
    wire N__10336;
    wire N__10335;
    wire N__10332;
    wire N__10329;
    wire N__10320;
    wire N__10319;
    wire N__10316;
    wire N__10313;
    wire N__10310;
    wire N__10307;
    wire N__10300;
    wire N__10297;
    wire N__10294;
    wire N__10291;
    wire N__10286;
    wire N__10283;
    wire N__10282;
    wire N__10281;
    wire N__10278;
    wire N__10277;
    wire N__10276;
    wire N__10273;
    wire N__10272;
    wire N__10269;
    wire N__10260;
    wire N__10259;
    wire N__10258;
    wire N__10255;
    wire N__10252;
    wire N__10251;
    wire N__10248;
    wire N__10245;
    wire N__10244;
    wire N__10239;
    wire N__10236;
    wire N__10233;
    wire N__10230;
    wire N__10227;
    wire N__10224;
    wire N__10217;
    wire N__10214;
    wire N__10209;
    wire N__10206;
    wire N__10203;
    wire N__10200;
    wire N__10197;
    wire N__10192;
    wire N__10187;
    wire N__10186;
    wire N__10185;
    wire N__10182;
    wire N__10181;
    wire N__10180;
    wire N__10179;
    wire N__10174;
    wire N__10171;
    wire N__10168;
    wire N__10167;
    wire N__10164;
    wire N__10161;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10151;
    wire N__10142;
    wire N__10141;
    wire N__10134;
    wire N__10131;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10121;
    wire N__10118;
    wire N__10115;
    wire N__10112;
    wire N__10107;
    wire N__10104;
    wire N__10097;
    wire N__10094;
    wire N__10091;
    wire N__10088;
    wire N__10085;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10075;
    wire N__10072;
    wire N__10069;
    wire N__10068;
    wire N__10067;
    wire N__10062;
    wire N__10059;
    wire N__10056;
    wire N__10053;
    wire N__10050;
    wire N__10047;
    wire N__10042;
    wire N__10039;
    wire N__10036;
    wire N__10033;
    wire N__10030;
    wire N__10025;
    wire N__10024;
    wire N__10023;
    wire N__10020;
    wire N__10019;
    wire N__10016;
    wire N__10013;
    wire N__10010;
    wire N__10007;
    wire N__10004;
    wire N__10001;
    wire N__9996;
    wire N__9993;
    wire N__9988;
    wire N__9985;
    wire N__9982;
    wire N__9979;
    wire N__9974;
    wire N__9971;
    wire N__9970;
    wire N__9969;
    wire N__9968;
    wire N__9965;
    wire N__9962;
    wire N__9961;
    wire N__9960;
    wire N__9959;
    wire N__9956;
    wire N__9955;
    wire N__9952;
    wire N__9951;
    wire N__9950;
    wire N__9949;
    wire N__9948;
    wire N__9945;
    wire N__9942;
    wire N__9939;
    wire N__9934;
    wire N__9933;
    wire N__9932;
    wire N__9929;
    wire N__9926;
    wire N__9925;
    wire N__9924;
    wire N__9921;
    wire N__9912;
    wire N__9911;
    wire N__9910;
    wire N__9909;
    wire N__9908;
    wire N__9907;
    wire N__9904;
    wire N__9897;
    wire N__9892;
    wire N__9889;
    wire N__9886;
    wire N__9881;
    wire N__9876;
    wire N__9867;
    wire N__9864;
    wire N__9857;
    wire N__9854;
    wire N__9851;
    wire N__9848;
    wire N__9839;
    wire N__9834;
    wire N__9831;
    wire N__9828;
    wire N__9825;
    wire N__9820;
    wire N__9817;
    wire N__9812;
    wire N__9809;
    wire N__9806;
    wire N__9803;
    wire N__9800;
    wire N__9799;
    wire N__9798;
    wire N__9797;
    wire N__9796;
    wire N__9785;
    wire N__9782;
    wire N__9779;
    wire N__9778;
    wire N__9777;
    wire N__9776;
    wire N__9775;
    wire N__9774;
    wire N__9773;
    wire N__9772;
    wire N__9771;
    wire N__9770;
    wire N__9749;
    wire N__9746;
    wire N__9743;
    wire N__9740;
    wire N__9739;
    wire N__9738;
    wire N__9737;
    wire N__9736;
    wire N__9735;
    wire N__9734;
    wire N__9733;
    wire N__9732;
    wire N__9731;
    wire N__9730;
    wire N__9729;
    wire N__9728;
    wire N__9727;
    wire N__9726;
    wire N__9725;
    wire N__9724;
    wire N__9723;
    wire N__9720;
    wire N__9719;
    wire N__9718;
    wire N__9717;
    wire N__9716;
    wire N__9715;
    wire N__9714;
    wire N__9713;
    wire N__9662;
    wire N__9659;
    wire N__9656;
    wire N__9655;
    wire N__9654;
    wire N__9651;
    wire N__9648;
    wire N__9647;
    wire N__9644;
    wire N__9639;
    wire N__9636;
    wire N__9631;
    wire N__9628;
    wire N__9623;
    wire N__9620;
    wire N__9617;
    wire N__9614;
    wire N__9613;
    wire N__9612;
    wire N__9611;
    wire N__9608;
    wire N__9603;
    wire N__9600;
    wire N__9597;
    wire N__9592;
    wire N__9589;
    wire N__9586;
    wire N__9583;
    wire N__9580;
    wire N__9577;
    wire N__9574;
    wire N__9569;
    wire N__9568;
    wire N__9563;
    wire N__9560;
    wire N__9557;
    wire N__9554;
    wire N__9553;
    wire N__9550;
    wire N__9547;
    wire N__9546;
    wire N__9541;
    wire N__9538;
    wire N__9537;
    wire N__9532;
    wire N__9529;
    wire N__9526;
    wire N__9523;
    wire N__9520;
    wire N__9517;
    wire N__9514;
    wire N__9511;
    wire N__9508;
    wire N__9503;
    wire N__9500;
    wire N__9497;
    wire N__9494;
    wire N__9491;
    wire N__9488;
    wire N__9485;
    wire N__9484;
    wire N__9481;
    wire N__9478;
    wire N__9477;
    wire N__9476;
    wire N__9473;
    wire N__9470;
    wire N__9465;
    wire N__9462;
    wire N__9459;
    wire N__9456;
    wire N__9451;
    wire N__9448;
    wire N__9445;
    wire N__9442;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9422;
    wire N__9419;
    wire N__9416;
    wire N__9413;
    wire N__9410;
    wire N__9407;
    wire N__9406;
    wire N__9403;
    wire N__9400;
    wire N__9399;
    wire N__9398;
    wire N__9393;
    wire N__9388;
    wire N__9383;
    wire N__9380;
    wire N__9377;
    wire N__9374;
    wire N__9371;
    wire N__9368;
    wire N__9365;
    wire N__9362;
    wire N__9359;
    wire N__9358;
    wire N__9357;
    wire N__9352;
    wire N__9351;
    wire N__9348;
    wire N__9345;
    wire N__9342;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9326;
    wire N__9325;
    wire N__9324;
    wire N__9323;
    wire N__9318;
    wire N__9315;
    wire N__9312;
    wire N__9309;
    wire N__9304;
    wire N__9301;
    wire N__9298;
    wire N__9295;
    wire N__9292;
    wire N__9289;
    wire N__9286;
    wire N__9281;
    wire N__9278;
    wire N__9275;
    wire N__9272;
    wire N__9269;
    wire N__9266;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9242;
    wire N__9239;
    wire N__9236;
    wire N__9233;
    wire N__9230;
    wire N__9227;
    wire N__9224;
    wire N__9221;
    wire N__9218;
    wire N__9215;
    wire N__9212;
    wire N__9209;
    wire N__9206;
    wire N__9203;
    wire N__9200;
    wire N__9197;
    wire N__9194;
    wire N__9191;
    wire N__9190;
    wire N__9187;
    wire N__9184;
    wire N__9183;
    wire N__9180;
    wire N__9177;
    wire N__9174;
    wire N__9173;
    wire N__9172;
    wire N__9171;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9140;
    wire N__9139;
    wire N__9138;
    wire N__9137;
    wire N__9136;
    wire N__9135;
    wire N__9134;
    wire N__9131;
    wire N__9128;
    wire N__9125;
    wire N__9124;
    wire N__9123;
    wire N__9122;
    wire N__9119;
    wire N__9118;
    wire N__9117;
    wire N__9116;
    wire N__9113;
    wire N__9110;
    wire N__9107;
    wire N__9104;
    wire N__9097;
    wire N__9094;
    wire N__9091;
    wire N__9090;
    wire N__9087;
    wire N__9080;
    wire N__9077;
    wire N__9076;
    wire N__9075;
    wire N__9072;
    wire N__9069;
    wire N__9068;
    wire N__9067;
    wire N__9066;
    wire N__9059;
    wire N__9054;
    wire N__9047;
    wire N__9044;
    wire N__9041;
    wire N__9040;
    wire N__9039;
    wire N__9038;
    wire N__9037;
    wire N__9032;
    wire N__9025;
    wire N__9020;
    wire N__9017;
    wire N__9014;
    wire N__9011;
    wire N__9002;
    wire N__8997;
    wire N__8994;
    wire N__8981;
    wire N__8980;
    wire N__8979;
    wire N__8976;
    wire N__8973;
    wire N__8972;
    wire N__8969;
    wire N__8966;
    wire N__8963;
    wire N__8960;
    wire N__8955;
    wire N__8952;
    wire N__8949;
    wire N__8946;
    wire N__8941;
    wire N__8936;
    wire N__8935;
    wire N__8932;
    wire N__8929;
    wire N__8928;
    wire N__8923;
    wire N__8920;
    wire N__8919;
    wire N__8916;
    wire N__8915;
    wire N__8914;
    wire N__8911;
    wire N__8908;
    wire N__8905;
    wire N__8902;
    wire N__8899;
    wire N__8894;
    wire N__8885;
    wire N__8882;
    wire N__8879;
    wire N__8876;
    wire N__8873;
    wire N__8870;
    wire N__8867;
    wire N__8864;
    wire N__8861;
    wire N__8858;
    wire N__8855;
    wire N__8852;
    wire N__8849;
    wire N__8846;
    wire N__8843;
    wire N__8840;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8828;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire N__8801;
    wire N__8798;
    wire N__8795;
    wire N__8792;
    wire N__8789;
    wire N__8786;
    wire N__8783;
    wire N__8780;
    wire N__8779;
    wire N__8778;
    wire N__8777;
    wire N__8776;
    wire N__8775;
    wire N__8774;
    wire N__8773;
    wire N__8770;
    wire N__8765;
    wire N__8762;
    wire N__8757;
    wire N__8754;
    wire N__8751;
    wire N__8750;
    wire N__8741;
    wire N__8734;
    wire N__8729;
    wire N__8728;
    wire N__8727;
    wire N__8726;
    wire N__8725;
    wire N__8722;
    wire N__8719;
    wire N__8718;
    wire N__8715;
    wire N__8712;
    wire N__8705;
    wire N__8698;
    wire N__8693;
    wire N__8690;
    wire N__8687;
    wire N__8684;
    wire N__8681;
    wire N__8678;
    wire N__8675;
    wire N__8672;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8641;
    wire N__8638;
    wire N__8635;
    wire N__8634;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8622;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8600;
    wire N__8597;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8584;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8570;
    wire N__8567;
    wire N__8564;
    wire N__8563;
    wire N__8558;
    wire N__8557;
    wire N__8556;
    wire N__8553;
    wire N__8548;
    wire N__8545;
    wire N__8542;
    wire N__8539;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8522;
    wire N__8521;
    wire N__8518;
    wire N__8515;
    wire N__8510;
    wire N__8507;
    wire N__8504;
    wire N__8501;
    wire N__8498;
    wire N__8495;
    wire N__8492;
    wire N__8491;
    wire N__8490;
    wire N__8489;
    wire N__8488;
    wire N__8485;
    wire N__8484;
    wire N__8481;
    wire N__8480;
    wire N__8479;
    wire N__8476;
    wire N__8469;
    wire N__8466;
    wire N__8463;
    wire N__8458;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8438;
    wire N__8435;
    wire N__8432;
    wire N__8429;
    wire N__8428;
    wire N__8425;
    wire N__8422;
    wire N__8421;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8399;
    wire N__8398;
    wire N__8395;
    wire N__8394;
    wire N__8393;
    wire N__8392;
    wire N__8385;
    wire N__8382;
    wire N__8379;
    wire N__8378;
    wire N__8377;
    wire N__8376;
    wire N__8375;
    wire N__8370;
    wire N__8367;
    wire N__8364;
    wire N__8359;
    wire N__8356;
    wire N__8353;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8333;
    wire N__8332;
    wire N__8331;
    wire N__8328;
    wire N__8327;
    wire N__8326;
    wire N__8323;
    wire N__8320;
    wire N__8319;
    wire N__8318;
    wire N__8317;
    wire N__8314;
    wire N__8309;
    wire N__8306;
    wire N__8303;
    wire N__8300;
    wire N__8295;
    wire N__8282;
    wire N__8281;
    wire N__8280;
    wire N__8277;
    wire N__8274;
    wire N__8271;
    wire N__8268;
    wire N__8261;
    wire N__8260;
    wire N__8259;
    wire N__8256;
    wire N__8255;
    wire N__8252;
    wire N__8251;
    wire N__8250;
    wire N__8249;
    wire N__8246;
    wire N__8243;
    wire N__8240;
    wire N__8237;
    wire N__8234;
    wire N__8229;
    wire N__8216;
    wire N__8215;
    wire N__8214;
    wire N__8213;
    wire N__8210;
    wire N__8203;
    wire N__8198;
    wire N__8195;
    wire N__8192;
    wire N__8189;
    wire N__8186;
    wire N__8183;
    wire N__8180;
    wire N__8177;
    wire N__8174;
    wire N__8171;
    wire N__8168;
    wire N__8165;
    wire N__8162;
    wire N__8159;
    wire N__8156;
    wire N__8153;
    wire N__8150;
    wire N__8147;
    wire N__8144;
    wire N__8141;
    wire N__8138;
    wire N__8135;
    wire N__8132;
    wire N__8129;
    wire N__8126;
    wire N__8123;
    wire N__8120;
    wire N__8117;
    wire N__8114;
    wire N__8111;
    wire N__8108;
    wire N__8105;
    wire N__8102;
    wire N__8099;
    wire N__8096;
    wire N__8093;
    wire N__8090;
    wire N__8087;
    wire N__8086;
    wire N__8085;
    wire N__8084;
    wire N__8083;
    wire N__8080;
    wire N__8077;
    wire N__8076;
    wire N__8073;
    wire N__8068;
    wire N__8063;
    wire N__8060;
    wire N__8051;
    wire N__8048;
    wire N__8045;
    wire N__8044;
    wire N__8041;
    wire N__8038;
    wire N__8035;
    wire N__8032;
    wire N__8029;
    wire N__8026;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8012;
    wire N__8011;
    wire N__8008;
    wire N__8005;
    wire N__8002;
    wire N__7999;
    wire N__7996;
    wire N__7993;
    wire N__7990;
    wire N__7987;
    wire N__7984;
    wire N__7981;
    wire N__7978;
    wire N__7975;
    wire N__7970;
    wire N__7969;
    wire N__7964;
    wire N__7961;
    wire N__7958;
    wire N__7957;
    wire N__7954;
    wire N__7951;
    wire N__7950;
    wire N__7947;
    wire N__7944;
    wire N__7941;
    wire N__7934;
    wire N__7931;
    wire N__7928;
    wire N__7927;
    wire N__7926;
    wire N__7923;
    wire N__7920;
    wire N__7919;
    wire N__7916;
    wire N__7913;
    wire N__7910;
    wire N__7905;
    wire N__7900;
    wire N__7897;
    wire N__7894;
    wire N__7891;
    wire N__7888;
    wire N__7885;
    wire N__7880;
    wire N__7879;
    wire N__7876;
    wire N__7875;
    wire N__7874;
    wire N__7873;
    wire N__7870;
    wire N__7867;
    wire N__7862;
    wire N__7859;
    wire N__7856;
    wire N__7851;
    wire N__7844;
    wire N__7841;
    wire N__7838;
    wire N__7835;
    wire N__7832;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7814;
    wire N__7811;
    wire N__7808;
    wire N__7805;
    wire N__7802;
    wire N__7799;
    wire N__7798;
    wire N__7795;
    wire N__7792;
    wire N__7787;
    wire N__7784;
    wire N__7783;
    wire N__7780;
    wire N__7777;
    wire N__7772;
    wire N__7769;
    wire N__7768;
    wire N__7765;
    wire N__7762;
    wire N__7757;
    wire N__7754;
    wire N__7753;
    wire N__7750;
    wire N__7747;
    wire N__7744;
    wire N__7739;
    wire N__7736;
    wire N__7735;
    wire N__7732;
    wire N__7729;
    wire N__7726;
    wire N__7721;
    wire N__7718;
    wire N__7717;
    wire N__7714;
    wire N__7711;
    wire N__7708;
    wire N__7703;
    wire N__7700;
    wire N__7697;
    wire N__7694;
    wire N__7693;
    wire N__7690;
    wire N__7687;
    wire N__7684;
    wire N__7679;
    wire N__7678;
    wire N__7677;
    wire N__7676;
    wire N__7675;
    wire N__7674;
    wire N__7673;
    wire N__7658;
    wire N__7655;
    wire N__7652;
    wire N__7649;
    wire N__7646;
    wire N__7643;
    wire N__7640;
    wire N__7637;
    wire N__7634;
    wire N__7633;
    wire N__7630;
    wire N__7627;
    wire N__7622;
    wire N__7619;
    wire N__7616;
    wire N__7613;
    wire N__7610;
    wire N__7607;
    wire N__7604;
    wire N__7601;
    wire N__7598;
    wire N__7595;
    wire N__7592;
    wire N__7589;
    wire N__7586;
    wire N__7583;
    wire N__7580;
    wire N__7577;
    wire N__7574;
    wire N__7571;
    wire N__7568;
    wire N__7565;
    wire N__7562;
    wire N__7559;
    wire N__7556;
    wire N__7553;
    wire N__7550;
    wire N__7547;
    wire N__7544;
    wire N__7541;
    wire N__7538;
    wire N__7535;
    wire N__7532;
    wire N__7529;
    wire N__7526;
    wire N__7523;
    wire N__7520;
    wire N__7517;
    wire N__7516;
    wire N__7513;
    wire N__7510;
    wire N__7507;
    wire N__7504;
    wire N__7501;
    wire N__7498;
    wire N__7495;
    wire N__7492;
    wire N__7489;
    wire N__7486;
    wire N__7481;
    wire N__7478;
    wire N__7475;
    wire N__7472;
    wire N__7469;
    wire N__7466;
    wire N__7463;
    wire N__7460;
    wire N__7457;
    wire N__7454;
    wire N__7451;
    wire N__7448;
    wire N__7445;
    wire N__7442;
    wire N__7441;
    wire N__7438;
    wire N__7435;
    wire N__7430;
    wire N__7427;
    wire N__7426;
    wire N__7423;
    wire N__7420;
    wire N__7419;
    wire N__7418;
    wire N__7417;
    wire N__7416;
    wire N__7411;
    wire N__7410;
    wire N__7407;
    wire N__7406;
    wire N__7401;
    wire N__7398;
    wire N__7395;
    wire N__7392;
    wire N__7389;
    wire N__7386;
    wire N__7381;
    wire N__7370;
    wire N__7367;
    wire N__7364;
    wire N__7361;
    wire N__7358;
    wire N__7355;
    wire N__7352;
    wire N__7349;
    wire N__7346;
    wire N__7343;
    wire N__7340;
    wire N__7337;
    wire N__7336;
    wire N__7335;
    wire N__7334;
    wire N__7331;
    wire N__7328;
    wire N__7325;
    wire N__7322;
    wire N__7313;
    wire N__7310;
    wire N__7307;
    wire N__7304;
    wire N__7301;
    wire N__7298;
    wire N__7295;
    wire N__7292;
    wire N__7289;
    wire N__7286;
    wire N__7283;
    wire N__7280;
    wire N__7277;
    wire N__7274;
    wire N__7271;
    wire N__7268;
    wire N__7265;
    wire N__7262;
    wire N__7259;
    wire N__7256;
    wire N__7253;
    wire N__7250;
    wire N__7247;
    wire N__7244;
    wire N__7241;
    wire N__7238;
    wire N__7235;
    wire N__7232;
    wire N__7229;
    wire N__7226;
    wire N__7223;
    wire N__7220;
    wire N__7217;
    wire N__7214;
    wire N__7213;
    wire N__7210;
    wire N__7207;
    wire N__7206;
    wire N__7205;
    wire N__7204;
    wire N__7203;
    wire N__7200;
    wire N__7197;
    wire N__7192;
    wire N__7187;
    wire N__7178;
    wire N__7175;
    wire N__7174;
    wire N__7171;
    wire N__7168;
    wire N__7163;
    wire N__7162;
    wire N__7157;
    wire N__7154;
    wire N__7151;
    wire N__7148;
    wire N__7145;
    wire N__7142;
    wire N__7139;
    wire N__7136;
    wire N__7133;
    wire N__7132;
    wire N__7129;
    wire N__7126;
    wire N__7123;
    wire N__7120;
    wire N__7117;
    wire N__7114;
    wire N__7109;
    wire N__7106;
    wire N__7103;
    wire N__7100;
    wire N__7097;
    wire N__7096;
    wire N__7091;
    wire N__7088;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7076;
    wire N__7073;
    wire N__7070;
    wire N__7067;
    wire N__7064;
    wire N__7061;
    wire N__7058;
    wire N__7055;
    wire N__7052;
    wire N__7049;
    wire N__7046;
    wire N__7043;
    wire N__7040;
    wire N__7039;
    wire N__7036;
    wire N__7033;
    wire N__7032;
    wire N__7031;
    wire N__7026;
    wire N__7023;
    wire N__7020;
    wire N__7013;
    wire N__7012;
    wire N__7009;
    wire N__7008;
    wire N__7005;
    wire N__7002;
    wire N__7001;
    wire N__7000;
    wire N__6997;
    wire N__6994;
    wire N__6991;
    wire N__6988;
    wire N__6987;
    wire N__6984;
    wire N__6981;
    wire N__6976;
    wire N__6973;
    wire N__6970;
    wire N__6967;
    wire N__6956;
    wire N__6953;
    wire N__6950;
    wire N__6947;
    wire N__6944;
    wire N__6943;
    wire N__6940;
    wire N__6937;
    wire N__6932;
    wire N__6929;
    wire N__6926;
    wire N__6923;
    wire N__6920;
    wire N__6917;
    wire N__6914;
    wire N__6911;
    wire N__6908;
    wire N__6905;
    wire N__6904;
    wire N__6899;
    wire N__6896;
    wire N__6893;
    wire N__6890;
    wire N__6887;
    wire N__6884;
    wire N__6881;
    wire N__6880;
    wire N__6879;
    wire N__6878;
    wire N__6875;
    wire N__6872;
    wire N__6869;
    wire N__6866;
    wire N__6865;
    wire N__6862;
    wire N__6857;
    wire N__6854;
    wire N__6851;
    wire N__6848;
    wire N__6843;
    wire N__6836;
    wire N__6835;
    wire N__6834;
    wire N__6831;
    wire N__6828;
    wire N__6825;
    wire N__6818;
    wire N__6815;
    wire N__6812;
    wire N__6811;
    wire N__6808;
    wire N__6805;
    wire N__6800;
    wire N__6799;
    wire N__6798;
    wire N__6793;
    wire N__6790;
    wire N__6785;
    wire N__6784;
    wire N__6781;
    wire N__6780;
    wire N__6777;
    wire N__6774;
    wire N__6771;
    wire N__6764;
    wire N__6761;
    wire N__6760;
    wire N__6757;
    wire N__6754;
    wire N__6753;
    wire N__6748;
    wire N__6745;
    wire N__6740;
    wire N__6739;
    wire N__6738;
    wire N__6737;
    wire N__6736;
    wire N__6735;
    wire N__6734;
    wire N__6731;
    wire N__6730;
    wire N__6729;
    wire N__6726;
    wire N__6721;
    wire N__6720;
    wire N__6719;
    wire N__6716;
    wire N__6711;
    wire N__6708;
    wire N__6703;
    wire N__6698;
    wire N__6695;
    wire N__6694;
    wire N__6693;
    wire N__6692;
    wire N__6689;
    wire N__6688;
    wire N__6687;
    wire N__6682;
    wire N__6677;
    wire N__6672;
    wire N__6665;
    wire N__6660;
    wire N__6657;
    wire N__6644;
    wire N__6641;
    wire N__6638;
    wire N__6635;
    wire N__6632;
    wire N__6629;
    wire N__6628;
    wire N__6627;
    wire N__6626;
    wire N__6623;
    wire N__6622;
    wire N__6621;
    wire N__6620;
    wire N__6619;
    wire N__6618;
    wire N__6617;
    wire N__6614;
    wire N__6613;
    wire N__6610;
    wire N__6607;
    wire N__6606;
    wire N__6603;
    wire N__6600;
    wire N__6599;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6583;
    wire N__6582;
    wire N__6581;
    wire N__6578;
    wire N__6575;
    wire N__6572;
    wire N__6571;
    wire N__6568;
    wire N__6567;
    wire N__6562;
    wire N__6559;
    wire N__6554;
    wire N__6551;
    wire N__6548;
    wire N__6543;
    wire N__6536;
    wire N__6533;
    wire N__6530;
    wire N__6527;
    wire N__6518;
    wire N__6503;
    wire N__6500;
    wire N__6497;
    wire N__6496;
    wire N__6495;
    wire N__6494;
    wire N__6491;
    wire N__6490;
    wire N__6489;
    wire N__6482;
    wire N__6479;
    wire N__6476;
    wire N__6475;
    wire N__6474;
    wire N__6473;
    wire N__6472;
    wire N__6471;
    wire N__6468;
    wire N__6461;
    wire N__6456;
    wire N__6453;
    wire N__6450;
    wire N__6447;
    wire N__6446;
    wire N__6445;
    wire N__6442;
    wire N__6439;
    wire N__6430;
    wire N__6425;
    wire N__6416;
    wire N__6415;
    wire N__6412;
    wire N__6409;
    wire N__6408;
    wire N__6407;
    wire N__6406;
    wire N__6405;
    wire N__6404;
    wire N__6403;
    wire N__6398;
    wire N__6393;
    wire N__6390;
    wire N__6389;
    wire N__6388;
    wire N__6385;
    wire N__6382;
    wire N__6379;
    wire N__6374;
    wire N__6373;
    wire N__6372;
    wire N__6371;
    wire N__6370;
    wire N__6367;
    wire N__6364;
    wire N__6361;
    wire N__6360;
    wire N__6359;
    wire N__6358;
    wire N__6355;
    wire N__6352;
    wire N__6349;
    wire N__6346;
    wire N__6341;
    wire N__6336;
    wire N__6329;
    wire N__6322;
    wire N__6305;
    wire N__6302;
    wire N__6299;
    wire N__6298;
    wire N__6297;
    wire N__6296;
    wire N__6295;
    wire N__6294;
    wire N__6293;
    wire N__6290;
    wire N__6287;
    wire N__6282;
    wire N__6277;
    wire N__6276;
    wire N__6273;
    wire N__6270;
    wire N__6269;
    wire N__6268;
    wire N__6267;
    wire N__6266;
    wire N__6259;
    wire N__6256;
    wire N__6253;
    wire N__6250;
    wire N__6245;
    wire N__6240;
    wire N__6235;
    wire N__6224;
    wire N__6223;
    wire N__6222;
    wire N__6221;
    wire N__6218;
    wire N__6215;
    wire N__6214;
    wire N__6213;
    wire N__6212;
    wire N__6211;
    wire N__6208;
    wire N__6207;
    wire N__6204;
    wire N__6203;
    wire N__6202;
    wire N__6201;
    wire N__6200;
    wire N__6197;
    wire N__6196;
    wire N__6195;
    wire N__6194;
    wire N__6193;
    wire N__6192;
    wire N__6189;
    wire N__6184;
    wire N__6181;
    wire N__6176;
    wire N__6173;
    wire N__6170;
    wire N__6165;
    wire N__6162;
    wire N__6161;
    wire N__6160;
    wire N__6157;
    wire N__6154;
    wire N__6147;
    wire N__6142;
    wire N__6133;
    wire N__6124;
    wire N__6121;
    wire N__6118;
    wire N__6101;
    wire N__6098;
    wire N__6097;
    wire N__6096;
    wire N__6095;
    wire N__6094;
    wire N__6093;
    wire N__6090;
    wire N__6087;
    wire N__6084;
    wire N__6081;
    wire N__6078;
    wire N__6077;
    wire N__6076;
    wire N__6073;
    wire N__6070;
    wire N__6067;
    wire N__6064;
    wire N__6057;
    wire N__6054;
    wire N__6041;
    wire N__6038;
    wire N__6035;
    wire N__6032;
    wire N__6029;
    wire N__6026;
    wire N__6023;
    wire N__6020;
    wire N__6017;
    wire N__6014;
    wire N__6011;
    wire N__6008;
    wire N__6005;
    wire N__6002;
    wire N__5999;
    wire N__5996;
    wire N__5993;
    wire N__5990;
    wire N__5987;
    wire N__5984;
    wire N__5981;
    wire N__5978;
    wire N__5975;
    wire N__5974;
    wire N__5971;
    wire N__5970;
    wire N__5967;
    wire N__5960;
    wire N__5957;
    wire N__5954;
    wire N__5953;
    wire N__5952;
    wire N__5951;
    wire N__5948;
    wire N__5941;
    wire N__5936;
    wire N__5935;
    wire N__5932;
    wire N__5929;
    wire N__5926;
    wire N__5923;
    wire N__5920;
    wire N__5917;
    wire N__5912;
    wire N__5909;
    wire N__5908;
    wire N__5907;
    wire N__5906;
    wire N__5905;
    wire N__5904;
    wire N__5901;
    wire N__5900;
    wire N__5897;
    wire N__5894;
    wire N__5893;
    wire N__5892;
    wire N__5891;
    wire N__5888;
    wire N__5885;
    wire N__5882;
    wire N__5879;
    wire N__5876;
    wire N__5873;
    wire N__5870;
    wire N__5863;
    wire N__5846;
    wire N__5843;
    wire N__5840;
    wire N__5839;
    wire N__5836;
    wire N__5835;
    wire N__5834;
    wire N__5833;
    wire N__5832;
    wire N__5829;
    wire N__5826;
    wire N__5823;
    wire N__5818;
    wire N__5813;
    wire N__5804;
    wire N__5801;
    wire N__5800;
    wire N__5797;
    wire N__5794;
    wire N__5789;
    wire N__5788;
    wire N__5785;
    wire N__5784;
    wire N__5781;
    wire N__5778;
    wire N__5775;
    wire N__5768;
    wire N__5765;
    wire N__5762;
    wire N__5759;
    wire N__5756;
    wire N__5755;
    wire N__5752;
    wire N__5749;
    wire N__5744;
    wire N__5741;
    wire N__5738;
    wire N__5737;
    wire N__5734;
    wire N__5731;
    wire N__5726;
    wire N__5723;
    wire N__5720;
    wire N__5717;
    wire N__5714;
    wire N__5711;
    wire N__5708;
    wire N__5705;
    wire N__5702;
    wire N__5699;
    wire N__5698;
    wire N__5693;
    wire N__5690;
    wire N__5687;
    wire N__5684;
    wire N__5681;
    wire N__5680;
    wire N__5677;
    wire N__5674;
    wire N__5671;
    wire N__5668;
    wire N__5663;
    wire N__5662;
    wire N__5659;
    wire N__5656;
    wire N__5651;
    wire N__5648;
    wire N__5645;
    wire N__5642;
    wire N__5639;
    wire N__5638;
    wire N__5635;
    wire N__5632;
    wire N__5629;
    wire N__5626;
    wire N__5623;
    wire N__5618;
    wire N__5617;
    wire N__5614;
    wire N__5611;
    wire N__5608;
    wire N__5607;
    wire N__5604;
    wire N__5601;
    wire N__5600;
    wire N__5597;
    wire N__5592;
    wire N__5589;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5570;
    wire N__5567;
    wire N__5566;
    wire N__5563;
    wire N__5560;
    wire N__5555;
    wire N__5552;
    wire N__5549;
    wire N__5546;
    wire N__5545;
    wire N__5542;
    wire N__5539;
    wire N__5534;
    wire N__5531;
    wire N__5528;
    wire N__5525;
    wire N__5524;
    wire N__5521;
    wire N__5518;
    wire N__5515;
    wire N__5512;
    wire N__5509;
    wire N__5506;
    wire N__5501;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5489;
    wire N__5486;
    wire N__5483;
    wire N__5480;
    wire N__5477;
    wire N__5476;
    wire N__5473;
    wire N__5470;
    wire N__5465;
    wire N__5462;
    wire N__5461;
    wire N__5458;
    wire N__5455;
    wire N__5450;
    wire N__5447;
    wire N__5444;
    wire N__5441;
    wire N__5438;
    wire N__5435;
    wire N__5432;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5396;
    wire N__5393;
    wire N__5390;
    wire N__5387;
    wire N__5384;
    wire N__5381;
    wire N__5378;
    wire N__5375;
    wire N__5372;
    wire N__5369;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5354;
    wire N__5351;
    wire N__5350;
    wire N__5347;
    wire N__5344;
    wire N__5341;
    wire N__5340;
    wire N__5339;
    wire N__5336;
    wire N__5333;
    wire N__5330;
    wire N__5327;
    wire N__5318;
    wire N__5315;
    wire N__5312;
    wire N__5309;
    wire N__5306;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5294;
    wire N__5291;
    wire N__5288;
    wire N__5285;
    wire N__5282;
    wire N__5279;
    wire N__5276;
    wire N__5273;
    wire N__5270;
    wire N__5267;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5255;
    wire N__5254;
    wire N__5251;
    wire N__5248;
    wire N__5245;
    wire N__5240;
    wire N__5237;
    wire N__5236;
    wire N__5235;
    wire N__5232;
    wire N__5227;
    wire N__5224;
    wire N__5219;
    wire N__5216;
    wire N__5215;
    wire N__5214;
    wire N__5211;
    wire N__5210;
    wire N__5209;
    wire N__5208;
    wire N__5207;
    wire N__5206;
    wire N__5205;
    wire N__5204;
    wire N__5201;
    wire N__5200;
    wire N__5197;
    wire N__5194;
    wire N__5189;
    wire N__5188;
    wire N__5187;
    wire N__5186;
    wire N__5185;
    wire N__5184;
    wire N__5183;
    wire N__5178;
    wire N__5171;
    wire N__5170;
    wire N__5169;
    wire N__5164;
    wire N__5161;
    wire N__5156;
    wire N__5153;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5135;
    wire N__5130;
    wire N__5129;
    wire N__5126;
    wire N__5121;
    wire N__5114;
    wire N__5107;
    wire N__5104;
    wire N__5093;
    wire N__5090;
    wire N__5087;
    wire N__5086;
    wire N__5085;
    wire N__5078;
    wire N__5077;
    wire N__5074;
    wire N__5071;
    wire N__5066;
    wire N__5063;
    wire N__5060;
    wire N__5057;
    wire N__5054;
    wire N__5053;
    wire N__5050;
    wire N__5047;
    wire N__5042;
    wire N__5041;
    wire N__5038;
    wire N__5037;
    wire N__5036;
    wire N__5035;
    wire N__5032;
    wire N__5029;
    wire N__5022;
    wire N__5019;
    wire N__5016;
    wire N__5013;
    wire N__5006;
    wire N__5003;
    wire N__5000;
    wire N__4997;
    wire N__4996;
    wire N__4993;
    wire N__4992;
    wire N__4989;
    wire N__4986;
    wire N__4983;
    wire N__4980;
    wire N__4975;
    wire N__4972;
    wire N__4969;
    wire N__4966;
    wire N__4963;
    wire N__4958;
    wire N__4955;
    wire N__4952;
    wire N__4949;
    wire N__4946;
    wire N__4943;
    wire N__4940;
    wire N__4937;
    wire N__4934;
    wire N__4931;
    wire N__4928;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4916;
    wire N__4913;
    wire N__4910;
    wire N__4907;
    wire N__4904;
    wire N__4901;
    wire N__4898;
    wire N__4895;
    wire N__4892;
    wire N__4891;
    wire N__4888;
    wire N__4885;
    wire N__4882;
    wire N__4879;
    wire N__4876;
    wire N__4873;
    wire N__4868;
    wire N__4865;
    wire N__4862;
    wire N__4859;
    wire N__4856;
    wire N__4853;
    wire N__4850;
    wire N__4847;
    wire N__4844;
    wire N__4841;
    wire N__4838;
    wire N__4835;
    wire N__4832;
    wire N__4831;
    wire N__4828;
    wire N__4825;
    wire N__4820;
    wire N__4817;
    wire N__4814;
    wire N__4811;
    wire N__4810;
    wire N__4809;
    wire N__4806;
    wire N__4801;
    wire N__4796;
    wire N__4795;
    wire N__4790;
    wire N__4787;
    wire N__4784;
    wire N__4781;
    wire N__4780;
    wire N__4777;
    wire N__4776;
    wire N__4773;
    wire N__4770;
    wire N__4767;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4748;
    wire N__4745;
    wire N__4742;
    wire N__4739;
    wire N__4736;
    wire N__4733;
    wire N__4730;
    wire N__4729;
    wire N__4724;
    wire N__4723;
    wire N__4722;
    wire N__4721;
    wire N__4720;
    wire N__4719;
    wire N__4718;
    wire N__4715;
    wire N__4708;
    wire N__4701;
    wire N__4694;
    wire N__4691;
    wire N__4688;
    wire N__4687;
    wire N__4686;
    wire N__4683;
    wire N__4680;
    wire N__4677;
    wire N__4674;
    wire N__4667;
    wire N__4664;
    wire N__4661;
    wire N__4660;
    wire N__4657;
    wire N__4656;
    wire N__4653;
    wire N__4650;
    wire N__4647;
    wire N__4644;
    wire N__4637;
    wire N__4634;
    wire N__4631;
    wire N__4628;
    wire N__4625;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4613;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4601;
    wire N__4598;
    wire N__4595;
    wire N__4592;
    wire N__4591;
    wire N__4588;
    wire N__4585;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4565;
    wire N__4562;
    wire N__4561;
    wire N__4558;
    wire N__4557;
    wire N__4554;
    wire N__4551;
    wire N__4548;
    wire N__4541;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4523;
    wire N__4520;
    wire N__4519;
    wire N__4516;
    wire N__4513;
    wire N__4508;
    wire N__4505;
    wire N__4504;
    wire N__4501;
    wire N__4498;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4486;
    wire N__4483;
    wire N__4480;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4463;
    wire N__4460;
    wire N__4457;
    wire N__4456;
    wire N__4453;
    wire N__4450;
    wire N__4445;
    wire N__4442;
    wire N__4441;
    wire N__4438;
    wire N__4435;
    wire N__4432;
    wire N__4429;
    wire N__4424;
    wire N__4421;
    wire N__4418;
    wire N__4415;
    wire N__4412;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4400;
    wire N__4397;
    wire N__4394;
    wire N__4391;
    wire N__4388;
    wire N__4387;
    wire N__4386;
    wire N__4383;
    wire N__4378;
    wire N__4375;
    wire N__4370;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4348;
    wire N__4345;
    wire N__4342;
    wire N__4337;
    wire N__4334;
    wire N__4331;
    wire N__4330;
    wire N__4327;
    wire N__4324;
    wire N__4321;
    wire N__4316;
    wire N__4315;
    wire N__4314;
    wire N__4311;
    wire N__4308;
    wire N__4305;
    wire N__4300;
    wire N__4297;
    wire N__4294;
    wire N__4291;
    wire N__4288;
    wire N__4285;
    wire N__4282;
    wire N__4279;
    wire N__4276;
    wire N__4271;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4258;
    wire N__4255;
    wire N__4250;
    wire N__4249;
    wire N__4248;
    wire N__4247;
    wire N__4246;
    wire N__4245;
    wire N__4244;
    wire N__4243;
    wire N__4240;
    wire N__4223;
    wire N__4220;
    wire N__4217;
    wire N__4216;
    wire N__4213;
    wire N__4210;
    wire N__4205;
    wire N__4204;
    wire N__4201;
    wire N__4198;
    wire N__4195;
    wire N__4192;
    wire N__4189;
    wire N__4186;
    wire N__4183;
    wire N__4180;
    wire N__4177;
    wire N__4174;
    wire N__4169;
    wire N__4166;
    wire N__4163;
    wire N__4160;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4148;
    wire N__4145;
    wire N__4142;
    wire N__4139;
    wire N__4136;
    wire N__4133;
    wire N__4130;
    wire N__4127;
    wire N__4124;
    wire N__4121;
    wire N__4118;
    wire N__4115;
    wire N__4112;
    wire N__4109;
    wire N__4106;
    wire N__4103;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4088;
    wire N__4085;
    wire N__4082;
    wire N__4079;
    wire N__4076;
    wire N__4073;
    wire N__4070;
    wire N__4067;
    wire N__4064;
    wire N__4061;
    wire N__4058;
    wire N__4055;
    wire N__4052;
    wire N__4049;
    wire N__4046;
    wire N__4043;
    wire N__4040;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire CLK80_PLL_i_i;
    wire \U712_CHIP_RAM.N_448_cascade_ ;
    wire \U712_CHIP_RAM.N_459_cascade_ ;
    wire \U712_CHIP_RAM.N_308_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_416_cascade_ ;
    wire \U712_CHIP_RAM.N_448 ;
    wire \U712_CHIP_RAM.N_261_cascade_ ;
    wire \U712_CHIP_RAM.N_404_cascade_ ;
    wire \U712_CHIP_RAM.N_413_cascade_ ;
    wire \U712_CHIP_RAM.N_414 ;
    wire \U712_CHIP_RAM.N_415_cascade_ ;
    wire \U712_CHIP_RAM.N_373_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_0 ;
    wire \U712_CHIP_RAM.N_373 ;
    wire N_48_i;
    wire RAMSPACEn_c;
    wire \U712_CHIP_RAM.N_355_cascade_ ;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0 ;
    wire TACK_OUTn;
    wire DBR_SYNCZ0Z_0;
    wire DBR_SYNCZ0Z_1;
    wire CLK40_PLL;
    wire \U712_BYTE_ENABLE.N_90 ;
    wire CLK40_PLL_g;
    wire CLK40_PLL_iso_i;
    wire LATCH_RAM;
    wire LATCH_CLK_0_i;
    wire \U712_CHIP_RAM.N_296_cascade_ ;
    wire \U712_CHIP_RAM.N_296 ;
    wire \U712_CHIP_RAM.N_63 ;
    wire bfn_8_8_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire BANK0_c;
    wire \U712_CHIP_RAM.N_404 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_ ;
    wire A_c_20;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_ ;
    wire \U712_CHIP_RAM.N_362 ;
    wire \U712_CHIP_RAM.N_470 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_1_0_cascade_ ;
    wire \U712_CHIP_RAM.N_344 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_i_i_a3_0_0 ;
    wire \U712_CHIP_RAM.N_344_cascade_ ;
    wire \U712_CHIP_RAM.N_267 ;
    wire \U712_CHIP_RAM.N_333 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_0_cascade_ ;
    wire \U712_CHIP_RAM.N_416 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0_a2_0_a3_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0_a2_0_a3_0 ;
    wire \U712_CHIP_RAM.N_45 ;
    wire \U712_CHIP_RAM.N_61_cascade_ ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.N_263 ;
    wire \U712_CHIP_RAM.N_271 ;
    wire \U712_CHIP_RAM.N_341_cascade_ ;
    wire \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_i_0_2 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_START_RNOZ0Z_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_2 ;
    wire \U712_CYCLE_TERM.TACK_STATE_r_sx_1 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire \U712_CYCLE_TERM.N_286_i_0_0_cascade_ ;
    wire \U712_CYCLE_TERM.N_286_i_0_en_cascade_ ;
    wire RESETn_c_i;
    wire CPU_TACK;
    wire \U712_CYCLE_TERM.N_286_i_0_en_0 ;
    wire DBRn_c;
    wire \U712_REG_SM.DBR_SYNCZ0Z_0 ;
    wire \INVU712_REG_SM.DBR_SYNC_1C_net ;
    wire TACK_EN_i_ess;
    wire N_977_i;
    wire VBENn_c;
    wire CONSTANT_ONE_NET;
    wire A_c_6;
    wire A_c_13;
    wire A_c_12;
    wire A_c_5;
    wire A_c_15;
    wire A_c_8;
    wire \U712_CHIP_RAM.N_261 ;
    wire A_c_11;
    wire A_c_4;
    wire \U712_CHIP_RAM.N_312 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_63_i_a2_0_i_0 ;
    wire \U712_CHIP_RAM.N_314 ;
    wire \U712_CHIP_RAM.N_459 ;
    wire \U712_CHIP_RAM.N_449 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i_1_cascade_ ;
    wire RESETn_c;
    wire \U712_CHIP_RAM.N_421 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_0_2 ;
    wire \U712_CHIP_RAM.N_421_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire \U712_CHIP_RAM.DMA_AZ0Z20 ;
    wire \INVU712_CHIP_RAM.DMA_A20C_net ;
    wire \U712_CHIP_RAM.N_18 ;
    wire \U712_CHIP_RAM.N_18_0 ;
    wire \U712_CHIP_RAM.N_113 ;
    wire \U712_CHIP_RAM.N_413 ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa ;
    wire \U712_CHIP_RAM.N_342 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0 ;
    wire AWEn_c;
    wire DBDIR_c;
    wire DBRn_c_i;
    wire DBRn_c_i_0;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_1_0_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_5 ;
    wire LATCH_REG;
    wire REG_CPU_CYCLE;
    wire \INVU712_REG_SM.STATE_COUNTER_5C_net ;
    wire \U712_REG_SM.STATE_COUNTERc_0_cascade_ ;
    wire \U712_REG_SM.REG_CPU_CYCLE_e_1 ;
    wire A_c_3;
    wire A_c_10;
    wire A_c_16;
    wire A_c_18;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ;
    wire \U712_CHIP_RAM.N_411_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_1_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_o3_0_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_1_0_cascade_ ;
    wire \U712_CHIP_RAM.N_294 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.N_316_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_101_i_a2_0_i_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_0 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER15 ;
    wire \U712_CHIP_RAM.N_109_i ;
    wire \U712_REG_SM.STATE_COUNTERc_0 ;
    wire \U712_REG_SM.un15_0_i_0_0 ;
    wire \U712_REG_SM.N_297 ;
    wire REG_TACK;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_6 ;
    wire REGENn_c;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_4 ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_3 ;
    wire \INVU712_REG_SM.REG_CYCLEC_net ;
    wire \U712_REG_SM.DBR_SYNCZ0Z_1 ;
    wire \INVU712_REG_SM.STATE_COUNTER_2C_net ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ;
    wire A_c_14;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ;
    wire DBENn_c;
    wire DMA_CYCLE;
    wire \U712_CHIP_RAM.REFRESH5lt7 ;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0Z0Z_0 ;
    wire N_49_i;
    wire \U712_BYTE_ENABLE.N_92 ;
    wire N_315;
    wire \U712_REG_SM.N_278_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_7 ;
    wire \U712_REG_SM.N_272 ;
    wire \U712_REG_SM.N_309 ;
    wire \U712_REG_SM.N_272_cascade_ ;
    wire C3_c;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire C1_c;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_REG_SM.LDSn_7_iv_i_0_0 ;
    wire \U712_REG_SM.N_278 ;
    wire ASn_c;
    wire \INVU712_REG_SM.C3_SYNC_0C_net ;
    wire WRITE_CYCLE;
    wire N_259;
    wire LDSn_c;
    wire \U712_REG_SM.N_467_cascade_ ;
    wire \U712_REG_SM.N_371 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ;
    wire CMA_c_5;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ;
    wire A_c_7;
    wire \U712_CHIP_RAM.N_329 ;
    wire A_c_2;
    wire A_c_9;
    wire \U712_CHIP_RAM.REFRESH5lto7_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire bfn_12_10_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire C1_c_g;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire \U712_REG_SM.UDSn_7_iv_i_0_0 ;
    wire \U712_REG_SM.C1_SYNC_RNI5ITS1Z0Z_1 ;
    wire \U712_REG_SM.LATCH_REG_0_sqmuxa ;
    wire \INVU712_REG_SM.UDSnC_net ;
    wire RAMENn_c;
    wire TSn_c;
    wire \U712_REG_SM.CYCLE_RUNZ0 ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_1 ;
    wire RnW_c;
    wire REG_WRITE_CYCLE;
    wire \INVU712_REG_SM.REG_CYCLE_STARTC_net ;
    wire \U712_CHIP_RAM.un1_CMA28_0_i_cascade_ ;
    wire CMA_c_0;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ;
    wire CMA_c_2;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ;
    wire CMA_c_7;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire DRA_c_1;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_0 ;
    wire \U712_REG_SM.N_369 ;
    wire UDSn_c;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_2 ;
    wire \U712_REG_SM.N_465 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.N_288 ;
    wire CASn_c;
    wire WEn_c;
    wire RASn_c;
    wire CRCSn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire CMA_c_10;
    wire A_c_17;
    wire CMA_c_8;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire CMA_c_3;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.CMA_5_sn_N_5_mux ;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ;
    wire CMA_c_4;
    wire A_c_19;
    wire \U712_CHIP_RAM.CMA_5_0_8 ;
    wire CMA_c_9;
    wire CLK80_PLL;
    wire \U712_CHIP_RAM.un1_CMA28_0_i_0 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire RAS0n_c;
    wire DRA_c_9;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire DRA_c_6;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire N_50_i;
    wire CPU_CYCLE;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0Z0Z_0 ;
    wire \U712_BYTE_ENABLE.N_91_cascade_ ;
    wire N_51_i;
    wire \U712_BYTE_ENABLE.N_89 ;
    wire N_90_i;
    wire N_92_i;
    wire N_91_i;
    wire SIZ_c_1;
    wire A_c_1;
    wire SIZ_c_0;
    wire A_c_0;
    wire N_89_i;
    wire DRA_c_3;
    wire DRA_c_2;
    wire AGNUS_REV_c;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire C3_c_g;
    wire DBRn_c_i_0_g;
    wire RESETn_c_i_g;
    wire REG_CYCLE;
    wire CASUn_c;
    wire CASLn_c;
    wire DRDENn_c;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL),
            .REFERENCECLK(N__4061),
            .RESETB(N__4901),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__11850),
            .DIN(N__11849),
            .DOUT(N__11848),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__11850),
            .PADOUT(N__11849),
            .PADIN(N__11848),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7052),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__11841),
            .DIN(N__11840),
            .DOUT(N__11839),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__11841),
            .PADOUT(N__11840),
            .PADIN(N__11839),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__11832),
            .DIN(N__11831),
            .DOUT(N__11830),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__11832),
            .PADOUT(N__11831),
            .PADIN(N__11830),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8198),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__11823),
            .DIN(N__11822),
            .DOUT(N__11821),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__11823),
            .PADOUT(N__11822),
            .PADIN(N__11821),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7241),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__11814),
            .DIN(N__11813),
            .DOUT(N__11812),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__11814),
            .PADOUT(N__11813),
            .PADIN(N__11812),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__11805),
            .DIN(N__11804),
            .DOUT(N__11803),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__11805),
            .PADOUT(N__11804),
            .PADIN(N__11803),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__11796),
            .DIN(N__11795),
            .DOUT(N__11794),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__11796),
            .PADOUT(N__11795),
            .PADIN(N__11794),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__11787),
            .DIN(N__11786),
            .DOUT(N__11785),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__11787),
            .PADOUT(N__11786),
            .PADIN(N__11785),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__11778),
            .DIN(N__11777),
            .DOUT(N__11776),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__11778),
            .PADOUT(N__11777),
            .PADIN(N__11776),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__11769),
            .DIN(N__11768),
            .DOUT(N__11767),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__11769),
            .PADOUT(N__11768),
            .PADIN(N__11767),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__11760),
            .DIN(N__11759),
            .DOUT(N__11758),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__11760),
            .PADOUT(N__11759),
            .PADIN(N__11758),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8171),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__11751),
            .DIN(N__11750),
            .DOUT(N__11749),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__11751),
            .PADOUT(N__11750),
            .PADIN(N__11749),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10436),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__11742),
            .DIN(N__11741),
            .DOUT(N__11740),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__11742),
            .PADOUT(N__11741),
            .PADIN(N__11740),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMENn_obuf_iopad (
            .OE(N__11733),
            .DIN(N__11732),
            .DOUT(N__11731),
            .PACKAGEPIN(RAMENn));
    defparam RAMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMENn_obuf_preio (
            .PADOEN(N__11733),
            .PADOUT(N__11732),
            .PADIN(N__11731),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8051),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__11724),
            .DIN(N__11723),
            .DOUT(N__11722),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__11724),
            .PADOUT(N__11723),
            .PADIN(N__11722),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__11715),
            .DIN(N__11714),
            .DOUT(N__11713),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__11715),
            .PADOUT(N__11714),
            .PADIN(N__11713),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__11706),
            .DIN(N__11705),
            .DOUT(N__11704),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__11706),
            .PADOUT(N__11705),
            .PADIN(N__11704),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4919),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__11697),
            .DIN(N__11696),
            .DOUT(N__11695),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__11697),
            .PADOUT(N__11696),
            .PADIN(N__11695),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__11688),
            .DIN(N__11687),
            .DOUT(N__11686),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__11688),
            .PADOUT(N__11687),
            .PADIN(N__11686),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__11679),
            .DIN(N__11678),
            .DOUT(N__11677),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__11679),
            .PADOUT(N__11678),
            .PADIN(N__11677),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7841),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__11670),
            .DIN(N__11669),
            .DOUT(N__11668),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__11670),
            .PADOUT(N__11669),
            .PADIN(N__11668),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__11661),
            .DIN(N__11660),
            .DOUT(N__11659),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__11661),
            .PADOUT(N__11660),
            .PADIN(N__11659),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9209),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__11652),
            .DIN(N__11651),
            .DOUT(N__11650),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__11652),
            .PADOUT(N__11651),
            .PADIN(N__11650),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__11643),
            .DIN(N__11642),
            .DOUT(N__11641),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__11643),
            .PADOUT(N__11642),
            .PADIN(N__11641),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10469),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__11634),
            .DIN(N__11633),
            .DOUT(N__11632),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__11634),
            .PADOUT(N__11633),
            .PADIN(N__11632),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__11625),
            .DIN(N__11624),
            .DOUT(N__11623),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__11625),
            .PADOUT(N__11624),
            .PADIN(N__11623),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__11616),
            .DIN(N__11615),
            .DOUT(N__11614),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__11616),
            .PADOUT(N__11615),
            .PADIN(N__11614),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__11607),
            .DIN(N__11606),
            .DOUT(N__11605),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__11607),
            .PADOUT(N__11606),
            .PADIN(N__11605),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__11598),
            .DIN(N__11597),
            .DOUT(N__11596),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__11598),
            .PADOUT(N__11597),
            .PADIN(N__11596),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_EN_obuf_iopad (
            .OE(N__11589),
            .DIN(N__11588),
            .DOUT(N__11587),
            .PACKAGEPIN(DMA_LATCH_EN));
    defparam DMA_LATCH_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_EN_obuf_preio (
            .PADOEN(N__11589),
            .PADOUT(N__11588),
            .PADIN(N__11587),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7370),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__11580),
            .DIN(N__11579),
            .DOUT(N__11578),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__11580),
            .PADOUT(N__11579),
            .PADIN(N__11578),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__11571),
            .DIN(N__11570),
            .DOUT(N__11569),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__11571),
            .PADOUT(N__11570),
            .PADIN(N__11569),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__11562),
            .DIN(N__11561),
            .DOUT(N__11560),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__11562),
            .PADOUT(N__11561),
            .PADIN(N__11560),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__11553),
            .DIN(N__11552),
            .DOUT(N__11551),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__11553),
            .PADOUT(N__11552),
            .PADIN(N__11551),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__11544),
            .DIN(N__11543),
            .DOUT(N__11542),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__11544),
            .PADOUT(N__11543),
            .PADIN(N__11542),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__11535),
            .DIN(N__11534),
            .DOUT(N__11533),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__11535),
            .PADOUT(N__11534),
            .PADIN(N__11533),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9227),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__11526),
            .DIN(N__11525),
            .DOUT(N__11524),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__11526),
            .PADOUT(N__11525),
            .PADIN(N__11524),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4475),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__11517),
            .DIN(N__11516),
            .DOUT(N__11515),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__11517),
            .PADOUT(N__11516),
            .PADIN(N__11515),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4216),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__11508),
            .DIN(N__11507),
            .DOUT(N__11506),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__11508),
            .PADOUT(N__11507),
            .PADIN(N__11506),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4091),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__11499),
            .DIN(N__11498),
            .DOUT(N__11497),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__11499),
            .PADOUT(N__11498),
            .PADIN(N__11497),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__11490),
            .DIN(N__11489),
            .DOUT(N__11488),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__11490),
            .PADOUT(N__11489),
            .PADIN(N__11488),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7457),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__11481),
            .DIN(N__11480),
            .DOUT(N__11479),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__11481),
            .PADOUT(N__11480),
            .PADIN(N__11479),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8822),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__11472),
            .DIN(N__11471),
            .DOUT(N__11470),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__11472),
            .PADOUT(N__11471),
            .PADIN(N__11470),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__11463),
            .DIN(N__11462),
            .DOUT(N__11461),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__11463),
            .PADOUT(N__11462),
            .PADIN(N__11461),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__11454),
            .DIN(N__11453),
            .DOUT(N__11452),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__11454),
            .PADOUT(N__11453),
            .PADIN(N__11452),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__11445),
            .DIN(N__11444),
            .DOUT(N__11443),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__11445),
            .PADOUT(N__11444),
            .PADIN(N__11443),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__11436),
            .DIN(N__11435),
            .DOUT(N__11434),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__11436),
            .PADOUT(N__11435),
            .PADIN(N__11434),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8885),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__11427),
            .DIN(N__11426),
            .DOUT(N__11425),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__11427),
            .PADOUT(N__11426),
            .PADIN(N__11425),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__11418),
            .DIN(N__11417),
            .DOUT(N__11416),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__11418),
            .PADOUT(N__11417),
            .PADIN(N__11416),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4204),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__11409),
            .DIN(N__11408),
            .DOUT(N__11407),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__11409),
            .PADOUT(N__11408),
            .PADIN(N__11407),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8687),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__11400),
            .DIN(N__11399),
            .DOUT(N__11398),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__11400),
            .PADOUT(N__11399),
            .PADIN(N__11398),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10715),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__11391),
            .DIN(N__11390),
            .DOUT(N__11389),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__11391),
            .PADOUT(N__11390),
            .PADIN(N__11389),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4142),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__11382),
            .DIN(N__11381),
            .DOUT(N__11380),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__11382),
            .PADOUT(N__11381),
            .PADIN(N__11380),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8615),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__11373),
            .DIN(N__11372),
            .DOUT(N__11371),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__11373),
            .PADOUT(N__11372),
            .PADIN(N__11371),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6818),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__11364),
            .DIN(N__11363),
            .DOUT(N__11362),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__11364),
            .PADOUT(N__11363),
            .PADIN(N__11362),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__11355),
            .DIN(N__11354),
            .DOUT(N__11353),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__11355),
            .PADOUT(N__11354),
            .PADIN(N__11353),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__11346),
            .DIN(N__11345),
            .DOUT(N__11344),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__11346),
            .PADOUT(N__11345),
            .PADIN(N__11344),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6929),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__11337),
            .DIN(N__11336),
            .DOUT(N__11335),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__11337),
            .PADOUT(N__11336),
            .PADIN(N__11335),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9245),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__11328),
            .DIN(N__11327),
            .DOUT(N__11326),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__11328),
            .PADOUT(N__11327),
            .PADIN(N__11326),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5492),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__11319),
            .DIN(N__11318),
            .DOUT(N__11317),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__11319),
            .PADOUT(N__11318),
            .PADIN(N__11317),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9269),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__11310),
            .DIN(N__11309),
            .DOUT(N__11308),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__11310),
            .PADOUT(N__11309),
            .PADIN(N__11308),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__11301),
            .DIN(N__11300),
            .DOUT(N__11299),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__11301),
            .PADOUT(N__11300),
            .PADIN(N__11299),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__11292),
            .DIN(N__11291),
            .DOUT(N__11290),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__11292),
            .PADOUT(N__11291),
            .PADIN(N__11290),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__11283),
            .DIN(N__11282),
            .DOUT(N__11281),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__11283),
            .PADOUT(N__11282),
            .PADIN(N__11281),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__11274),
            .DIN(N__11273),
            .DOUT(N__11272),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__11274),
            .PADOUT(N__11273),
            .PADIN(N__11272),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7298),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__11265),
            .DIN(N__11264),
            .DOUT(N__11263),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__11265),
            .PADOUT(N__11264),
            .PADIN(N__11263),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10454),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__11256),
            .DIN(N__11255),
            .DOUT(N__11254),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__11256),
            .PADOUT(N__11255),
            .PADIN(N__11254),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__11247),
            .DIN(N__11246),
            .DOUT(N__11245),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__11247),
            .PADOUT(N__11246),
            .PADIN(N__11245),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10496),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__11238),
            .DIN(N__11237),
            .DOUT(N__11236),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__11238),
            .PADOUT(N__11237),
            .PADIN(N__11236),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4940),
            .DIN0(),
            .DOUT0(N__4364),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__11229),
            .DIN(N__11228),
            .DOUT(N__11227),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__11229),
            .PADOUT(N__11228),
            .PADIN(N__11227),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7817),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__11220),
            .DIN(N__11219),
            .DOUT(N__11218),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__11220),
            .PADOUT(N__11219),
            .PADIN(N__11218),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__11211),
            .DIN(N__11210),
            .DOUT(N__11209),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__11211),
            .PADOUT(N__11210),
            .PADIN(N__11209),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__11202),
            .DIN(N__11201),
            .DOUT(N__11200),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__11202),
            .PADOUT(N__11201),
            .PADIN(N__11200),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8852),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__11193),
            .DIN(N__11192),
            .DOUT(N__11191),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__11193),
            .PADOUT(N__11192),
            .PADIN(N__11191),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__11184),
            .DIN(N__11183),
            .DOUT(N__11182),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__11184),
            .PADOUT(N__11183),
            .PADIN(N__11182),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__11175),
            .DIN(N__11174),
            .DOUT(N__11173),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__11175),
            .PADOUT(N__11174),
            .PADIN(N__11173),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__11166),
            .DIN(N__11165),
            .DOUT(N__11164),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__11166),
            .PADOUT(N__11165),
            .PADIN(N__11164),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__11157),
            .DIN(N__11156),
            .DOUT(N__11155),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__11157),
            .PADOUT(N__11156),
            .PADIN(N__11155),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7277),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__11148),
            .DIN(N__11147),
            .DOUT(N__11146),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__11148),
            .PADOUT(N__11147),
            .PADIN(N__11146),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8441),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__11139),
            .DIN(N__11138),
            .DOUT(N__11137),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__11139),
            .PADOUT(N__11138),
            .PADIN(N__11137),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10094),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__11130),
            .DIN(N__11129),
            .DOUT(N__11128),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__11130),
            .PADOUT(N__11129),
            .PADIN(N__11128),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5582),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__11121),
            .DIN(N__11120),
            .DOUT(N__11119),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__11121),
            .PADOUT(N__11120),
            .PADIN(N__11119),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__11112),
            .DIN(N__11111),
            .DOUT(N__11110),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__11112),
            .PADOUT(N__11111),
            .PADIN(N__11110),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__11103),
            .DIN(N__11102),
            .DOUT(N__11101),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__11103),
            .PADOUT(N__11102),
            .PADIN(N__11101),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8801),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__11094),
            .DIN(N__11093),
            .DOUT(N__11092),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__11094),
            .PADOUT(N__11093),
            .PADIN(N__11092),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__11085),
            .DIN(N__11084),
            .DOUT(N__11083),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__11085),
            .PADOUT(N__11084),
            .PADIN(N__11083),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__11076),
            .DIN(N__11075),
            .DOUT(N__11074),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__11076),
            .PADOUT(N__11075),
            .PADIN(N__11074),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4424),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__11067),
            .DIN(N__11066),
            .DOUT(N__11065),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__11067),
            .PADOUT(N__11066),
            .PADIN(N__11065),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7352),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__11058),
            .DIN(N__11057),
            .DOUT(N__11056),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__11058),
            .PADOUT(N__11057),
            .PADIN(N__11056),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4217),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__11049),
            .DIN(N__11048),
            .DOUT(N__11047),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__11049),
            .PADOUT(N__11048),
            .PADIN(N__11047),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2684 (
            .O(N__11030),
            .I(N__11024));
    InMux I__2683 (
            .O(N__11029),
            .I(N__11021));
    InMux I__2682 (
            .O(N__11028),
            .I(N__11018));
    InMux I__2681 (
            .O(N__11027),
            .I(N__11015));
    LocalMux I__2680 (
            .O(N__11024),
            .I(N__11009));
    LocalMux I__2679 (
            .O(N__11021),
            .I(N__11004));
    LocalMux I__2678 (
            .O(N__11018),
            .I(N__10996));
    LocalMux I__2677 (
            .O(N__11015),
            .I(N__10984));
    SRMux I__2676 (
            .O(N__11014),
            .I(N__10901));
    SRMux I__2675 (
            .O(N__11013),
            .I(N__10901));
    SRMux I__2674 (
            .O(N__11012),
            .I(N__10901));
    Glb2LocalMux I__2673 (
            .O(N__11009),
            .I(N__10901));
    SRMux I__2672 (
            .O(N__11008),
            .I(N__10901));
    SRMux I__2671 (
            .O(N__11007),
            .I(N__10901));
    Glb2LocalMux I__2670 (
            .O(N__11004),
            .I(N__10901));
    SRMux I__2669 (
            .O(N__11003),
            .I(N__10901));
    SRMux I__2668 (
            .O(N__11002),
            .I(N__10901));
    SRMux I__2667 (
            .O(N__11001),
            .I(N__10901));
    SRMux I__2666 (
            .O(N__11000),
            .I(N__10901));
    SRMux I__2665 (
            .O(N__10999),
            .I(N__10901));
    Glb2LocalMux I__2664 (
            .O(N__10996),
            .I(N__10901));
    SRMux I__2663 (
            .O(N__10995),
            .I(N__10901));
    SRMux I__2662 (
            .O(N__10994),
            .I(N__10901));
    SRMux I__2661 (
            .O(N__10993),
            .I(N__10901));
    SRMux I__2660 (
            .O(N__10992),
            .I(N__10901));
    SRMux I__2659 (
            .O(N__10991),
            .I(N__10901));
    SRMux I__2658 (
            .O(N__10990),
            .I(N__10901));
    SRMux I__2657 (
            .O(N__10989),
            .I(N__10901));
    SRMux I__2656 (
            .O(N__10988),
            .I(N__10901));
    SRMux I__2655 (
            .O(N__10987),
            .I(N__10901));
    Glb2LocalMux I__2654 (
            .O(N__10984),
            .I(N__10901));
    SRMux I__2653 (
            .O(N__10983),
            .I(N__10901));
    SRMux I__2652 (
            .O(N__10982),
            .I(N__10901));
    SRMux I__2651 (
            .O(N__10981),
            .I(N__10901));
    SRMux I__2650 (
            .O(N__10980),
            .I(N__10901));
    SRMux I__2649 (
            .O(N__10979),
            .I(N__10901));
    SRMux I__2648 (
            .O(N__10978),
            .I(N__10901));
    SRMux I__2647 (
            .O(N__10977),
            .I(N__10901));
    SRMux I__2646 (
            .O(N__10976),
            .I(N__10901));
    SRMux I__2645 (
            .O(N__10975),
            .I(N__10901));
    SRMux I__2644 (
            .O(N__10974),
            .I(N__10901));
    SRMux I__2643 (
            .O(N__10973),
            .I(N__10901));
    SRMux I__2642 (
            .O(N__10972),
            .I(N__10901));
    GlobalMux I__2641 (
            .O(N__10901),
            .I(N__10898));
    gio2CtrlBuf I__2640 (
            .O(N__10898),
            .I(RESETn_c_i_g));
    InMux I__2639 (
            .O(N__10895),
            .I(N__10892));
    LocalMux I__2638 (
            .O(N__10892),
            .I(N__10889));
    Span4Mux_h I__2637 (
            .O(N__10889),
            .I(N__10886));
    Span4Mux_h I__2636 (
            .O(N__10886),
            .I(N__10883));
    Span4Mux_h I__2635 (
            .O(N__10883),
            .I(N__10880));
    Span4Mux_v I__2634 (
            .O(N__10880),
            .I(N__10876));
    InMux I__2633 (
            .O(N__10879),
            .I(N__10873));
    Odrv4 I__2632 (
            .O(N__10876),
            .I(REG_CYCLE));
    LocalMux I__2631 (
            .O(N__10873),
            .I(REG_CYCLE));
    InMux I__2630 (
            .O(N__10868),
            .I(N__10865));
    LocalMux I__2629 (
            .O(N__10865),
            .I(N__10861));
    InMux I__2628 (
            .O(N__10864),
            .I(N__10858));
    Span4Mux_v I__2627 (
            .O(N__10861),
            .I(N__10854));
    LocalMux I__2626 (
            .O(N__10858),
            .I(N__10851));
    InMux I__2625 (
            .O(N__10857),
            .I(N__10848));
    Span4Mux_h I__2624 (
            .O(N__10854),
            .I(N__10841));
    Span4Mux_v I__2623 (
            .O(N__10851),
            .I(N__10841));
    LocalMux I__2622 (
            .O(N__10848),
            .I(N__10841));
    Span4Mux_v I__2621 (
            .O(N__10841),
            .I(N__10838));
    Span4Mux_h I__2620 (
            .O(N__10838),
            .I(N__10833));
    InMux I__2619 (
            .O(N__10837),
            .I(N__10829));
    InMux I__2618 (
            .O(N__10836),
            .I(N__10826));
    Span4Mux_h I__2617 (
            .O(N__10833),
            .I(N__10823));
    InMux I__2616 (
            .O(N__10832),
            .I(N__10820));
    LocalMux I__2615 (
            .O(N__10829),
            .I(N__10817));
    LocalMux I__2614 (
            .O(N__10826),
            .I(N__10814));
    Span4Mux_h I__2613 (
            .O(N__10823),
            .I(N__10809));
    LocalMux I__2612 (
            .O(N__10820),
            .I(N__10809));
    Span12Mux_h I__2611 (
            .O(N__10817),
            .I(N__10806));
    Span12Mux_v I__2610 (
            .O(N__10814),
            .I(N__10803));
    Span4Mux_h I__2609 (
            .O(N__10809),
            .I(N__10800));
    Span12Mux_v I__2608 (
            .O(N__10806),
            .I(N__10797));
    Span12Mux_h I__2607 (
            .O(N__10803),
            .I(N__10794));
    Span4Mux_v I__2606 (
            .O(N__10800),
            .I(N__10791));
    Odrv12 I__2605 (
            .O(N__10797),
            .I(CASUn_c));
    Odrv12 I__2604 (
            .O(N__10794),
            .I(CASUn_c));
    Odrv4 I__2603 (
            .O(N__10791),
            .I(CASUn_c));
    InMux I__2602 (
            .O(N__10784),
            .I(N__10779));
    InMux I__2601 (
            .O(N__10783),
            .I(N__10776));
    CascadeMux I__2600 (
            .O(N__10782),
            .I(N__10772));
    LocalMux I__2599 (
            .O(N__10779),
            .I(N__10767));
    LocalMux I__2598 (
            .O(N__10776),
            .I(N__10767));
    InMux I__2597 (
            .O(N__10775),
            .I(N__10764));
    InMux I__2596 (
            .O(N__10772),
            .I(N__10760));
    Span4Mux_v I__2595 (
            .O(N__10767),
            .I(N__10755));
    LocalMux I__2594 (
            .O(N__10764),
            .I(N__10755));
    InMux I__2593 (
            .O(N__10763),
            .I(N__10752));
    LocalMux I__2592 (
            .O(N__10760),
            .I(N__10749));
    Span4Mux_h I__2591 (
            .O(N__10755),
            .I(N__10744));
    LocalMux I__2590 (
            .O(N__10752),
            .I(N__10744));
    Span4Mux_v I__2589 (
            .O(N__10749),
            .I(N__10741));
    Sp12to4 I__2588 (
            .O(N__10744),
            .I(N__10737));
    Sp12to4 I__2587 (
            .O(N__10741),
            .I(N__10734));
    InMux I__2586 (
            .O(N__10740),
            .I(N__10731));
    Span12Mux_v I__2585 (
            .O(N__10737),
            .I(N__10728));
    Span12Mux_h I__2584 (
            .O(N__10734),
            .I(N__10723));
    LocalMux I__2583 (
            .O(N__10731),
            .I(N__10723));
    Span12Mux_h I__2582 (
            .O(N__10728),
            .I(N__10718));
    Span12Mux_v I__2581 (
            .O(N__10723),
            .I(N__10718));
    Odrv12 I__2580 (
            .O(N__10718),
            .I(CASLn_c));
    IoInMux I__2579 (
            .O(N__10715),
            .I(N__10712));
    LocalMux I__2578 (
            .O(N__10712),
            .I(N__10709));
    Span4Mux_s3_v I__2577 (
            .O(N__10709),
            .I(N__10706));
    Span4Mux_v I__2576 (
            .O(N__10706),
            .I(N__10703));
    Sp12to4 I__2575 (
            .O(N__10703),
            .I(N__10700));
    Odrv12 I__2574 (
            .O(N__10700),
            .I(DRDENn_c));
    CascadeMux I__2573 (
            .O(N__10697),
            .I(N__10694));
    InMux I__2572 (
            .O(N__10694),
            .I(N__10687));
    CascadeMux I__2571 (
            .O(N__10693),
            .I(N__10683));
    CascadeMux I__2570 (
            .O(N__10692),
            .I(N__10680));
    CascadeMux I__2569 (
            .O(N__10691),
            .I(N__10675));
    InMux I__2568 (
            .O(N__10690),
            .I(N__10667));
    LocalMux I__2567 (
            .O(N__10687),
            .I(N__10664));
    InMux I__2566 (
            .O(N__10686),
            .I(N__10661));
    InMux I__2565 (
            .O(N__10683),
            .I(N__10656));
    InMux I__2564 (
            .O(N__10680),
            .I(N__10656));
    InMux I__2563 (
            .O(N__10679),
            .I(N__10651));
    InMux I__2562 (
            .O(N__10678),
            .I(N__10648));
    InMux I__2561 (
            .O(N__10675),
            .I(N__10642));
    CascadeMux I__2560 (
            .O(N__10674),
            .I(N__10636));
    InMux I__2559 (
            .O(N__10673),
            .I(N__10626));
    InMux I__2558 (
            .O(N__10672),
            .I(N__10626));
    InMux I__2557 (
            .O(N__10671),
            .I(N__10626));
    InMux I__2556 (
            .O(N__10670),
            .I(N__10626));
    LocalMux I__2555 (
            .O(N__10667),
            .I(N__10617));
    Span4Mux_h I__2554 (
            .O(N__10664),
            .I(N__10617));
    LocalMux I__2553 (
            .O(N__10661),
            .I(N__10617));
    LocalMux I__2552 (
            .O(N__10656),
            .I(N__10617));
    InMux I__2551 (
            .O(N__10655),
            .I(N__10612));
    InMux I__2550 (
            .O(N__10654),
            .I(N__10612));
    LocalMux I__2549 (
            .O(N__10651),
            .I(N__10607));
    LocalMux I__2548 (
            .O(N__10648),
            .I(N__10607));
    InMux I__2547 (
            .O(N__10647),
            .I(N__10604));
    InMux I__2546 (
            .O(N__10646),
            .I(N__10599));
    InMux I__2545 (
            .O(N__10645),
            .I(N__10599));
    LocalMux I__2544 (
            .O(N__10642),
            .I(N__10596));
    InMux I__2543 (
            .O(N__10641),
            .I(N__10591));
    InMux I__2542 (
            .O(N__10640),
            .I(N__10591));
    InMux I__2541 (
            .O(N__10639),
            .I(N__10588));
    InMux I__2540 (
            .O(N__10636),
            .I(N__10585));
    InMux I__2539 (
            .O(N__10635),
            .I(N__10582));
    LocalMux I__2538 (
            .O(N__10626),
            .I(N__10575));
    Span4Mux_h I__2537 (
            .O(N__10617),
            .I(N__10575));
    LocalMux I__2536 (
            .O(N__10612),
            .I(N__10575));
    Span4Mux_v I__2535 (
            .O(N__10607),
            .I(N__10570));
    LocalMux I__2534 (
            .O(N__10604),
            .I(N__10567));
    LocalMux I__2533 (
            .O(N__10599),
            .I(N__10564));
    Span4Mux_h I__2532 (
            .O(N__10596),
            .I(N__10555));
    LocalMux I__2531 (
            .O(N__10591),
            .I(N__10555));
    LocalMux I__2530 (
            .O(N__10588),
            .I(N__10555));
    LocalMux I__2529 (
            .O(N__10585),
            .I(N__10555));
    LocalMux I__2528 (
            .O(N__10582),
            .I(N__10552));
    Span4Mux_v I__2527 (
            .O(N__10575),
            .I(N__10549));
    InMux I__2526 (
            .O(N__10574),
            .I(N__10546));
    InMux I__2525 (
            .O(N__10573),
            .I(N__10543));
    Span4Mux_h I__2524 (
            .O(N__10570),
            .I(N__10536));
    Span4Mux_v I__2523 (
            .O(N__10567),
            .I(N__10536));
    Span4Mux_v I__2522 (
            .O(N__10564),
            .I(N__10536));
    Span4Mux_h I__2521 (
            .O(N__10555),
            .I(N__10533));
    Span4Mux_h I__2520 (
            .O(N__10552),
            .I(N__10528));
    Span4Mux_h I__2519 (
            .O(N__10549),
            .I(N__10528));
    LocalMux I__2518 (
            .O(N__10546),
            .I(CPU_CYCLE));
    LocalMux I__2517 (
            .O(N__10543),
            .I(CPU_CYCLE));
    Odrv4 I__2516 (
            .O(N__10536),
            .I(CPU_CYCLE));
    Odrv4 I__2515 (
            .O(N__10533),
            .I(CPU_CYCLE));
    Odrv4 I__2514 (
            .O(N__10528),
            .I(CPU_CYCLE));
    InMux I__2513 (
            .O(N__10517),
            .I(N__10513));
    InMux I__2512 (
            .O(N__10516),
            .I(N__10510));
    LocalMux I__2511 (
            .O(N__10513),
            .I(N__10505));
    LocalMux I__2510 (
            .O(N__10510),
            .I(N__10505));
    Span4Mux_v I__2509 (
            .O(N__10505),
            .I(N__10502));
    Odrv4 I__2508 (
            .O(N__10502),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0Z0Z_0 ));
    CascadeMux I__2507 (
            .O(N__10499),
            .I(\U712_BYTE_ENABLE.N_91_cascade_ ));
    IoInMux I__2506 (
            .O(N__10496),
            .I(N__10493));
    LocalMux I__2505 (
            .O(N__10493),
            .I(N__10490));
    Span4Mux_s2_h I__2504 (
            .O(N__10490),
            .I(N__10487));
    Sp12to4 I__2503 (
            .O(N__10487),
            .I(N__10484));
    Span12Mux_v I__2502 (
            .O(N__10484),
            .I(N__10481));
    Span12Mux_h I__2501 (
            .O(N__10481),
            .I(N__10478));
    Odrv12 I__2500 (
            .O(N__10478),
            .I(N_51_i));
    InMux I__2499 (
            .O(N__10475),
            .I(N__10472));
    LocalMux I__2498 (
            .O(N__10472),
            .I(\U712_BYTE_ENABLE.N_89 ));
    IoInMux I__2497 (
            .O(N__10469),
            .I(N__10466));
    LocalMux I__2496 (
            .O(N__10466),
            .I(N__10463));
    IoSpan4Mux I__2495 (
            .O(N__10463),
            .I(N__10460));
    Span4Mux_s3_v I__2494 (
            .O(N__10460),
            .I(N__10457));
    Odrv4 I__2493 (
            .O(N__10457),
            .I(N_90_i));
    IoInMux I__2492 (
            .O(N__10454),
            .I(N__10451));
    LocalMux I__2491 (
            .O(N__10451),
            .I(N__10448));
    IoSpan4Mux I__2490 (
            .O(N__10448),
            .I(N__10445));
    Span4Mux_s2_v I__2489 (
            .O(N__10445),
            .I(N__10442));
    Span4Mux_v I__2488 (
            .O(N__10442),
            .I(N__10439));
    Odrv4 I__2487 (
            .O(N__10439),
            .I(N_92_i));
    IoInMux I__2486 (
            .O(N__10436),
            .I(N__10433));
    LocalMux I__2485 (
            .O(N__10433),
            .I(N__10430));
    Span4Mux_s3_v I__2484 (
            .O(N__10430),
            .I(N__10427));
    Odrv4 I__2483 (
            .O(N__10427),
            .I(N_91_i));
    CascadeMux I__2482 (
            .O(N__10424),
            .I(N__10420));
    CascadeMux I__2481 (
            .O(N__10423),
            .I(N__10417));
    InMux I__2480 (
            .O(N__10420),
            .I(N__10413));
    InMux I__2479 (
            .O(N__10417),
            .I(N__10408));
    InMux I__2478 (
            .O(N__10416),
            .I(N__10408));
    LocalMux I__2477 (
            .O(N__10413),
            .I(N__10400));
    LocalMux I__2476 (
            .O(N__10408),
            .I(N__10397));
    InMux I__2475 (
            .O(N__10407),
            .I(N__10394));
    InMux I__2474 (
            .O(N__10406),
            .I(N__10385));
    InMux I__2473 (
            .O(N__10405),
            .I(N__10385));
    InMux I__2472 (
            .O(N__10404),
            .I(N__10385));
    InMux I__2471 (
            .O(N__10403),
            .I(N__10385));
    Span4Mux_v I__2470 (
            .O(N__10400),
            .I(N__10382));
    Sp12to4 I__2469 (
            .O(N__10397),
            .I(N__10377));
    LocalMux I__2468 (
            .O(N__10394),
            .I(N__10377));
    LocalMux I__2467 (
            .O(N__10385),
            .I(N__10374));
    Span4Mux_v I__2466 (
            .O(N__10382),
            .I(N__10371));
    Span12Mux_h I__2465 (
            .O(N__10377),
            .I(N__10368));
    Span12Mux_v I__2464 (
            .O(N__10374),
            .I(N__10365));
    Span4Mux_v I__2463 (
            .O(N__10371),
            .I(N__10362));
    Span12Mux_v I__2462 (
            .O(N__10368),
            .I(N__10357));
    Span12Mux_h I__2461 (
            .O(N__10365),
            .I(N__10357));
    Sp12to4 I__2460 (
            .O(N__10362),
            .I(N__10354));
    Odrv12 I__2459 (
            .O(N__10357),
            .I(SIZ_c_1));
    Odrv12 I__2458 (
            .O(N__10354),
            .I(SIZ_c_1));
    InMux I__2457 (
            .O(N__10349),
            .I(N__10342));
    InMux I__2456 (
            .O(N__10348),
            .I(N__10342));
    InMux I__2455 (
            .O(N__10347),
            .I(N__10339));
    LocalMux I__2454 (
            .O(N__10342),
            .I(N__10332));
    LocalMux I__2453 (
            .O(N__10339),
            .I(N__10329));
    InMux I__2452 (
            .O(N__10338),
            .I(N__10320));
    InMux I__2451 (
            .O(N__10337),
            .I(N__10320));
    InMux I__2450 (
            .O(N__10336),
            .I(N__10320));
    InMux I__2449 (
            .O(N__10335),
            .I(N__10320));
    Span4Mux_v I__2448 (
            .O(N__10332),
            .I(N__10316));
    Span4Mux_v I__2447 (
            .O(N__10329),
            .I(N__10313));
    LocalMux I__2446 (
            .O(N__10320),
            .I(N__10310));
    InMux I__2445 (
            .O(N__10319),
            .I(N__10307));
    Span4Mux_v I__2444 (
            .O(N__10316),
            .I(N__10300));
    Span4Mux_v I__2443 (
            .O(N__10313),
            .I(N__10300));
    Span4Mux_v I__2442 (
            .O(N__10310),
            .I(N__10300));
    LocalMux I__2441 (
            .O(N__10307),
            .I(N__10297));
    Sp12to4 I__2440 (
            .O(N__10300),
            .I(N__10294));
    Sp12to4 I__2439 (
            .O(N__10297),
            .I(N__10291));
    Span12Mux_h I__2438 (
            .O(N__10294),
            .I(N__10286));
    Span12Mux_v I__2437 (
            .O(N__10291),
            .I(N__10286));
    Odrv12 I__2436 (
            .O(N__10286),
            .I(A_c_1));
    CascadeMux I__2435 (
            .O(N__10283),
            .I(N__10278));
    CascadeMux I__2434 (
            .O(N__10282),
            .I(N__10273));
    InMux I__2433 (
            .O(N__10281),
            .I(N__10269));
    InMux I__2432 (
            .O(N__10278),
            .I(N__10260));
    InMux I__2431 (
            .O(N__10277),
            .I(N__10260));
    InMux I__2430 (
            .O(N__10276),
            .I(N__10260));
    InMux I__2429 (
            .O(N__10273),
            .I(N__10260));
    CascadeMux I__2428 (
            .O(N__10272),
            .I(N__10255));
    LocalMux I__2427 (
            .O(N__10269),
            .I(N__10252));
    LocalMux I__2426 (
            .O(N__10260),
            .I(N__10248));
    InMux I__2425 (
            .O(N__10259),
            .I(N__10245));
    InMux I__2424 (
            .O(N__10258),
            .I(N__10239));
    InMux I__2423 (
            .O(N__10255),
            .I(N__10239));
    Span4Mux_v I__2422 (
            .O(N__10252),
            .I(N__10236));
    InMux I__2421 (
            .O(N__10251),
            .I(N__10233));
    Span4Mux_h I__2420 (
            .O(N__10248),
            .I(N__10230));
    LocalMux I__2419 (
            .O(N__10245),
            .I(N__10227));
    InMux I__2418 (
            .O(N__10244),
            .I(N__10224));
    LocalMux I__2417 (
            .O(N__10239),
            .I(N__10217));
    Sp12to4 I__2416 (
            .O(N__10236),
            .I(N__10217));
    LocalMux I__2415 (
            .O(N__10233),
            .I(N__10217));
    Span4Mux_v I__2414 (
            .O(N__10230),
            .I(N__10214));
    Span4Mux_h I__2413 (
            .O(N__10227),
            .I(N__10209));
    LocalMux I__2412 (
            .O(N__10224),
            .I(N__10209));
    Span12Mux_h I__2411 (
            .O(N__10217),
            .I(N__10206));
    Span4Mux_h I__2410 (
            .O(N__10214),
            .I(N__10203));
    Sp12to4 I__2409 (
            .O(N__10209),
            .I(N__10200));
    Span12Mux_v I__2408 (
            .O(N__10206),
            .I(N__10197));
    Sp12to4 I__2407 (
            .O(N__10203),
            .I(N__10192));
    Span12Mux_v I__2406 (
            .O(N__10200),
            .I(N__10192));
    Odrv12 I__2405 (
            .O(N__10197),
            .I(SIZ_c_0));
    Odrv12 I__2404 (
            .O(N__10192),
            .I(SIZ_c_0));
    CascadeMux I__2403 (
            .O(N__10187),
            .I(N__10182));
    InMux I__2402 (
            .O(N__10186),
            .I(N__10174));
    InMux I__2401 (
            .O(N__10185),
            .I(N__10174));
    InMux I__2400 (
            .O(N__10182),
            .I(N__10171));
    CascadeMux I__2399 (
            .O(N__10181),
            .I(N__10168));
    CascadeMux I__2398 (
            .O(N__10180),
            .I(N__10164));
    CascadeMux I__2397 (
            .O(N__10179),
            .I(N__10161));
    LocalMux I__2396 (
            .O(N__10174),
            .I(N__10157));
    LocalMux I__2395 (
            .O(N__10171),
            .I(N__10154));
    InMux I__2394 (
            .O(N__10168),
            .I(N__10151));
    InMux I__2393 (
            .O(N__10167),
            .I(N__10142));
    InMux I__2392 (
            .O(N__10164),
            .I(N__10142));
    InMux I__2391 (
            .O(N__10161),
            .I(N__10142));
    InMux I__2390 (
            .O(N__10160),
            .I(N__10142));
    Span4Mux_h I__2389 (
            .O(N__10157),
            .I(N__10134));
    Span4Mux_v I__2388 (
            .O(N__10154),
            .I(N__10134));
    LocalMux I__2387 (
            .O(N__10151),
            .I(N__10134));
    LocalMux I__2386 (
            .O(N__10142),
            .I(N__10131));
    InMux I__2385 (
            .O(N__10141),
            .I(N__10127));
    Span4Mux_h I__2384 (
            .O(N__10134),
            .I(N__10124));
    Span4Mux_v I__2383 (
            .O(N__10131),
            .I(N__10121));
    InMux I__2382 (
            .O(N__10130),
            .I(N__10118));
    LocalMux I__2381 (
            .O(N__10127),
            .I(N__10115));
    Span4Mux_v I__2380 (
            .O(N__10124),
            .I(N__10112));
    Sp12to4 I__2379 (
            .O(N__10121),
            .I(N__10107));
    LocalMux I__2378 (
            .O(N__10118),
            .I(N__10107));
    Span4Mux_v I__2377 (
            .O(N__10115),
            .I(N__10104));
    Sp12to4 I__2376 (
            .O(N__10112),
            .I(N__10097));
    Span12Mux_h I__2375 (
            .O(N__10107),
            .I(N__10097));
    Sp12to4 I__2374 (
            .O(N__10104),
            .I(N__10097));
    Odrv12 I__2373 (
            .O(N__10097),
            .I(A_c_0));
    IoInMux I__2372 (
            .O(N__10094),
            .I(N__10091));
    LocalMux I__2371 (
            .O(N__10091),
            .I(N__10088));
    Span4Mux_s2_v I__2370 (
            .O(N__10088),
            .I(N__10085));
    Span4Mux_h I__2369 (
            .O(N__10085),
            .I(N__10082));
    Span4Mux_v I__2368 (
            .O(N__10082),
            .I(N__10079));
    Odrv4 I__2367 (
            .O(N__10079),
            .I(N_89_i));
    InMux I__2366 (
            .O(N__10076),
            .I(N__10072));
    InMux I__2365 (
            .O(N__10075),
            .I(N__10069));
    LocalMux I__2364 (
            .O(N__10072),
            .I(N__10062));
    LocalMux I__2363 (
            .O(N__10069),
            .I(N__10062));
    InMux I__2362 (
            .O(N__10068),
            .I(N__10059));
    InMux I__2361 (
            .O(N__10067),
            .I(N__10056));
    Span4Mux_v I__2360 (
            .O(N__10062),
            .I(N__10053));
    LocalMux I__2359 (
            .O(N__10059),
            .I(N__10050));
    LocalMux I__2358 (
            .O(N__10056),
            .I(N__10047));
    Span4Mux_h I__2357 (
            .O(N__10053),
            .I(N__10042));
    Span4Mux_v I__2356 (
            .O(N__10050),
            .I(N__10042));
    Span12Mux_v I__2355 (
            .O(N__10047),
            .I(N__10039));
    Span4Mux_v I__2354 (
            .O(N__10042),
            .I(N__10036));
    Span12Mux_h I__2353 (
            .O(N__10039),
            .I(N__10033));
    Sp12to4 I__2352 (
            .O(N__10036),
            .I(N__10030));
    Odrv12 I__2351 (
            .O(N__10033),
            .I(DRA_c_3));
    Odrv12 I__2350 (
            .O(N__10030),
            .I(DRA_c_3));
    InMux I__2349 (
            .O(N__10025),
            .I(N__10020));
    InMux I__2348 (
            .O(N__10024),
            .I(N__10016));
    InMux I__2347 (
            .O(N__10023),
            .I(N__10013));
    LocalMux I__2346 (
            .O(N__10020),
            .I(N__10010));
    InMux I__2345 (
            .O(N__10019),
            .I(N__10007));
    LocalMux I__2344 (
            .O(N__10016),
            .I(N__10004));
    LocalMux I__2343 (
            .O(N__10013),
            .I(N__10001));
    Span4Mux_h I__2342 (
            .O(N__10010),
            .I(N__9996));
    LocalMux I__2341 (
            .O(N__10007),
            .I(N__9996));
    Span4Mux_v I__2340 (
            .O(N__10004),
            .I(N__9993));
    Sp12to4 I__2339 (
            .O(N__10001),
            .I(N__9988));
    Sp12to4 I__2338 (
            .O(N__9996),
            .I(N__9988));
    Sp12to4 I__2337 (
            .O(N__9993),
            .I(N__9985));
    Span12Mux_v I__2336 (
            .O(N__9988),
            .I(N__9982));
    Span12Mux_h I__2335 (
            .O(N__9985),
            .I(N__9979));
    Span12Mux_h I__2334 (
            .O(N__9982),
            .I(N__9974));
    Span12Mux_v I__2333 (
            .O(N__9979),
            .I(N__9974));
    Odrv12 I__2332 (
            .O(N__9974),
            .I(DRA_c_2));
    InMux I__2331 (
            .O(N__9971),
            .I(N__9965));
    InMux I__2330 (
            .O(N__9970),
            .I(N__9962));
    InMux I__2329 (
            .O(N__9969),
            .I(N__9956));
    InMux I__2328 (
            .O(N__9968),
            .I(N__9952));
    LocalMux I__2327 (
            .O(N__9965),
            .I(N__9945));
    LocalMux I__2326 (
            .O(N__9962),
            .I(N__9942));
    InMux I__2325 (
            .O(N__9961),
            .I(N__9939));
    InMux I__2324 (
            .O(N__9960),
            .I(N__9934));
    InMux I__2323 (
            .O(N__9959),
            .I(N__9934));
    LocalMux I__2322 (
            .O(N__9956),
            .I(N__9929));
    InMux I__2321 (
            .O(N__9955),
            .I(N__9926));
    LocalMux I__2320 (
            .O(N__9952),
            .I(N__9921));
    InMux I__2319 (
            .O(N__9951),
            .I(N__9912));
    InMux I__2318 (
            .O(N__9950),
            .I(N__9912));
    InMux I__2317 (
            .O(N__9949),
            .I(N__9912));
    InMux I__2316 (
            .O(N__9948),
            .I(N__9912));
    Span4Mux_h I__2315 (
            .O(N__9945),
            .I(N__9904));
    Span4Mux_h I__2314 (
            .O(N__9942),
            .I(N__9897));
    LocalMux I__2313 (
            .O(N__9939),
            .I(N__9897));
    LocalMux I__2312 (
            .O(N__9934),
            .I(N__9897));
    InMux I__2311 (
            .O(N__9933),
            .I(N__9892));
    InMux I__2310 (
            .O(N__9932),
            .I(N__9892));
    Span4Mux_v I__2309 (
            .O(N__9929),
            .I(N__9889));
    LocalMux I__2308 (
            .O(N__9926),
            .I(N__9886));
    InMux I__2307 (
            .O(N__9925),
            .I(N__9881));
    InMux I__2306 (
            .O(N__9924),
            .I(N__9881));
    Span4Mux_h I__2305 (
            .O(N__9921),
            .I(N__9876));
    LocalMux I__2304 (
            .O(N__9912),
            .I(N__9876));
    InMux I__2303 (
            .O(N__9911),
            .I(N__9867));
    InMux I__2302 (
            .O(N__9910),
            .I(N__9867));
    InMux I__2301 (
            .O(N__9909),
            .I(N__9867));
    InMux I__2300 (
            .O(N__9908),
            .I(N__9867));
    InMux I__2299 (
            .O(N__9907),
            .I(N__9864));
    Span4Mux_h I__2298 (
            .O(N__9904),
            .I(N__9857));
    Span4Mux_h I__2297 (
            .O(N__9897),
            .I(N__9857));
    LocalMux I__2296 (
            .O(N__9892),
            .I(N__9857));
    Span4Mux_h I__2295 (
            .O(N__9889),
            .I(N__9854));
    Span4Mux_v I__2294 (
            .O(N__9886),
            .I(N__9851));
    LocalMux I__2293 (
            .O(N__9881),
            .I(N__9848));
    Sp12to4 I__2292 (
            .O(N__9876),
            .I(N__9839));
    LocalMux I__2291 (
            .O(N__9867),
            .I(N__9839));
    LocalMux I__2290 (
            .O(N__9864),
            .I(N__9839));
    Sp12to4 I__2289 (
            .O(N__9857),
            .I(N__9839));
    Sp12to4 I__2288 (
            .O(N__9854),
            .I(N__9834));
    Sp12to4 I__2287 (
            .O(N__9851),
            .I(N__9834));
    Span12Mux_h I__2286 (
            .O(N__9848),
            .I(N__9831));
    Span12Mux_v I__2285 (
            .O(N__9839),
            .I(N__9828));
    Span12Mux_h I__2284 (
            .O(N__9834),
            .I(N__9825));
    Span12Mux_v I__2283 (
            .O(N__9831),
            .I(N__9820));
    Span12Mux_h I__2282 (
            .O(N__9828),
            .I(N__9820));
    Span12Mux_v I__2281 (
            .O(N__9825),
            .I(N__9817));
    Odrv12 I__2280 (
            .O(N__9820),
            .I(AGNUS_REV_c));
    Odrv12 I__2279 (
            .O(N__9817),
            .I(AGNUS_REV_c));
    InMux I__2278 (
            .O(N__9812),
            .I(N__9809));
    LocalMux I__2277 (
            .O(N__9809),
            .I(N__9806));
    Span4Mux_h I__2276 (
            .O(N__9806),
            .I(N__9803));
    Odrv4 I__2275 (
            .O(N__9803),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    ClkMux I__2274 (
            .O(N__9800),
            .I(N__9785));
    ClkMux I__2273 (
            .O(N__9799),
            .I(N__9785));
    ClkMux I__2272 (
            .O(N__9798),
            .I(N__9785));
    ClkMux I__2271 (
            .O(N__9797),
            .I(N__9785));
    ClkMux I__2270 (
            .O(N__9796),
            .I(N__9785));
    GlobalMux I__2269 (
            .O(N__9785),
            .I(N__9782));
    gio2CtrlBuf I__2268 (
            .O(N__9782),
            .I(C3_c_g));
    CEMux I__2267 (
            .O(N__9779),
            .I(N__9749));
    CEMux I__2266 (
            .O(N__9778),
            .I(N__9749));
    CEMux I__2265 (
            .O(N__9777),
            .I(N__9749));
    CEMux I__2264 (
            .O(N__9776),
            .I(N__9749));
    CEMux I__2263 (
            .O(N__9775),
            .I(N__9749));
    CEMux I__2262 (
            .O(N__9774),
            .I(N__9749));
    CEMux I__2261 (
            .O(N__9773),
            .I(N__9749));
    CEMux I__2260 (
            .O(N__9772),
            .I(N__9749));
    CEMux I__2259 (
            .O(N__9771),
            .I(N__9749));
    CEMux I__2258 (
            .O(N__9770),
            .I(N__9749));
    GlobalMux I__2257 (
            .O(N__9749),
            .I(N__9746));
    gio2CtrlBuf I__2256 (
            .O(N__9746),
            .I(DBRn_c_i_0_g));
    InMux I__2255 (
            .O(N__9743),
            .I(N__9740));
    LocalMux I__2254 (
            .O(N__9740),
            .I(N__9720));
    ClkMux I__2253 (
            .O(N__9739),
            .I(N__9662));
    ClkMux I__2252 (
            .O(N__9738),
            .I(N__9662));
    ClkMux I__2251 (
            .O(N__9737),
            .I(N__9662));
    ClkMux I__2250 (
            .O(N__9736),
            .I(N__9662));
    ClkMux I__2249 (
            .O(N__9735),
            .I(N__9662));
    ClkMux I__2248 (
            .O(N__9734),
            .I(N__9662));
    ClkMux I__2247 (
            .O(N__9733),
            .I(N__9662));
    ClkMux I__2246 (
            .O(N__9732),
            .I(N__9662));
    ClkMux I__2245 (
            .O(N__9731),
            .I(N__9662));
    ClkMux I__2244 (
            .O(N__9730),
            .I(N__9662));
    ClkMux I__2243 (
            .O(N__9729),
            .I(N__9662));
    ClkMux I__2242 (
            .O(N__9728),
            .I(N__9662));
    ClkMux I__2241 (
            .O(N__9727),
            .I(N__9662));
    ClkMux I__2240 (
            .O(N__9726),
            .I(N__9662));
    ClkMux I__2239 (
            .O(N__9725),
            .I(N__9662));
    ClkMux I__2238 (
            .O(N__9724),
            .I(N__9662));
    ClkMux I__2237 (
            .O(N__9723),
            .I(N__9662));
    Glb2LocalMux I__2236 (
            .O(N__9720),
            .I(N__9662));
    ClkMux I__2235 (
            .O(N__9719),
            .I(N__9662));
    ClkMux I__2234 (
            .O(N__9718),
            .I(N__9662));
    ClkMux I__2233 (
            .O(N__9717),
            .I(N__9662));
    ClkMux I__2232 (
            .O(N__9716),
            .I(N__9662));
    ClkMux I__2231 (
            .O(N__9715),
            .I(N__9662));
    ClkMux I__2230 (
            .O(N__9714),
            .I(N__9662));
    ClkMux I__2229 (
            .O(N__9713),
            .I(N__9662));
    GlobalMux I__2228 (
            .O(N__9662),
            .I(CLK80_PLL));
    CEMux I__2227 (
            .O(N__9659),
            .I(N__9656));
    LocalMux I__2226 (
            .O(N__9656),
            .I(N__9651));
    CEMux I__2225 (
            .O(N__9655),
            .I(N__9648));
    CEMux I__2224 (
            .O(N__9654),
            .I(N__9644));
    Span4Mux_h I__2223 (
            .O(N__9651),
            .I(N__9639));
    LocalMux I__2222 (
            .O(N__9648),
            .I(N__9639));
    CEMux I__2221 (
            .O(N__9647),
            .I(N__9636));
    LocalMux I__2220 (
            .O(N__9644),
            .I(N__9631));
    Span4Mux_h I__2219 (
            .O(N__9639),
            .I(N__9631));
    LocalMux I__2218 (
            .O(N__9636),
            .I(N__9628));
    Odrv4 I__2217 (
            .O(N__9631),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv4 I__2216 (
            .O(N__9628),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    InMux I__2215 (
            .O(N__9623),
            .I(N__9620));
    LocalMux I__2214 (
            .O(N__9620),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__2213 (
            .O(N__9617),
            .I(N__9614));
    LocalMux I__2212 (
            .O(N__9614),
            .I(N__9608));
    InMux I__2211 (
            .O(N__9613),
            .I(N__9603));
    InMux I__2210 (
            .O(N__9612),
            .I(N__9603));
    InMux I__2209 (
            .O(N__9611),
            .I(N__9600));
    Span4Mux_v I__2208 (
            .O(N__9608),
            .I(N__9597));
    LocalMux I__2207 (
            .O(N__9603),
            .I(N__9592));
    LocalMux I__2206 (
            .O(N__9600),
            .I(N__9592));
    Span4Mux_v I__2205 (
            .O(N__9597),
            .I(N__9589));
    Sp12to4 I__2204 (
            .O(N__9592),
            .I(N__9586));
    Sp12to4 I__2203 (
            .O(N__9589),
            .I(N__9583));
    Span12Mux_v I__2202 (
            .O(N__9586),
            .I(N__9580));
    Span12Mux_h I__2201 (
            .O(N__9583),
            .I(N__9577));
    Span12Mux_h I__2200 (
            .O(N__9580),
            .I(N__9574));
    Odrv12 I__2199 (
            .O(N__9577),
            .I(DRA_c_5));
    Odrv12 I__2198 (
            .O(N__9574),
            .I(DRA_c_5));
    InMux I__2197 (
            .O(N__9569),
            .I(N__9563));
    InMux I__2196 (
            .O(N__9568),
            .I(N__9563));
    LocalMux I__2195 (
            .O(N__9563),
            .I(N__9560));
    Span4Mux_h I__2194 (
            .O(N__9560),
            .I(N__9557));
    Odrv4 I__2193 (
            .O(N__9557),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__2192 (
            .O(N__9554),
            .I(N__9550));
    InMux I__2191 (
            .O(N__9553),
            .I(N__9547));
    LocalMux I__2190 (
            .O(N__9550),
            .I(N__9541));
    LocalMux I__2189 (
            .O(N__9547),
            .I(N__9541));
    InMux I__2188 (
            .O(N__9546),
            .I(N__9538));
    Span4Mux_h I__2187 (
            .O(N__9541),
            .I(N__9532));
    LocalMux I__2186 (
            .O(N__9538),
            .I(N__9532));
    InMux I__2185 (
            .O(N__9537),
            .I(N__9529));
    Span4Mux_v I__2184 (
            .O(N__9532),
            .I(N__9526));
    LocalMux I__2183 (
            .O(N__9529),
            .I(N__9523));
    Span4Mux_v I__2182 (
            .O(N__9526),
            .I(N__9520));
    Span12Mux_v I__2181 (
            .O(N__9523),
            .I(N__9517));
    Sp12to4 I__2180 (
            .O(N__9520),
            .I(N__9514));
    Span12Mux_h I__2179 (
            .O(N__9517),
            .I(N__9511));
    Span12Mux_h I__2178 (
            .O(N__9514),
            .I(N__9508));
    Odrv12 I__2177 (
            .O(N__9511),
            .I(DRA_c_4));
    Odrv12 I__2176 (
            .O(N__9508),
            .I(DRA_c_4));
    InMux I__2175 (
            .O(N__9503),
            .I(N__9500));
    LocalMux I__2174 (
            .O(N__9500),
            .I(N__9497));
    Odrv4 I__2173 (
            .O(N__9497),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__2172 (
            .O(N__9494),
            .I(N__9491));
    LocalMux I__2171 (
            .O(N__9491),
            .I(N__9488));
    Odrv4 I__2170 (
            .O(N__9488),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__2169 (
            .O(N__9485),
            .I(N__9481));
    InMux I__2168 (
            .O(N__9484),
            .I(N__9478));
    LocalMux I__2167 (
            .O(N__9481),
            .I(N__9473));
    LocalMux I__2166 (
            .O(N__9478),
            .I(N__9470));
    InMux I__2165 (
            .O(N__9477),
            .I(N__9465));
    InMux I__2164 (
            .O(N__9476),
            .I(N__9465));
    Span4Mux_v I__2163 (
            .O(N__9473),
            .I(N__9462));
    Span4Mux_v I__2162 (
            .O(N__9470),
            .I(N__9459));
    LocalMux I__2161 (
            .O(N__9465),
            .I(N__9456));
    Sp12to4 I__2160 (
            .O(N__9462),
            .I(N__9451));
    Sp12to4 I__2159 (
            .O(N__9459),
            .I(N__9451));
    Span12Mux_v I__2158 (
            .O(N__9456),
            .I(N__9448));
    Span12Mux_h I__2157 (
            .O(N__9451),
            .I(N__9445));
    Span12Mux_h I__2156 (
            .O(N__9448),
            .I(N__9442));
    Odrv12 I__2155 (
            .O(N__9445),
            .I(DRA_c_8));
    Odrv12 I__2154 (
            .O(N__9442),
            .I(DRA_c_8));
    CascadeMux I__2153 (
            .O(N__9437),
            .I(N__9434));
    InMux I__2152 (
            .O(N__9434),
            .I(N__9431));
    LocalMux I__2151 (
            .O(N__9431),
            .I(N__9428));
    Odrv4 I__2150 (
            .O(N__9428),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__2149 (
            .O(N__9425),
            .I(N__9422));
    LocalMux I__2148 (
            .O(N__9422),
            .I(N__9419));
    Span12Mux_h I__2147 (
            .O(N__9419),
            .I(N__9416));
    Odrv12 I__2146 (
            .O(N__9416),
            .I(RAS0n_c));
    CascadeMux I__2145 (
            .O(N__9413),
            .I(N__9410));
    InMux I__2144 (
            .O(N__9410),
            .I(N__9407));
    LocalMux I__2143 (
            .O(N__9407),
            .I(N__9403));
    InMux I__2142 (
            .O(N__9406),
            .I(N__9400));
    Span4Mux_v I__2141 (
            .O(N__9403),
            .I(N__9393));
    LocalMux I__2140 (
            .O(N__9400),
            .I(N__9393));
    InMux I__2139 (
            .O(N__9399),
            .I(N__9388));
    InMux I__2138 (
            .O(N__9398),
            .I(N__9388));
    Span4Mux_h I__2137 (
            .O(N__9393),
            .I(N__9383));
    LocalMux I__2136 (
            .O(N__9388),
            .I(N__9383));
    Span4Mux_h I__2135 (
            .O(N__9383),
            .I(N__9380));
    Span4Mux_v I__2134 (
            .O(N__9380),
            .I(N__9377));
    Sp12to4 I__2133 (
            .O(N__9377),
            .I(N__9374));
    Span12Mux_v I__2132 (
            .O(N__9374),
            .I(N__9371));
    Odrv12 I__2131 (
            .O(N__9371),
            .I(DRA_c_9));
    InMux I__2130 (
            .O(N__9368),
            .I(N__9365));
    LocalMux I__2129 (
            .O(N__9365),
            .I(N__9362));
    Odrv4 I__2128 (
            .O(N__9362),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    InMux I__2127 (
            .O(N__9359),
            .I(N__9352));
    InMux I__2126 (
            .O(N__9358),
            .I(N__9352));
    InMux I__2125 (
            .O(N__9357),
            .I(N__9348));
    LocalMux I__2124 (
            .O(N__9352),
            .I(N__9345));
    InMux I__2123 (
            .O(N__9351),
            .I(N__9342));
    LocalMux I__2122 (
            .O(N__9348),
            .I(N__9335));
    Sp12to4 I__2121 (
            .O(N__9345),
            .I(N__9335));
    LocalMux I__2120 (
            .O(N__9342),
            .I(N__9335));
    Span12Mux_v I__2119 (
            .O(N__9335),
            .I(N__9332));
    Span12Mux_h I__2118 (
            .O(N__9332),
            .I(N__9329));
    Odrv12 I__2117 (
            .O(N__9329),
            .I(DRA_c_6));
    InMux I__2116 (
            .O(N__9326),
            .I(N__9318));
    InMux I__2115 (
            .O(N__9325),
            .I(N__9318));
    InMux I__2114 (
            .O(N__9324),
            .I(N__9315));
    InMux I__2113 (
            .O(N__9323),
            .I(N__9312));
    LocalMux I__2112 (
            .O(N__9318),
            .I(N__9309));
    LocalMux I__2111 (
            .O(N__9315),
            .I(N__9304));
    LocalMux I__2110 (
            .O(N__9312),
            .I(N__9304));
    Span4Mux_v I__2109 (
            .O(N__9309),
            .I(N__9301));
    Span4Mux_v I__2108 (
            .O(N__9304),
            .I(N__9298));
    Sp12to4 I__2107 (
            .O(N__9301),
            .I(N__9295));
    Sp12to4 I__2106 (
            .O(N__9298),
            .I(N__9292));
    Span12Mux_h I__2105 (
            .O(N__9295),
            .I(N__9289));
    Span12Mux_h I__2104 (
            .O(N__9292),
            .I(N__9286));
    Odrv12 I__2103 (
            .O(N__9289),
            .I(DRA_c_7));
    Odrv12 I__2102 (
            .O(N__9286),
            .I(DRA_c_7));
    CascadeMux I__2101 (
            .O(N__9281),
            .I(N__9278));
    InMux I__2100 (
            .O(N__9278),
            .I(N__9275));
    LocalMux I__2099 (
            .O(N__9275),
            .I(N__9272));
    Odrv12 I__2098 (
            .O(N__9272),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    IoInMux I__2097 (
            .O(N__9269),
            .I(N__9266));
    LocalMux I__2096 (
            .O(N__9266),
            .I(N__9263));
    Span4Mux_s2_h I__2095 (
            .O(N__9263),
            .I(N__9260));
    Sp12to4 I__2094 (
            .O(N__9260),
            .I(N__9257));
    Span12Mux_v I__2093 (
            .O(N__9257),
            .I(N__9254));
    Span12Mux_v I__2092 (
            .O(N__9254),
            .I(N__9251));
    Span12Mux_h I__2091 (
            .O(N__9251),
            .I(N__9248));
    Odrv12 I__2090 (
            .O(N__9248),
            .I(N_50_i));
    IoInMux I__2089 (
            .O(N__9245),
            .I(N__9242));
    LocalMux I__2088 (
            .O(N__9242),
            .I(N__9239));
    IoSpan4Mux I__2087 (
            .O(N__9239),
            .I(N__9236));
    Sp12to4 I__2086 (
            .O(N__9236),
            .I(N__9233));
    Span12Mux_s7_v I__2085 (
            .O(N__9233),
            .I(N__9230));
    Odrv12 I__2084 (
            .O(N__9230),
            .I(WEn_c));
    IoInMux I__2083 (
            .O(N__9227),
            .I(N__9224));
    LocalMux I__2082 (
            .O(N__9224),
            .I(N__9221));
    Span4Mux_s3_v I__2081 (
            .O(N__9221),
            .I(N__9218));
    Span4Mux_v I__2080 (
            .O(N__9218),
            .I(N__9215));
    Span4Mux_h I__2079 (
            .O(N__9215),
            .I(N__9212));
    Odrv4 I__2078 (
            .O(N__9212),
            .I(RASn_c));
    IoInMux I__2077 (
            .O(N__9209),
            .I(N__9206));
    LocalMux I__2076 (
            .O(N__9206),
            .I(N__9203));
    Span4Mux_s0_v I__2075 (
            .O(N__9203),
            .I(N__9200));
    Sp12to4 I__2074 (
            .O(N__9200),
            .I(N__9197));
    Span12Mux_h I__2073 (
            .O(N__9197),
            .I(N__9194));
    Odrv12 I__2072 (
            .O(N__9194),
            .I(CRCSn_c));
    InMux I__2071 (
            .O(N__9191),
            .I(N__9187));
    InMux I__2070 (
            .O(N__9190),
            .I(N__9184));
    LocalMux I__2069 (
            .O(N__9187),
            .I(N__9180));
    LocalMux I__2068 (
            .O(N__9184),
            .I(N__9177));
    InMux I__2067 (
            .O(N__9183),
            .I(N__9174));
    Span4Mux_v I__2066 (
            .O(N__9180),
            .I(N__9164));
    Span4Mux_h I__2065 (
            .O(N__9177),
            .I(N__9164));
    LocalMux I__2064 (
            .O(N__9174),
            .I(N__9164));
    InMux I__2063 (
            .O(N__9173),
            .I(N__9161));
    InMux I__2062 (
            .O(N__9172),
            .I(N__9158));
    InMux I__2061 (
            .O(N__9171),
            .I(N__9155));
    Span4Mux_h I__2060 (
            .O(N__9164),
            .I(N__9152));
    LocalMux I__2059 (
            .O(N__9161),
            .I(N__9149));
    LocalMux I__2058 (
            .O(N__9158),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__2057 (
            .O(N__9155),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__2056 (
            .O(N__9152),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv12 I__2055 (
            .O(N__9149),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    CascadeMux I__2054 (
            .O(N__9140),
            .I(N__9131));
    CascadeMux I__2053 (
            .O(N__9139),
            .I(N__9128));
    CascadeMux I__2052 (
            .O(N__9138),
            .I(N__9125));
    CascadeMux I__2051 (
            .O(N__9137),
            .I(N__9119));
    CascadeMux I__2050 (
            .O(N__9136),
            .I(N__9113));
    InMux I__2049 (
            .O(N__9135),
            .I(N__9110));
    InMux I__2048 (
            .O(N__9134),
            .I(N__9107));
    InMux I__2047 (
            .O(N__9131),
            .I(N__9104));
    InMux I__2046 (
            .O(N__9128),
            .I(N__9097));
    InMux I__2045 (
            .O(N__9125),
            .I(N__9097));
    InMux I__2044 (
            .O(N__9124),
            .I(N__9097));
    InMux I__2043 (
            .O(N__9123),
            .I(N__9094));
    CascadeMux I__2042 (
            .O(N__9122),
            .I(N__9091));
    InMux I__2041 (
            .O(N__9119),
            .I(N__9087));
    InMux I__2040 (
            .O(N__9118),
            .I(N__9080));
    InMux I__2039 (
            .O(N__9117),
            .I(N__9080));
    InMux I__2038 (
            .O(N__9116),
            .I(N__9080));
    InMux I__2037 (
            .O(N__9113),
            .I(N__9077));
    LocalMux I__2036 (
            .O(N__9110),
            .I(N__9072));
    LocalMux I__2035 (
            .O(N__9107),
            .I(N__9069));
    LocalMux I__2034 (
            .O(N__9104),
            .I(N__9059));
    LocalMux I__2033 (
            .O(N__9097),
            .I(N__9059));
    LocalMux I__2032 (
            .O(N__9094),
            .I(N__9059));
    InMux I__2031 (
            .O(N__9091),
            .I(N__9054));
    InMux I__2030 (
            .O(N__9090),
            .I(N__9054));
    LocalMux I__2029 (
            .O(N__9087),
            .I(N__9047));
    LocalMux I__2028 (
            .O(N__9080),
            .I(N__9047));
    LocalMux I__2027 (
            .O(N__9077),
            .I(N__9047));
    InMux I__2026 (
            .O(N__9076),
            .I(N__9044));
    InMux I__2025 (
            .O(N__9075),
            .I(N__9041));
    Span4Mux_v I__2024 (
            .O(N__9072),
            .I(N__9032));
    Span4Mux_h I__2023 (
            .O(N__9069),
            .I(N__9032));
    InMux I__2022 (
            .O(N__9068),
            .I(N__9025));
    InMux I__2021 (
            .O(N__9067),
            .I(N__9025));
    InMux I__2020 (
            .O(N__9066),
            .I(N__9025));
    Span4Mux_v I__2019 (
            .O(N__9059),
            .I(N__9020));
    LocalMux I__2018 (
            .O(N__9054),
            .I(N__9020));
    Span4Mux_v I__2017 (
            .O(N__9047),
            .I(N__9017));
    LocalMux I__2016 (
            .O(N__9044),
            .I(N__9014));
    LocalMux I__2015 (
            .O(N__9041),
            .I(N__9011));
    InMux I__2014 (
            .O(N__9040),
            .I(N__9002));
    InMux I__2013 (
            .O(N__9039),
            .I(N__9002));
    InMux I__2012 (
            .O(N__9038),
            .I(N__9002));
    InMux I__2011 (
            .O(N__9037),
            .I(N__9002));
    Span4Mux_h I__2010 (
            .O(N__9032),
            .I(N__8997));
    LocalMux I__2009 (
            .O(N__9025),
            .I(N__8997));
    Span4Mux_h I__2008 (
            .O(N__9020),
            .I(N__8994));
    Odrv4 I__2007 (
            .O(N__9017),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2006 (
            .O(N__9014),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2005 (
            .O(N__9011),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2004 (
            .O(N__9002),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2003 (
            .O(N__8997),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2002 (
            .O(N__8994),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    CascadeMux I__2001 (
            .O(N__8981),
            .I(N__8976));
    CascadeMux I__2000 (
            .O(N__8980),
            .I(N__8973));
    InMux I__1999 (
            .O(N__8979),
            .I(N__8969));
    InMux I__1998 (
            .O(N__8976),
            .I(N__8966));
    InMux I__1997 (
            .O(N__8973),
            .I(N__8963));
    CascadeMux I__1996 (
            .O(N__8972),
            .I(N__8960));
    LocalMux I__1995 (
            .O(N__8969),
            .I(N__8955));
    LocalMux I__1994 (
            .O(N__8966),
            .I(N__8955));
    LocalMux I__1993 (
            .O(N__8963),
            .I(N__8952));
    InMux I__1992 (
            .O(N__8960),
            .I(N__8949));
    Span4Mux_v I__1991 (
            .O(N__8955),
            .I(N__8946));
    Span4Mux_v I__1990 (
            .O(N__8952),
            .I(N__8941));
    LocalMux I__1989 (
            .O(N__8949),
            .I(N__8941));
    Odrv4 I__1988 (
            .O(N__8946),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__1987 (
            .O(N__8941),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    InMux I__1986 (
            .O(N__8936),
            .I(N__8932));
    InMux I__1985 (
            .O(N__8935),
            .I(N__8929));
    LocalMux I__1984 (
            .O(N__8932),
            .I(N__8923));
    LocalMux I__1983 (
            .O(N__8929),
            .I(N__8923));
    InMux I__1982 (
            .O(N__8928),
            .I(N__8920));
    Span4Mux_v I__1981 (
            .O(N__8923),
            .I(N__8916));
    LocalMux I__1980 (
            .O(N__8920),
            .I(N__8911));
    InMux I__1979 (
            .O(N__8919),
            .I(N__8908));
    Span4Mux_h I__1978 (
            .O(N__8916),
            .I(N__8905));
    InMux I__1977 (
            .O(N__8915),
            .I(N__8902));
    InMux I__1976 (
            .O(N__8914),
            .I(N__8899));
    Span4Mux_v I__1975 (
            .O(N__8911),
            .I(N__8894));
    LocalMux I__1974 (
            .O(N__8908),
            .I(N__8894));
    Odrv4 I__1973 (
            .O(N__8905),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1972 (
            .O(N__8902),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1971 (
            .O(N__8899),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1970 (
            .O(N__8894),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    IoInMux I__1969 (
            .O(N__8885),
            .I(N__8882));
    LocalMux I__1968 (
            .O(N__8882),
            .I(N__8879));
    Span12Mux_s10_v I__1967 (
            .O(N__8879),
            .I(N__8876));
    Odrv12 I__1966 (
            .O(N__8876),
            .I(CMA_c_10));
    InMux I__1965 (
            .O(N__8873),
            .I(N__8870));
    LocalMux I__1964 (
            .O(N__8870),
            .I(N__8867));
    Span4Mux_v I__1963 (
            .O(N__8867),
            .I(N__8864));
    Span4Mux_v I__1962 (
            .O(N__8864),
            .I(N__8861));
    Sp12to4 I__1961 (
            .O(N__8861),
            .I(N__8858));
    Span12Mux_h I__1960 (
            .O(N__8858),
            .I(N__8855));
    Odrv12 I__1959 (
            .O(N__8855),
            .I(A_c_17));
    IoInMux I__1958 (
            .O(N__8852),
            .I(N__8849));
    LocalMux I__1957 (
            .O(N__8849),
            .I(N__8846));
    IoSpan4Mux I__1956 (
            .O(N__8846),
            .I(N__8843));
    IoSpan4Mux I__1955 (
            .O(N__8843),
            .I(N__8840));
    Span4Mux_s3_h I__1954 (
            .O(N__8840),
            .I(N__8837));
    Sp12to4 I__1953 (
            .O(N__8837),
            .I(N__8834));
    Odrv12 I__1952 (
            .O(N__8834),
            .I(CMA_c_8));
    InMux I__1951 (
            .O(N__8831),
            .I(N__8828));
    LocalMux I__1950 (
            .O(N__8828),
            .I(N__8825));
    Odrv12 I__1949 (
            .O(N__8825),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    IoInMux I__1948 (
            .O(N__8822),
            .I(N__8819));
    LocalMux I__1947 (
            .O(N__8819),
            .I(N__8816));
    Span12Mux_s2_h I__1946 (
            .O(N__8816),
            .I(N__8813));
    Span12Mux_h I__1945 (
            .O(N__8813),
            .I(N__8810));
    Odrv12 I__1944 (
            .O(N__8810),
            .I(CMA_c_3));
    InMux I__1943 (
            .O(N__8807),
            .I(N__8804));
    LocalMux I__1942 (
            .O(N__8804),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ));
    IoInMux I__1941 (
            .O(N__8801),
            .I(N__8798));
    LocalMux I__1940 (
            .O(N__8798),
            .I(N__8795));
    Span4Mux_s2_h I__1939 (
            .O(N__8795),
            .I(N__8792));
    Sp12to4 I__1938 (
            .O(N__8792),
            .I(N__8789));
    Span12Mux_s10_v I__1937 (
            .O(N__8789),
            .I(N__8786));
    Span12Mux_h I__1936 (
            .O(N__8786),
            .I(N__8783));
    Odrv12 I__1935 (
            .O(N__8783),
            .I(CMA_c_6));
    InMux I__1934 (
            .O(N__8780),
            .I(N__8770));
    InMux I__1933 (
            .O(N__8779),
            .I(N__8765));
    InMux I__1932 (
            .O(N__8778),
            .I(N__8765));
    InMux I__1931 (
            .O(N__8777),
            .I(N__8762));
    InMux I__1930 (
            .O(N__8776),
            .I(N__8757));
    InMux I__1929 (
            .O(N__8775),
            .I(N__8757));
    CascadeMux I__1928 (
            .O(N__8774),
            .I(N__8754));
    CascadeMux I__1927 (
            .O(N__8773),
            .I(N__8751));
    LocalMux I__1926 (
            .O(N__8770),
            .I(N__8741));
    LocalMux I__1925 (
            .O(N__8765),
            .I(N__8741));
    LocalMux I__1924 (
            .O(N__8762),
            .I(N__8741));
    LocalMux I__1923 (
            .O(N__8757),
            .I(N__8741));
    InMux I__1922 (
            .O(N__8754),
            .I(N__8734));
    InMux I__1921 (
            .O(N__8751),
            .I(N__8734));
    InMux I__1920 (
            .O(N__8750),
            .I(N__8734));
    Odrv12 I__1919 (
            .O(N__8741),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__1918 (
            .O(N__8734),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    CascadeMux I__1917 (
            .O(N__8729),
            .I(N__8722));
    CascadeMux I__1916 (
            .O(N__8728),
            .I(N__8719));
    CascadeMux I__1915 (
            .O(N__8727),
            .I(N__8715));
    CascadeMux I__1914 (
            .O(N__8726),
            .I(N__8712));
    InMux I__1913 (
            .O(N__8725),
            .I(N__8705));
    InMux I__1912 (
            .O(N__8722),
            .I(N__8705));
    InMux I__1911 (
            .O(N__8719),
            .I(N__8705));
    InMux I__1910 (
            .O(N__8718),
            .I(N__8698));
    InMux I__1909 (
            .O(N__8715),
            .I(N__8698));
    InMux I__1908 (
            .O(N__8712),
            .I(N__8698));
    LocalMux I__1907 (
            .O(N__8705),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1 ));
    LocalMux I__1906 (
            .O(N__8698),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1 ));
    InMux I__1905 (
            .O(N__8693),
            .I(N__8690));
    LocalMux I__1904 (
            .O(N__8690),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ));
    IoInMux I__1903 (
            .O(N__8687),
            .I(N__8684));
    LocalMux I__1902 (
            .O(N__8684),
            .I(N__8681));
    IoSpan4Mux I__1901 (
            .O(N__8681),
            .I(N__8678));
    Span4Mux_s3_h I__1900 (
            .O(N__8678),
            .I(N__8675));
    Sp12to4 I__1899 (
            .O(N__8675),
            .I(N__8672));
    Span12Mux_h I__1898 (
            .O(N__8672),
            .I(N__8669));
    Odrv12 I__1897 (
            .O(N__8669),
            .I(CMA_c_4));
    InMux I__1896 (
            .O(N__8666),
            .I(N__8663));
    LocalMux I__1895 (
            .O(N__8663),
            .I(N__8660));
    Span4Mux_v I__1894 (
            .O(N__8660),
            .I(N__8657));
    Span4Mux_v I__1893 (
            .O(N__8657),
            .I(N__8654));
    Sp12to4 I__1892 (
            .O(N__8654),
            .I(N__8651));
    Span12Mux_h I__1891 (
            .O(N__8651),
            .I(N__8648));
    Odrv12 I__1890 (
            .O(N__8648),
            .I(A_c_19));
    InMux I__1889 (
            .O(N__8645),
            .I(N__8642));
    LocalMux I__1888 (
            .O(N__8642),
            .I(N__8638));
    InMux I__1887 (
            .O(N__8641),
            .I(N__8635));
    Span4Mux_v I__1886 (
            .O(N__8638),
            .I(N__8630));
    LocalMux I__1885 (
            .O(N__8635),
            .I(N__8627));
    InMux I__1884 (
            .O(N__8634),
            .I(N__8622));
    InMux I__1883 (
            .O(N__8633),
            .I(N__8622));
    Odrv4 I__1882 (
            .O(N__8630),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    Odrv12 I__1881 (
            .O(N__8627),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    LocalMux I__1880 (
            .O(N__8622),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    IoInMux I__1879 (
            .O(N__8615),
            .I(N__8612));
    LocalMux I__1878 (
            .O(N__8612),
            .I(N__8609));
    IoSpan4Mux I__1877 (
            .O(N__8609),
            .I(N__8606));
    IoSpan4Mux I__1876 (
            .O(N__8606),
            .I(N__8603));
    Span4Mux_s3_h I__1875 (
            .O(N__8603),
            .I(N__8600));
    Sp12to4 I__1874 (
            .O(N__8600),
            .I(N__8597));
    Odrv12 I__1873 (
            .O(N__8597),
            .I(CMA_c_9));
    InMux I__1872 (
            .O(N__8594),
            .I(N__8591));
    LocalMux I__1871 (
            .O(N__8591),
            .I(N__8588));
    Odrv4 I__1870 (
            .O(N__8588),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__1869 (
            .O(N__8585),
            .I(N__8579));
    InMux I__1868 (
            .O(N__8584),
            .I(N__8579));
    LocalMux I__1867 (
            .O(N__8579),
            .I(N__8576));
    Odrv4 I__1866 (
            .O(N__8576),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__1865 (
            .O(N__8573),
            .I(N__8570));
    LocalMux I__1864 (
            .O(N__8570),
            .I(N__8567));
    Odrv4 I__1863 (
            .O(N__8567),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__1862 (
            .O(N__8564),
            .I(N__8558));
    InMux I__1861 (
            .O(N__8563),
            .I(N__8558));
    LocalMux I__1860 (
            .O(N__8558),
            .I(N__8553));
    InMux I__1859 (
            .O(N__8557),
            .I(N__8548));
    InMux I__1858 (
            .O(N__8556),
            .I(N__8548));
    Span4Mux_v I__1857 (
            .O(N__8553),
            .I(N__8545));
    LocalMux I__1856 (
            .O(N__8548),
            .I(N__8542));
    Span4Mux_h I__1855 (
            .O(N__8545),
            .I(N__8539));
    Span12Mux_h I__1854 (
            .O(N__8542),
            .I(N__8534));
    Sp12to4 I__1853 (
            .O(N__8539),
            .I(N__8534));
    Span12Mux_v I__1852 (
            .O(N__8534),
            .I(N__8531));
    Odrv12 I__1851 (
            .O(N__8531),
            .I(DRA_c_1));
    InMux I__1850 (
            .O(N__8528),
            .I(N__8525));
    LocalMux I__1849 (
            .O(N__8525),
            .I(N__8522));
    Span4Mux_v I__1848 (
            .O(N__8522),
            .I(N__8518));
    InMux I__1847 (
            .O(N__8521),
            .I(N__8515));
    Sp12to4 I__1846 (
            .O(N__8518),
            .I(N__8510));
    LocalMux I__1845 (
            .O(N__8515),
            .I(N__8510));
    Span12Mux_h I__1844 (
            .O(N__8510),
            .I(N__8507));
    Span12Mux_v I__1843 (
            .O(N__8507),
            .I(N__8504));
    Odrv12 I__1842 (
            .O(N__8504),
            .I(DRA_c_0));
    InMux I__1841 (
            .O(N__8501),
            .I(N__8498));
    LocalMux I__1840 (
            .O(N__8498),
            .I(N__8495));
    Odrv12 I__1839 (
            .O(N__8495),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    CascadeMux I__1838 (
            .O(N__8492),
            .I(N__8485));
    InMux I__1837 (
            .O(N__8491),
            .I(N__8481));
    InMux I__1836 (
            .O(N__8490),
            .I(N__8476));
    InMux I__1835 (
            .O(N__8489),
            .I(N__8469));
    InMux I__1834 (
            .O(N__8488),
            .I(N__8469));
    InMux I__1833 (
            .O(N__8485),
            .I(N__8469));
    InMux I__1832 (
            .O(N__8484),
            .I(N__8466));
    LocalMux I__1831 (
            .O(N__8481),
            .I(N__8463));
    InMux I__1830 (
            .O(N__8480),
            .I(N__8458));
    InMux I__1829 (
            .O(N__8479),
            .I(N__8458));
    LocalMux I__1828 (
            .O(N__8476),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_0 ));
    LocalMux I__1827 (
            .O(N__8469),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_0 ));
    LocalMux I__1826 (
            .O(N__8466),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_0 ));
    Odrv4 I__1825 (
            .O(N__8463),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_0 ));
    LocalMux I__1824 (
            .O(N__8458),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_0 ));
    InMux I__1823 (
            .O(N__8447),
            .I(N__8444));
    LocalMux I__1822 (
            .O(N__8444),
            .I(\U712_REG_SM.N_369 ));
    IoInMux I__1821 (
            .O(N__8441),
            .I(N__8438));
    LocalMux I__1820 (
            .O(N__8438),
            .I(N__8435));
    IoSpan4Mux I__1819 (
            .O(N__8435),
            .I(N__8432));
    Span4Mux_s3_v I__1818 (
            .O(N__8432),
            .I(N__8429));
    Sp12to4 I__1817 (
            .O(N__8429),
            .I(N__8425));
    CascadeMux I__1816 (
            .O(N__8428),
            .I(N__8422));
    Span12Mux_h I__1815 (
            .O(N__8425),
            .I(N__8417));
    InMux I__1814 (
            .O(N__8422),
            .I(N__8414));
    InMux I__1813 (
            .O(N__8421),
            .I(N__8411));
    InMux I__1812 (
            .O(N__8420),
            .I(N__8408));
    Odrv12 I__1811 (
            .O(N__8417),
            .I(UDSn_c));
    LocalMux I__1810 (
            .O(N__8414),
            .I(UDSn_c));
    LocalMux I__1809 (
            .O(N__8411),
            .I(UDSn_c));
    LocalMux I__1808 (
            .O(N__8408),
            .I(UDSn_c));
    CascadeMux I__1807 (
            .O(N__8399),
            .I(N__8395));
    InMux I__1806 (
            .O(N__8398),
            .I(N__8385));
    InMux I__1805 (
            .O(N__8395),
            .I(N__8385));
    InMux I__1804 (
            .O(N__8394),
            .I(N__8385));
    InMux I__1803 (
            .O(N__8393),
            .I(N__8382));
    CascadeMux I__1802 (
            .O(N__8392),
            .I(N__8379));
    LocalMux I__1801 (
            .O(N__8385),
            .I(N__8370));
    LocalMux I__1800 (
            .O(N__8382),
            .I(N__8370));
    InMux I__1799 (
            .O(N__8379),
            .I(N__8367));
    InMux I__1798 (
            .O(N__8378),
            .I(N__8364));
    InMux I__1797 (
            .O(N__8377),
            .I(N__8359));
    InMux I__1796 (
            .O(N__8376),
            .I(N__8359));
    InMux I__1795 (
            .O(N__8375),
            .I(N__8356));
    Span4Mux_h I__1794 (
            .O(N__8370),
            .I(N__8353));
    LocalMux I__1793 (
            .O(N__8367),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_2 ));
    LocalMux I__1792 (
            .O(N__8364),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_2 ));
    LocalMux I__1791 (
            .O(N__8359),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_2 ));
    LocalMux I__1790 (
            .O(N__8356),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_2 ));
    Odrv4 I__1789 (
            .O(N__8353),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_2 ));
    InMux I__1788 (
            .O(N__8342),
            .I(N__8339));
    LocalMux I__1787 (
            .O(N__8339),
            .I(\U712_REG_SM.N_465 ));
    CascadeMux I__1786 (
            .O(N__8336),
            .I(N__8333));
    InMux I__1785 (
            .O(N__8333),
            .I(N__8328));
    CascadeMux I__1784 (
            .O(N__8332),
            .I(N__8323));
    InMux I__1783 (
            .O(N__8331),
            .I(N__8320));
    LocalMux I__1782 (
            .O(N__8328),
            .I(N__8314));
    InMux I__1781 (
            .O(N__8327),
            .I(N__8309));
    InMux I__1780 (
            .O(N__8326),
            .I(N__8309));
    InMux I__1779 (
            .O(N__8323),
            .I(N__8306));
    LocalMux I__1778 (
            .O(N__8320),
            .I(N__8303));
    InMux I__1777 (
            .O(N__8319),
            .I(N__8300));
    InMux I__1776 (
            .O(N__8318),
            .I(N__8295));
    InMux I__1775 (
            .O(N__8317),
            .I(N__8295));
    Odrv4 I__1774 (
            .O(N__8314),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1773 (
            .O(N__8309),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1772 (
            .O(N__8306),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__1771 (
            .O(N__8303),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1770 (
            .O(N__8300),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1769 (
            .O(N__8295),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    CascadeMux I__1768 (
            .O(N__8282),
            .I(N__8277));
    InMux I__1767 (
            .O(N__8281),
            .I(N__8274));
    InMux I__1766 (
            .O(N__8280),
            .I(N__8271));
    InMux I__1765 (
            .O(N__8277),
            .I(N__8268));
    LocalMux I__1764 (
            .O(N__8274),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__1763 (
            .O(N__8271),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__1762 (
            .O(N__8268),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    CascadeMux I__1761 (
            .O(N__8261),
            .I(N__8256));
    InMux I__1760 (
            .O(N__8260),
            .I(N__8252));
    InMux I__1759 (
            .O(N__8259),
            .I(N__8246));
    InMux I__1758 (
            .O(N__8256),
            .I(N__8243));
    InMux I__1757 (
            .O(N__8255),
            .I(N__8240));
    LocalMux I__1756 (
            .O(N__8252),
            .I(N__8237));
    InMux I__1755 (
            .O(N__8251),
            .I(N__8234));
    InMux I__1754 (
            .O(N__8250),
            .I(N__8229));
    InMux I__1753 (
            .O(N__8249),
            .I(N__8229));
    LocalMux I__1752 (
            .O(N__8246),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1751 (
            .O(N__8243),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1750 (
            .O(N__8240),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__1749 (
            .O(N__8237),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1748 (
            .O(N__8234),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1747 (
            .O(N__8229),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    InMux I__1746 (
            .O(N__8216),
            .I(N__8210));
    InMux I__1745 (
            .O(N__8215),
            .I(N__8203));
    InMux I__1744 (
            .O(N__8214),
            .I(N__8203));
    InMux I__1743 (
            .O(N__8213),
            .I(N__8203));
    LocalMux I__1742 (
            .O(N__8210),
            .I(\U712_REG_SM.N_288 ));
    LocalMux I__1741 (
            .O(N__8203),
            .I(\U712_REG_SM.N_288 ));
    IoInMux I__1740 (
            .O(N__8198),
            .I(N__8195));
    LocalMux I__1739 (
            .O(N__8195),
            .I(N__8192));
    IoSpan4Mux I__1738 (
            .O(N__8192),
            .I(N__8189));
    Sp12to4 I__1737 (
            .O(N__8189),
            .I(N__8186));
    Span12Mux_s7_v I__1736 (
            .O(N__8186),
            .I(N__8183));
    Odrv12 I__1735 (
            .O(N__8183),
            .I(CASn_c));
    InMux I__1734 (
            .O(N__8180),
            .I(N__8177));
    LocalMux I__1733 (
            .O(N__8177),
            .I(N__8174));
    Odrv4 I__1732 (
            .O(N__8174),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ));
    IoInMux I__1731 (
            .O(N__8171),
            .I(N__8168));
    LocalMux I__1730 (
            .O(N__8168),
            .I(N__8165));
    IoSpan4Mux I__1729 (
            .O(N__8165),
            .I(N__8162));
    Sp12to4 I__1728 (
            .O(N__8162),
            .I(N__8159));
    Span12Mux_s3_h I__1727 (
            .O(N__8159),
            .I(N__8156));
    Span12Mux_h I__1726 (
            .O(N__8156),
            .I(N__8153));
    Odrv12 I__1725 (
            .O(N__8153),
            .I(CMA_c_7));
    InMux I__1724 (
            .O(N__8150),
            .I(N__8147));
    LocalMux I__1723 (
            .O(N__8147),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ));
    InMux I__1722 (
            .O(N__8144),
            .I(N__8141));
    LocalMux I__1721 (
            .O(N__8141),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ));
    InMux I__1720 (
            .O(N__8138),
            .I(N__8135));
    LocalMux I__1719 (
            .O(N__8135),
            .I(N__8132));
    Odrv12 I__1718 (
            .O(N__8132),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ));
    InMux I__1717 (
            .O(N__8129),
            .I(N__8126));
    LocalMux I__1716 (
            .O(N__8126),
            .I(N__8123));
    Odrv12 I__1715 (
            .O(N__8123),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ));
    InMux I__1714 (
            .O(N__8120),
            .I(N__8117));
    LocalMux I__1713 (
            .O(N__8117),
            .I(N__8114));
    Span4Mux_h I__1712 (
            .O(N__8114),
            .I(N__8111));
    Odrv4 I__1711 (
            .O(N__8111),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__1710 (
            .O(N__8108),
            .I(N__8105));
    LocalMux I__1709 (
            .O(N__8105),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    CascadeMux I__1708 (
            .O(N__8102),
            .I(N__8099));
    InMux I__1707 (
            .O(N__8099),
            .I(N__8096));
    LocalMux I__1706 (
            .O(N__8096),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__1705 (
            .O(N__8093),
            .I(N__8090));
    LocalMux I__1704 (
            .O(N__8090),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__1703 (
            .O(N__8087),
            .I(N__8080));
    InMux I__1702 (
            .O(N__8086),
            .I(N__8077));
    InMux I__1701 (
            .O(N__8085),
            .I(N__8073));
    InMux I__1700 (
            .O(N__8084),
            .I(N__8068));
    InMux I__1699 (
            .O(N__8083),
            .I(N__8068));
    LocalMux I__1698 (
            .O(N__8080),
            .I(N__8063));
    LocalMux I__1697 (
            .O(N__8077),
            .I(N__8063));
    InMux I__1696 (
            .O(N__8076),
            .I(N__8060));
    LocalMux I__1695 (
            .O(N__8073),
            .I(\U712_REG_SM.LATCH_REG_0_sqmuxa ));
    LocalMux I__1694 (
            .O(N__8068),
            .I(\U712_REG_SM.LATCH_REG_0_sqmuxa ));
    Odrv4 I__1693 (
            .O(N__8063),
            .I(\U712_REG_SM.LATCH_REG_0_sqmuxa ));
    LocalMux I__1692 (
            .O(N__8060),
            .I(\U712_REG_SM.LATCH_REG_0_sqmuxa ));
    IoInMux I__1691 (
            .O(N__8051),
            .I(N__8048));
    LocalMux I__1690 (
            .O(N__8048),
            .I(N__8045));
    Span4Mux_s1_v I__1689 (
            .O(N__8045),
            .I(N__8041));
    InMux I__1688 (
            .O(N__8044),
            .I(N__8038));
    Sp12to4 I__1687 (
            .O(N__8041),
            .I(N__8035));
    LocalMux I__1686 (
            .O(N__8038),
            .I(N__8032));
    Span12Mux_h I__1685 (
            .O(N__8035),
            .I(N__8029));
    Span4Mux_v I__1684 (
            .O(N__8032),
            .I(N__8026));
    Span12Mux_v I__1683 (
            .O(N__8029),
            .I(N__8021));
    Sp12to4 I__1682 (
            .O(N__8026),
            .I(N__8021));
    Span12Mux_h I__1681 (
            .O(N__8021),
            .I(N__8018));
    Span12Mux_v I__1680 (
            .O(N__8018),
            .I(N__8015));
    Odrv12 I__1679 (
            .O(N__8015),
            .I(RAMENn_c));
    CascadeMux I__1678 (
            .O(N__8012),
            .I(N__8008));
    InMux I__1677 (
            .O(N__8011),
            .I(N__8005));
    InMux I__1676 (
            .O(N__8008),
            .I(N__8002));
    LocalMux I__1675 (
            .O(N__8005),
            .I(N__7999));
    LocalMux I__1674 (
            .O(N__8002),
            .I(N__7996));
    Span4Mux_v I__1673 (
            .O(N__7999),
            .I(N__7993));
    Span4Mux_v I__1672 (
            .O(N__7996),
            .I(N__7990));
    Span4Mux_h I__1671 (
            .O(N__7993),
            .I(N__7987));
    Sp12to4 I__1670 (
            .O(N__7990),
            .I(N__7984));
    Sp12to4 I__1669 (
            .O(N__7987),
            .I(N__7981));
    Span12Mux_h I__1668 (
            .O(N__7984),
            .I(N__7978));
    Span12Mux_v I__1667 (
            .O(N__7981),
            .I(N__7975));
    Odrv12 I__1666 (
            .O(N__7978),
            .I(TSn_c));
    Odrv12 I__1665 (
            .O(N__7975),
            .I(TSn_c));
    InMux I__1664 (
            .O(N__7970),
            .I(N__7964));
    InMux I__1663 (
            .O(N__7969),
            .I(N__7964));
    LocalMux I__1662 (
            .O(N__7964),
            .I(\U712_REG_SM.CYCLE_RUNZ0 ));
    InMux I__1661 (
            .O(N__7961),
            .I(N__7958));
    LocalMux I__1660 (
            .O(N__7958),
            .I(N__7954));
    InMux I__1659 (
            .O(N__7957),
            .I(N__7951));
    Span4Mux_h I__1658 (
            .O(N__7954),
            .I(N__7947));
    LocalMux I__1657 (
            .O(N__7951),
            .I(N__7944));
    InMux I__1656 (
            .O(N__7950),
            .I(N__7941));
    Odrv4 I__1655 (
            .O(N__7947),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_1 ));
    Odrv4 I__1654 (
            .O(N__7944),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_1 ));
    LocalMux I__1653 (
            .O(N__7941),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_1 ));
    InMux I__1652 (
            .O(N__7934),
            .I(N__7931));
    LocalMux I__1651 (
            .O(N__7931),
            .I(N__7928));
    Span4Mux_v I__1650 (
            .O(N__7928),
            .I(N__7923));
    InMux I__1649 (
            .O(N__7927),
            .I(N__7920));
    CascadeMux I__1648 (
            .O(N__7926),
            .I(N__7916));
    Span4Mux_v I__1647 (
            .O(N__7923),
            .I(N__7913));
    LocalMux I__1646 (
            .O(N__7920),
            .I(N__7910));
    InMux I__1645 (
            .O(N__7919),
            .I(N__7905));
    InMux I__1644 (
            .O(N__7916),
            .I(N__7905));
    Span4Mux_v I__1643 (
            .O(N__7913),
            .I(N__7900));
    Span4Mux_v I__1642 (
            .O(N__7910),
            .I(N__7900));
    LocalMux I__1641 (
            .O(N__7905),
            .I(N__7897));
    Sp12to4 I__1640 (
            .O(N__7900),
            .I(N__7894));
    Span12Mux_v I__1639 (
            .O(N__7897),
            .I(N__7891));
    Span12Mux_h I__1638 (
            .O(N__7894),
            .I(N__7888));
    Span12Mux_h I__1637 (
            .O(N__7891),
            .I(N__7885));
    Odrv12 I__1636 (
            .O(N__7888),
            .I(RnW_c));
    Odrv12 I__1635 (
            .O(N__7885),
            .I(RnW_c));
    InMux I__1634 (
            .O(N__7880),
            .I(N__7876));
    CascadeMux I__1633 (
            .O(N__7879),
            .I(N__7870));
    LocalMux I__1632 (
            .O(N__7876),
            .I(N__7867));
    InMux I__1631 (
            .O(N__7875),
            .I(N__7862));
    InMux I__1630 (
            .O(N__7874),
            .I(N__7862));
    InMux I__1629 (
            .O(N__7873),
            .I(N__7859));
    InMux I__1628 (
            .O(N__7870),
            .I(N__7856));
    Span4Mux_v I__1627 (
            .O(N__7867),
            .I(N__7851));
    LocalMux I__1626 (
            .O(N__7862),
            .I(N__7851));
    LocalMux I__1625 (
            .O(N__7859),
            .I(REG_WRITE_CYCLE));
    LocalMux I__1624 (
            .O(N__7856),
            .I(REG_WRITE_CYCLE));
    Odrv4 I__1623 (
            .O(N__7851),
            .I(REG_WRITE_CYCLE));
    CascadeMux I__1622 (
            .O(N__7844),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_cascade_ ));
    IoInMux I__1621 (
            .O(N__7841),
            .I(N__7838));
    LocalMux I__1620 (
            .O(N__7838),
            .I(N__7835));
    Span4Mux_s3_v I__1619 (
            .O(N__7835),
            .I(N__7832));
    Span4Mux_v I__1618 (
            .O(N__7832),
            .I(N__7829));
    Span4Mux_h I__1617 (
            .O(N__7829),
            .I(N__7826));
    Odrv4 I__1616 (
            .O(N__7826),
            .I(CMA_c_0));
    InMux I__1615 (
            .O(N__7823),
            .I(N__7820));
    LocalMux I__1614 (
            .O(N__7820),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ));
    IoInMux I__1613 (
            .O(N__7817),
            .I(N__7814));
    LocalMux I__1612 (
            .O(N__7814),
            .I(N__7811));
    Span4Mux_s3_v I__1611 (
            .O(N__7811),
            .I(N__7808));
    Span4Mux_v I__1610 (
            .O(N__7808),
            .I(N__7805));
    Span4Mux_v I__1609 (
            .O(N__7805),
            .I(N__7802));
    Odrv4 I__1608 (
            .O(N__7802),
            .I(CMA_c_2));
    InMux I__1607 (
            .O(N__7799),
            .I(N__7795));
    InMux I__1606 (
            .O(N__7798),
            .I(N__7792));
    LocalMux I__1605 (
            .O(N__7795),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    LocalMux I__1604 (
            .O(N__7792),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    InMux I__1603 (
            .O(N__7787),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__1602 (
            .O(N__7784),
            .I(N__7780));
    InMux I__1601 (
            .O(N__7783),
            .I(N__7777));
    LocalMux I__1600 (
            .O(N__7780),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    LocalMux I__1599 (
            .O(N__7777),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    InMux I__1598 (
            .O(N__7772),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__1597 (
            .O(N__7769),
            .I(N__7765));
    InMux I__1596 (
            .O(N__7768),
            .I(N__7762));
    LocalMux I__1595 (
            .O(N__7765),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__1594 (
            .O(N__7762),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__1593 (
            .O(N__7757),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    CascadeMux I__1592 (
            .O(N__7754),
            .I(N__7750));
    InMux I__1591 (
            .O(N__7753),
            .I(N__7747));
    InMux I__1590 (
            .O(N__7750),
            .I(N__7744));
    LocalMux I__1589 (
            .O(N__7747),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__1588 (
            .O(N__7744),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__1587 (
            .O(N__7739),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__1586 (
            .O(N__7736),
            .I(N__7732));
    InMux I__1585 (
            .O(N__7735),
            .I(N__7729));
    LocalMux I__1584 (
            .O(N__7732),
            .I(N__7726));
    LocalMux I__1583 (
            .O(N__7729),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    Odrv4 I__1582 (
            .O(N__7726),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__1581 (
            .O(N__7721),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__1580 (
            .O(N__7718),
            .I(N__7714));
    InMux I__1579 (
            .O(N__7717),
            .I(N__7711));
    LocalMux I__1578 (
            .O(N__7714),
            .I(N__7708));
    LocalMux I__1577 (
            .O(N__7711),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    Odrv4 I__1576 (
            .O(N__7708),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__1575 (
            .O(N__7703),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__1574 (
            .O(N__7700),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    InMux I__1573 (
            .O(N__7697),
            .I(N__7694));
    LocalMux I__1572 (
            .O(N__7694),
            .I(N__7690));
    InMux I__1571 (
            .O(N__7693),
            .I(N__7687));
    Span4Mux_h I__1570 (
            .O(N__7690),
            .I(N__7684));
    LocalMux I__1569 (
            .O(N__7687),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    Odrv4 I__1568 (
            .O(N__7684),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    ClkMux I__1567 (
            .O(N__7679),
            .I(N__7658));
    ClkMux I__1566 (
            .O(N__7678),
            .I(N__7658));
    ClkMux I__1565 (
            .O(N__7677),
            .I(N__7658));
    ClkMux I__1564 (
            .O(N__7676),
            .I(N__7658));
    ClkMux I__1563 (
            .O(N__7675),
            .I(N__7658));
    ClkMux I__1562 (
            .O(N__7674),
            .I(N__7658));
    ClkMux I__1561 (
            .O(N__7673),
            .I(N__7658));
    GlobalMux I__1560 (
            .O(N__7658),
            .I(N__7655));
    gio2CtrlBuf I__1559 (
            .O(N__7655),
            .I(C1_c_g));
    SRMux I__1558 (
            .O(N__7652),
            .I(N__7649));
    LocalMux I__1557 (
            .O(N__7649),
            .I(N__7646));
    Span4Mux_h I__1556 (
            .O(N__7646),
            .I(N__7643));
    Odrv4 I__1555 (
            .O(N__7643),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    InMux I__1554 (
            .O(N__7640),
            .I(N__7637));
    LocalMux I__1553 (
            .O(N__7637),
            .I(\U712_REG_SM.UDSn_7_iv_i_0_0 ));
    InMux I__1552 (
            .O(N__7634),
            .I(N__7630));
    InMux I__1551 (
            .O(N__7633),
            .I(N__7627));
    LocalMux I__1550 (
            .O(N__7630),
            .I(\U712_REG_SM.C1_SYNC_RNI5ITS1Z0Z_1 ));
    LocalMux I__1549 (
            .O(N__7627),
            .I(\U712_REG_SM.C1_SYNC_RNI5ITS1Z0Z_1 ));
    InMux I__1548 (
            .O(N__7622),
            .I(N__7619));
    LocalMux I__1547 (
            .O(N__7619),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ));
    InMux I__1546 (
            .O(N__7616),
            .I(N__7613));
    LocalMux I__1545 (
            .O(N__7613),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ));
    InMux I__1544 (
            .O(N__7610),
            .I(N__7607));
    LocalMux I__1543 (
            .O(N__7607),
            .I(N__7604));
    Odrv12 I__1542 (
            .O(N__7604),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ));
    InMux I__1541 (
            .O(N__7601),
            .I(N__7598));
    LocalMux I__1540 (
            .O(N__7598),
            .I(N__7595));
    Span12Mux_v I__1539 (
            .O(N__7595),
            .I(N__7592));
    Span12Mux_h I__1538 (
            .O(N__7592),
            .I(N__7589));
    Odrv12 I__1537 (
            .O(N__7589),
            .I(A_c_7));
    InMux I__1536 (
            .O(N__7586),
            .I(N__7583));
    LocalMux I__1535 (
            .O(N__7583),
            .I(\U712_CHIP_RAM.N_329 ));
    InMux I__1534 (
            .O(N__7580),
            .I(N__7577));
    LocalMux I__1533 (
            .O(N__7577),
            .I(N__7574));
    Sp12to4 I__1532 (
            .O(N__7574),
            .I(N__7571));
    Span12Mux_v I__1531 (
            .O(N__7571),
            .I(N__7568));
    Span12Mux_h I__1530 (
            .O(N__7568),
            .I(N__7565));
    Odrv12 I__1529 (
            .O(N__7565),
            .I(A_c_2));
    InMux I__1528 (
            .O(N__7562),
            .I(N__7559));
    LocalMux I__1527 (
            .O(N__7559),
            .I(N__7556));
    Span12Mux_v I__1526 (
            .O(N__7556),
            .I(N__7553));
    Span12Mux_h I__1525 (
            .O(N__7553),
            .I(N__7550));
    Odrv12 I__1524 (
            .O(N__7550),
            .I(A_c_9));
    InMux I__1523 (
            .O(N__7547),
            .I(N__7544));
    LocalMux I__1522 (
            .O(N__7544),
            .I(N__7541));
    Span4Mux_h I__1521 (
            .O(N__7541),
            .I(N__7538));
    Odrv4 I__1520 (
            .O(N__7538),
            .I(\U712_CHIP_RAM.REFRESH5lto7_0 ));
    InMux I__1519 (
            .O(N__7535),
            .I(N__7532));
    LocalMux I__1518 (
            .O(N__7532),
            .I(N__7529));
    Odrv4 I__1517 (
            .O(N__7529),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__1516 (
            .O(N__7526),
            .I(N__7523));
    LocalMux I__1515 (
            .O(N__7523),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__1514 (
            .O(N__7520),
            .I(bfn_12_10_0_));
    InMux I__1513 (
            .O(N__7517),
            .I(N__7513));
    IoInMux I__1512 (
            .O(N__7516),
            .I(N__7510));
    LocalMux I__1511 (
            .O(N__7513),
            .I(N__7507));
    LocalMux I__1510 (
            .O(N__7510),
            .I(N__7504));
    Span4Mux_v I__1509 (
            .O(N__7507),
            .I(N__7501));
    IoSpan4Mux I__1508 (
            .O(N__7504),
            .I(N__7498));
    Sp12to4 I__1507 (
            .O(N__7501),
            .I(N__7495));
    IoSpan4Mux I__1506 (
            .O(N__7498),
            .I(N__7492));
    Span12Mux_h I__1505 (
            .O(N__7495),
            .I(N__7489));
    IoSpan4Mux I__1504 (
            .O(N__7492),
            .I(N__7486));
    Odrv12 I__1503 (
            .O(N__7489),
            .I(C1_c));
    Odrv4 I__1502 (
            .O(N__7486),
            .I(C1_c));
    InMux I__1501 (
            .O(N__7481),
            .I(N__7478));
    LocalMux I__1500 (
            .O(N__7478),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    CascadeMux I__1499 (
            .O(N__7475),
            .I(N__7472));
    InMux I__1498 (
            .O(N__7472),
            .I(N__7469));
    LocalMux I__1497 (
            .O(N__7469),
            .I(N__7466));
    Odrv4 I__1496 (
            .O(N__7466),
            .I(\U712_REG_SM.LDSn_7_iv_i_0_0 ));
    InMux I__1495 (
            .O(N__7463),
            .I(N__7460));
    LocalMux I__1494 (
            .O(N__7460),
            .I(\U712_REG_SM.N_278 ));
    IoInMux I__1493 (
            .O(N__7457),
            .I(N__7454));
    LocalMux I__1492 (
            .O(N__7454),
            .I(N__7451));
    IoSpan4Mux I__1491 (
            .O(N__7451),
            .I(N__7448));
    Span4Mux_s3_v I__1490 (
            .O(N__7448),
            .I(N__7445));
    Sp12to4 I__1489 (
            .O(N__7445),
            .I(N__7442));
    Span12Mux_s11_v I__1488 (
            .O(N__7442),
            .I(N__7438));
    InMux I__1487 (
            .O(N__7441),
            .I(N__7435));
    Odrv12 I__1486 (
            .O(N__7438),
            .I(ASn_c));
    LocalMux I__1485 (
            .O(N__7435),
            .I(ASn_c));
    CascadeMux I__1484 (
            .O(N__7430),
            .I(N__7427));
    InMux I__1483 (
            .O(N__7427),
            .I(N__7423));
    InMux I__1482 (
            .O(N__7426),
            .I(N__7420));
    LocalMux I__1481 (
            .O(N__7423),
            .I(N__7411));
    LocalMux I__1480 (
            .O(N__7420),
            .I(N__7411));
    InMux I__1479 (
            .O(N__7419),
            .I(N__7407));
    InMux I__1478 (
            .O(N__7418),
            .I(N__7401));
    InMux I__1477 (
            .O(N__7417),
            .I(N__7401));
    InMux I__1476 (
            .O(N__7416),
            .I(N__7398));
    Span12Mux_v I__1475 (
            .O(N__7411),
            .I(N__7395));
    InMux I__1474 (
            .O(N__7410),
            .I(N__7392));
    LocalMux I__1473 (
            .O(N__7407),
            .I(N__7389));
    InMux I__1472 (
            .O(N__7406),
            .I(N__7386));
    LocalMux I__1471 (
            .O(N__7401),
            .I(N__7381));
    LocalMux I__1470 (
            .O(N__7398),
            .I(N__7381));
    Odrv12 I__1469 (
            .O(N__7395),
            .I(WRITE_CYCLE));
    LocalMux I__1468 (
            .O(N__7392),
            .I(WRITE_CYCLE));
    Odrv4 I__1467 (
            .O(N__7389),
            .I(WRITE_CYCLE));
    LocalMux I__1466 (
            .O(N__7386),
            .I(WRITE_CYCLE));
    Odrv4 I__1465 (
            .O(N__7381),
            .I(WRITE_CYCLE));
    IoInMux I__1464 (
            .O(N__7370),
            .I(N__7367));
    LocalMux I__1463 (
            .O(N__7367),
            .I(N__7364));
    Span4Mux_s0_v I__1462 (
            .O(N__7364),
            .I(N__7361));
    Sp12to4 I__1461 (
            .O(N__7361),
            .I(N__7358));
    Span12Mux_h I__1460 (
            .O(N__7358),
            .I(N__7355));
    Odrv12 I__1459 (
            .O(N__7355),
            .I(N_259));
    IoInMux I__1458 (
            .O(N__7352),
            .I(N__7349));
    LocalMux I__1457 (
            .O(N__7349),
            .I(N__7346));
    IoSpan4Mux I__1456 (
            .O(N__7346),
            .I(N__7343));
    Sp12to4 I__1455 (
            .O(N__7343),
            .I(N__7340));
    Span12Mux_v I__1454 (
            .O(N__7340),
            .I(N__7337));
    Span12Mux_h I__1453 (
            .O(N__7337),
            .I(N__7331));
    InMux I__1452 (
            .O(N__7336),
            .I(N__7328));
    InMux I__1451 (
            .O(N__7335),
            .I(N__7325));
    InMux I__1450 (
            .O(N__7334),
            .I(N__7322));
    Odrv12 I__1449 (
            .O(N__7331),
            .I(LDSn_c));
    LocalMux I__1448 (
            .O(N__7328),
            .I(LDSn_c));
    LocalMux I__1447 (
            .O(N__7325),
            .I(LDSn_c));
    LocalMux I__1446 (
            .O(N__7322),
            .I(LDSn_c));
    CascadeMux I__1445 (
            .O(N__7313),
            .I(\U712_REG_SM.N_467_cascade_ ));
    InMux I__1444 (
            .O(N__7310),
            .I(N__7307));
    LocalMux I__1443 (
            .O(N__7307),
            .I(\U712_REG_SM.N_371 ));
    InMux I__1442 (
            .O(N__7304),
            .I(N__7301));
    LocalMux I__1441 (
            .O(N__7301),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ));
    IoInMux I__1440 (
            .O(N__7298),
            .I(N__7295));
    LocalMux I__1439 (
            .O(N__7295),
            .I(N__7292));
    Odrv12 I__1438 (
            .O(N__7292),
            .I(CMA_c_1));
    InMux I__1437 (
            .O(N__7289),
            .I(N__7286));
    LocalMux I__1436 (
            .O(N__7286),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ));
    InMux I__1435 (
            .O(N__7283),
            .I(N__7280));
    LocalMux I__1434 (
            .O(N__7280),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ));
    IoInMux I__1433 (
            .O(N__7277),
            .I(N__7274));
    LocalMux I__1432 (
            .O(N__7274),
            .I(N__7271));
    IoSpan4Mux I__1431 (
            .O(N__7271),
            .I(N__7268));
    Span4Mux_s2_h I__1430 (
            .O(N__7268),
            .I(N__7265));
    Sp12to4 I__1429 (
            .O(N__7265),
            .I(N__7262));
    Span12Mux_h I__1428 (
            .O(N__7262),
            .I(N__7259));
    Odrv12 I__1427 (
            .O(N__7259),
            .I(CMA_c_5));
    InMux I__1426 (
            .O(N__7256),
            .I(N__7253));
    LocalMux I__1425 (
            .O(N__7253),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ));
    CascadeMux I__1424 (
            .O(N__7250),
            .I(N__7247));
    InMux I__1423 (
            .O(N__7247),
            .I(N__7244));
    LocalMux I__1422 (
            .O(N__7244),
            .I(\U712_BYTE_ENABLE.N_92 ));
    IoInMux I__1421 (
            .O(N__7241),
            .I(N__7238));
    LocalMux I__1420 (
            .O(N__7238),
            .I(N__7235));
    IoSpan4Mux I__1419 (
            .O(N__7235),
            .I(N__7232));
    Span4Mux_s2_h I__1418 (
            .O(N__7232),
            .I(N__7229));
    Sp12to4 I__1417 (
            .O(N__7229),
            .I(N__7226));
    Span12Mux_s9_h I__1416 (
            .O(N__7226),
            .I(N__7223));
    Span12Mux_v I__1415 (
            .O(N__7223),
            .I(N__7220));
    Odrv12 I__1414 (
            .O(N__7220),
            .I(N_315));
    CascadeMux I__1413 (
            .O(N__7217),
            .I(\U712_REG_SM.N_278_cascade_ ));
    CascadeMux I__1412 (
            .O(N__7214),
            .I(N__7210));
    CascadeMux I__1411 (
            .O(N__7213),
            .I(N__7207));
    InMux I__1410 (
            .O(N__7210),
            .I(N__7200));
    InMux I__1409 (
            .O(N__7207),
            .I(N__7197));
    InMux I__1408 (
            .O(N__7206),
            .I(N__7192));
    InMux I__1407 (
            .O(N__7205),
            .I(N__7192));
    InMux I__1406 (
            .O(N__7204),
            .I(N__7187));
    InMux I__1405 (
            .O(N__7203),
            .I(N__7187));
    LocalMux I__1404 (
            .O(N__7200),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_7 ));
    LocalMux I__1403 (
            .O(N__7197),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_7 ));
    LocalMux I__1402 (
            .O(N__7192),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_7 ));
    LocalMux I__1401 (
            .O(N__7187),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_7 ));
    InMux I__1400 (
            .O(N__7178),
            .I(N__7175));
    LocalMux I__1399 (
            .O(N__7175),
            .I(N__7171));
    InMux I__1398 (
            .O(N__7174),
            .I(N__7168));
    Odrv4 I__1397 (
            .O(N__7171),
            .I(\U712_REG_SM.N_272 ));
    LocalMux I__1396 (
            .O(N__7168),
            .I(\U712_REG_SM.N_272 ));
    InMux I__1395 (
            .O(N__7163),
            .I(N__7157));
    InMux I__1394 (
            .O(N__7162),
            .I(N__7157));
    LocalMux I__1393 (
            .O(N__7157),
            .I(\U712_REG_SM.N_309 ));
    CascadeMux I__1392 (
            .O(N__7154),
            .I(\U712_REG_SM.N_272_cascade_ ));
    IoInMux I__1391 (
            .O(N__7151),
            .I(N__7148));
    LocalMux I__1390 (
            .O(N__7148),
            .I(N__7145));
    IoSpan4Mux I__1389 (
            .O(N__7145),
            .I(N__7142));
    Span4Mux_s3_h I__1388 (
            .O(N__7142),
            .I(N__7139));
    Span4Mux_h I__1387 (
            .O(N__7139),
            .I(N__7136));
    Sp12to4 I__1386 (
            .O(N__7136),
            .I(N__7133));
    Span12Mux_h I__1385 (
            .O(N__7133),
            .I(N__7129));
    InMux I__1384 (
            .O(N__7132),
            .I(N__7126));
    Span12Mux_h I__1383 (
            .O(N__7129),
            .I(N__7123));
    LocalMux I__1382 (
            .O(N__7126),
            .I(N__7120));
    Span12Mux_v I__1381 (
            .O(N__7123),
            .I(N__7117));
    Span12Mux_h I__1380 (
            .O(N__7120),
            .I(N__7114));
    Odrv12 I__1379 (
            .O(N__7117),
            .I(C3_c));
    Odrv12 I__1378 (
            .O(N__7114),
            .I(C3_c));
    InMux I__1377 (
            .O(N__7109),
            .I(N__7106));
    LocalMux I__1376 (
            .O(N__7106),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    InMux I__1375 (
            .O(N__7103),
            .I(N__7100));
    LocalMux I__1374 (
            .O(N__7100),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ));
    InMux I__1373 (
            .O(N__7097),
            .I(N__7091));
    InMux I__1372 (
            .O(N__7096),
            .I(N__7091));
    LocalMux I__1371 (
            .O(N__7091),
            .I(N__7088));
    Span4Mux_v I__1370 (
            .O(N__7088),
            .I(N__7085));
    Span4Mux_v I__1369 (
            .O(N__7085),
            .I(N__7082));
    Sp12to4 I__1368 (
            .O(N__7082),
            .I(N__7079));
    Span12Mux_h I__1367 (
            .O(N__7079),
            .I(N__7076));
    Odrv12 I__1366 (
            .O(N__7076),
            .I(A_c_14));
    InMux I__1365 (
            .O(N__7073),
            .I(N__7070));
    LocalMux I__1364 (
            .O(N__7070),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ));
    InMux I__1363 (
            .O(N__7067),
            .I(N__7064));
    LocalMux I__1362 (
            .O(N__7064),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__1361 (
            .O(N__7061),
            .I(N__7058));
    LocalMux I__1360 (
            .O(N__7058),
            .I(N__7055));
    Odrv4 I__1359 (
            .O(N__7055),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    IoInMux I__1358 (
            .O(N__7052),
            .I(N__7049));
    LocalMux I__1357 (
            .O(N__7049),
            .I(N__7046));
    Span4Mux_s2_v I__1356 (
            .O(N__7046),
            .I(N__7043));
    Span4Mux_h I__1355 (
            .O(N__7043),
            .I(N__7040));
    Sp12to4 I__1354 (
            .O(N__7040),
            .I(N__7036));
    InMux I__1353 (
            .O(N__7039),
            .I(N__7033));
    Span12Mux_v I__1352 (
            .O(N__7036),
            .I(N__7026));
    LocalMux I__1351 (
            .O(N__7033),
            .I(N__7026));
    InMux I__1350 (
            .O(N__7032),
            .I(N__7023));
    InMux I__1349 (
            .O(N__7031),
            .I(N__7020));
    Odrv12 I__1348 (
            .O(N__7026),
            .I(DBENn_c));
    LocalMux I__1347 (
            .O(N__7023),
            .I(DBENn_c));
    LocalMux I__1346 (
            .O(N__7020),
            .I(DBENn_c));
    CascadeMux I__1345 (
            .O(N__7013),
            .I(N__7009));
    InMux I__1344 (
            .O(N__7012),
            .I(N__7005));
    InMux I__1343 (
            .O(N__7009),
            .I(N__7002));
    InMux I__1342 (
            .O(N__7008),
            .I(N__6997));
    LocalMux I__1341 (
            .O(N__7005),
            .I(N__6994));
    LocalMux I__1340 (
            .O(N__7002),
            .I(N__6991));
    InMux I__1339 (
            .O(N__7001),
            .I(N__6988));
    InMux I__1338 (
            .O(N__7000),
            .I(N__6984));
    LocalMux I__1337 (
            .O(N__6997),
            .I(N__6981));
    Span4Mux_v I__1336 (
            .O(N__6994),
            .I(N__6976));
    Span4Mux_v I__1335 (
            .O(N__6991),
            .I(N__6976));
    LocalMux I__1334 (
            .O(N__6988),
            .I(N__6973));
    InMux I__1333 (
            .O(N__6987),
            .I(N__6970));
    LocalMux I__1332 (
            .O(N__6984),
            .I(N__6967));
    Odrv12 I__1331 (
            .O(N__6981),
            .I(DMA_CYCLE));
    Odrv4 I__1330 (
            .O(N__6976),
            .I(DMA_CYCLE));
    Odrv4 I__1329 (
            .O(N__6973),
            .I(DMA_CYCLE));
    LocalMux I__1328 (
            .O(N__6970),
            .I(DMA_CYCLE));
    Odrv4 I__1327 (
            .O(N__6967),
            .I(DMA_CYCLE));
    InMux I__1326 (
            .O(N__6956),
            .I(N__6953));
    LocalMux I__1325 (
            .O(N__6953),
            .I(N__6950));
    Span4Mux_h I__1324 (
            .O(N__6950),
            .I(N__6947));
    Odrv4 I__1323 (
            .O(N__6947),
            .I(\U712_CHIP_RAM.REFRESH5lt7 ));
    InMux I__1322 (
            .O(N__6944),
            .I(N__6940));
    InMux I__1321 (
            .O(N__6943),
            .I(N__6937));
    LocalMux I__1320 (
            .O(N__6940),
            .I(N__6932));
    LocalMux I__1319 (
            .O(N__6937),
            .I(N__6932));
    Odrv12 I__1318 (
            .O(N__6932),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0Z0Z_0 ));
    IoInMux I__1317 (
            .O(N__6929),
            .I(N__6926));
    LocalMux I__1316 (
            .O(N__6926),
            .I(N__6923));
    IoSpan4Mux I__1315 (
            .O(N__6923),
            .I(N__6920));
    Span4Mux_s3_h I__1314 (
            .O(N__6920),
            .I(N__6917));
    Sp12to4 I__1313 (
            .O(N__6917),
            .I(N__6914));
    Span12Mux_h I__1312 (
            .O(N__6914),
            .I(N__6911));
    Span12Mux_v I__1311 (
            .O(N__6911),
            .I(N__6908));
    Odrv12 I__1310 (
            .O(N__6908),
            .I(N_49_i));
    InMux I__1309 (
            .O(N__6905),
            .I(N__6899));
    InMux I__1308 (
            .O(N__6904),
            .I(N__6899));
    LocalMux I__1307 (
            .O(N__6899),
            .I(\U712_REG_SM.STATE_COUNTERc_0 ));
    InMux I__1306 (
            .O(N__6896),
            .I(N__6893));
    LocalMux I__1305 (
            .O(N__6893),
            .I(\U712_REG_SM.un15_0_i_0_0 ));
    CascadeMux I__1304 (
            .O(N__6890),
            .I(N__6887));
    InMux I__1303 (
            .O(N__6887),
            .I(N__6884));
    LocalMux I__1302 (
            .O(N__6884),
            .I(\U712_REG_SM.N_297 ));
    InMux I__1301 (
            .O(N__6881),
            .I(N__6875));
    InMux I__1300 (
            .O(N__6880),
            .I(N__6872));
    InMux I__1299 (
            .O(N__6879),
            .I(N__6869));
    InMux I__1298 (
            .O(N__6878),
            .I(N__6866));
    LocalMux I__1297 (
            .O(N__6875),
            .I(N__6862));
    LocalMux I__1296 (
            .O(N__6872),
            .I(N__6857));
    LocalMux I__1295 (
            .O(N__6869),
            .I(N__6857));
    LocalMux I__1294 (
            .O(N__6866),
            .I(N__6854));
    InMux I__1293 (
            .O(N__6865),
            .I(N__6851));
    Span4Mux_v I__1292 (
            .O(N__6862),
            .I(N__6848));
    Span4Mux_h I__1291 (
            .O(N__6857),
            .I(N__6843));
    Span4Mux_h I__1290 (
            .O(N__6854),
            .I(N__6843));
    LocalMux I__1289 (
            .O(N__6851),
            .I(REG_TACK));
    Odrv4 I__1288 (
            .O(N__6848),
            .I(REG_TACK));
    Odrv4 I__1287 (
            .O(N__6843),
            .I(REG_TACK));
    InMux I__1286 (
            .O(N__6836),
            .I(N__6831));
    InMux I__1285 (
            .O(N__6835),
            .I(N__6828));
    InMux I__1284 (
            .O(N__6834),
            .I(N__6825));
    LocalMux I__1283 (
            .O(N__6831),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_6 ));
    LocalMux I__1282 (
            .O(N__6828),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_6 ));
    LocalMux I__1281 (
            .O(N__6825),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_6 ));
    IoInMux I__1280 (
            .O(N__6818),
            .I(N__6815));
    LocalMux I__1279 (
            .O(N__6815),
            .I(N__6812));
    Span12Mux_s11_v I__1278 (
            .O(N__6812),
            .I(N__6808));
    InMux I__1277 (
            .O(N__6811),
            .I(N__6805));
    Odrv12 I__1276 (
            .O(N__6808),
            .I(REGENn_c));
    LocalMux I__1275 (
            .O(N__6805),
            .I(REGENn_c));
    InMux I__1274 (
            .O(N__6800),
            .I(N__6793));
    InMux I__1273 (
            .O(N__6799),
            .I(N__6793));
    InMux I__1272 (
            .O(N__6798),
            .I(N__6790));
    LocalMux I__1271 (
            .O(N__6793),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_4 ));
    LocalMux I__1270 (
            .O(N__6790),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_4 ));
    CascadeMux I__1269 (
            .O(N__6785),
            .I(N__6781));
    InMux I__1268 (
            .O(N__6784),
            .I(N__6777));
    InMux I__1267 (
            .O(N__6781),
            .I(N__6774));
    InMux I__1266 (
            .O(N__6780),
            .I(N__6771));
    LocalMux I__1265 (
            .O(N__6777),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_3 ));
    LocalMux I__1264 (
            .O(N__6774),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_3 ));
    LocalMux I__1263 (
            .O(N__6771),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_3 ));
    InMux I__1262 (
            .O(N__6764),
            .I(N__6761));
    LocalMux I__1261 (
            .O(N__6761),
            .I(N__6757));
    InMux I__1260 (
            .O(N__6760),
            .I(N__6754));
    Span4Mux_v I__1259 (
            .O(N__6757),
            .I(N__6748));
    LocalMux I__1258 (
            .O(N__6754),
            .I(N__6748));
    InMux I__1257 (
            .O(N__6753),
            .I(N__6745));
    Odrv4 I__1256 (
            .O(N__6748),
            .I(\U712_REG_SM.DBR_SYNCZ0Z_1 ));
    LocalMux I__1255 (
            .O(N__6745),
            .I(\U712_REG_SM.DBR_SYNCZ0Z_1 ));
    CascadeMux I__1254 (
            .O(N__6740),
            .I(N__6731));
    InMux I__1253 (
            .O(N__6739),
            .I(N__6726));
    InMux I__1252 (
            .O(N__6738),
            .I(N__6721));
    InMux I__1251 (
            .O(N__6737),
            .I(N__6721));
    InMux I__1250 (
            .O(N__6736),
            .I(N__6716));
    InMux I__1249 (
            .O(N__6735),
            .I(N__6711));
    InMux I__1248 (
            .O(N__6734),
            .I(N__6711));
    InMux I__1247 (
            .O(N__6731),
            .I(N__6708));
    InMux I__1246 (
            .O(N__6730),
            .I(N__6703));
    InMux I__1245 (
            .O(N__6729),
            .I(N__6703));
    LocalMux I__1244 (
            .O(N__6726),
            .I(N__6698));
    LocalMux I__1243 (
            .O(N__6721),
            .I(N__6698));
    InMux I__1242 (
            .O(N__6720),
            .I(N__6695));
    CascadeMux I__1241 (
            .O(N__6719),
            .I(N__6689));
    LocalMux I__1240 (
            .O(N__6716),
            .I(N__6682));
    LocalMux I__1239 (
            .O(N__6711),
            .I(N__6682));
    LocalMux I__1238 (
            .O(N__6708),
            .I(N__6677));
    LocalMux I__1237 (
            .O(N__6703),
            .I(N__6677));
    Span4Mux_h I__1236 (
            .O(N__6698),
            .I(N__6672));
    LocalMux I__1235 (
            .O(N__6695),
            .I(N__6672));
    InMux I__1234 (
            .O(N__6694),
            .I(N__6665));
    InMux I__1233 (
            .O(N__6693),
            .I(N__6665));
    InMux I__1232 (
            .O(N__6692),
            .I(N__6665));
    InMux I__1231 (
            .O(N__6689),
            .I(N__6660));
    InMux I__1230 (
            .O(N__6688),
            .I(N__6660));
    InMux I__1229 (
            .O(N__6687),
            .I(N__6657));
    Odrv4 I__1228 (
            .O(N__6682),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv12 I__1227 (
            .O(N__6677),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1226 (
            .O(N__6672),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1225 (
            .O(N__6665),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1224 (
            .O(N__6660),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1223 (
            .O(N__6657),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    CascadeMux I__1222 (
            .O(N__6644),
            .I(\U712_CHIP_RAM.N_316_cascade_ ));
    InMux I__1221 (
            .O(N__6641),
            .I(N__6638));
    LocalMux I__1220 (
            .O(N__6638),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_1 ));
    InMux I__1219 (
            .O(N__6635),
            .I(N__6632));
    LocalMux I__1218 (
            .O(N__6632),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_101_i_a2_0_i_1 ));
    CascadeMux I__1217 (
            .O(N__6629),
            .I(N__6623));
    InMux I__1216 (
            .O(N__6628),
            .I(N__6614));
    CascadeMux I__1215 (
            .O(N__6627),
            .I(N__6610));
    InMux I__1214 (
            .O(N__6626),
            .I(N__6607));
    InMux I__1213 (
            .O(N__6623),
            .I(N__6603));
    InMux I__1212 (
            .O(N__6622),
            .I(N__6600));
    InMux I__1211 (
            .O(N__6621),
            .I(N__6592));
    InMux I__1210 (
            .O(N__6620),
            .I(N__6592));
    InMux I__1209 (
            .O(N__6619),
            .I(N__6592));
    InMux I__1208 (
            .O(N__6618),
            .I(N__6589));
    InMux I__1207 (
            .O(N__6617),
            .I(N__6586));
    LocalMux I__1206 (
            .O(N__6614),
            .I(N__6583));
    InMux I__1205 (
            .O(N__6613),
            .I(N__6578));
    InMux I__1204 (
            .O(N__6610),
            .I(N__6575));
    LocalMux I__1203 (
            .O(N__6607),
            .I(N__6572));
    CascadeMux I__1202 (
            .O(N__6606),
            .I(N__6568));
    LocalMux I__1201 (
            .O(N__6603),
            .I(N__6562));
    LocalMux I__1200 (
            .O(N__6600),
            .I(N__6562));
    InMux I__1199 (
            .O(N__6599),
            .I(N__6559));
    LocalMux I__1198 (
            .O(N__6592),
            .I(N__6554));
    LocalMux I__1197 (
            .O(N__6589),
            .I(N__6554));
    LocalMux I__1196 (
            .O(N__6586),
            .I(N__6551));
    Span4Mux_v I__1195 (
            .O(N__6583),
            .I(N__6548));
    InMux I__1194 (
            .O(N__6582),
            .I(N__6543));
    InMux I__1193 (
            .O(N__6581),
            .I(N__6543));
    LocalMux I__1192 (
            .O(N__6578),
            .I(N__6536));
    LocalMux I__1191 (
            .O(N__6575),
            .I(N__6536));
    Span4Mux_h I__1190 (
            .O(N__6572),
            .I(N__6536));
    InMux I__1189 (
            .O(N__6571),
            .I(N__6533));
    InMux I__1188 (
            .O(N__6568),
            .I(N__6530));
    InMux I__1187 (
            .O(N__6567),
            .I(N__6527));
    Span4Mux_v I__1186 (
            .O(N__6562),
            .I(N__6518));
    LocalMux I__1185 (
            .O(N__6559),
            .I(N__6518));
    Span4Mux_h I__1184 (
            .O(N__6554),
            .I(N__6518));
    Span4Mux_h I__1183 (
            .O(N__6551),
            .I(N__6518));
    Odrv4 I__1182 (
            .O(N__6548),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1181 (
            .O(N__6543),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1180 (
            .O(N__6536),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1179 (
            .O(N__6533),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1178 (
            .O(N__6530),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1177 (
            .O(N__6527),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1176 (
            .O(N__6518),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__1175 (
            .O(N__6503),
            .I(N__6500));
    LocalMux I__1174 (
            .O(N__6500),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_0 ));
    CascadeMux I__1173 (
            .O(N__6497),
            .I(N__6491));
    InMux I__1172 (
            .O(N__6496),
            .I(N__6482));
    InMux I__1171 (
            .O(N__6495),
            .I(N__6482));
    InMux I__1170 (
            .O(N__6494),
            .I(N__6482));
    InMux I__1169 (
            .O(N__6491),
            .I(N__6479));
    InMux I__1168 (
            .O(N__6490),
            .I(N__6476));
    CascadeMux I__1167 (
            .O(N__6489),
            .I(N__6468));
    LocalMux I__1166 (
            .O(N__6482),
            .I(N__6461));
    LocalMux I__1165 (
            .O(N__6479),
            .I(N__6461));
    LocalMux I__1164 (
            .O(N__6476),
            .I(N__6461));
    InMux I__1163 (
            .O(N__6475),
            .I(N__6456));
    InMux I__1162 (
            .O(N__6474),
            .I(N__6456));
    InMux I__1161 (
            .O(N__6473),
            .I(N__6453));
    InMux I__1160 (
            .O(N__6472),
            .I(N__6450));
    InMux I__1159 (
            .O(N__6471),
            .I(N__6447));
    InMux I__1158 (
            .O(N__6468),
            .I(N__6442));
    Span4Mux_v I__1157 (
            .O(N__6461),
            .I(N__6439));
    LocalMux I__1156 (
            .O(N__6456),
            .I(N__6430));
    LocalMux I__1155 (
            .O(N__6453),
            .I(N__6430));
    LocalMux I__1154 (
            .O(N__6450),
            .I(N__6430));
    LocalMux I__1153 (
            .O(N__6447),
            .I(N__6430));
    InMux I__1152 (
            .O(N__6446),
            .I(N__6425));
    InMux I__1151 (
            .O(N__6445),
            .I(N__6425));
    LocalMux I__1150 (
            .O(N__6442),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1149 (
            .O(N__6439),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1148 (
            .O(N__6430),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1147 (
            .O(N__6425),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    CascadeMux I__1146 (
            .O(N__6416),
            .I(N__6412));
    CascadeMux I__1145 (
            .O(N__6415),
            .I(N__6409));
    InMux I__1144 (
            .O(N__6412),
            .I(N__6398));
    InMux I__1143 (
            .O(N__6409),
            .I(N__6398));
    InMux I__1142 (
            .O(N__6408),
            .I(N__6393));
    InMux I__1141 (
            .O(N__6407),
            .I(N__6393));
    CascadeMux I__1140 (
            .O(N__6406),
            .I(N__6390));
    CascadeMux I__1139 (
            .O(N__6405),
            .I(N__6385));
    CascadeMux I__1138 (
            .O(N__6404),
            .I(N__6382));
    InMux I__1137 (
            .O(N__6403),
            .I(N__6379));
    LocalMux I__1136 (
            .O(N__6398),
            .I(N__6374));
    LocalMux I__1135 (
            .O(N__6393),
            .I(N__6374));
    InMux I__1134 (
            .O(N__6390),
            .I(N__6367));
    InMux I__1133 (
            .O(N__6389),
            .I(N__6364));
    InMux I__1132 (
            .O(N__6388),
            .I(N__6361));
    InMux I__1131 (
            .O(N__6385),
            .I(N__6355));
    InMux I__1130 (
            .O(N__6382),
            .I(N__6352));
    LocalMux I__1129 (
            .O(N__6379),
            .I(N__6349));
    Span4Mux_v I__1128 (
            .O(N__6374),
            .I(N__6346));
    InMux I__1127 (
            .O(N__6373),
            .I(N__6341));
    InMux I__1126 (
            .O(N__6372),
            .I(N__6341));
    InMux I__1125 (
            .O(N__6371),
            .I(N__6336));
    InMux I__1124 (
            .O(N__6370),
            .I(N__6336));
    LocalMux I__1123 (
            .O(N__6367),
            .I(N__6329));
    LocalMux I__1122 (
            .O(N__6364),
            .I(N__6329));
    LocalMux I__1121 (
            .O(N__6361),
            .I(N__6329));
    InMux I__1120 (
            .O(N__6360),
            .I(N__6322));
    InMux I__1119 (
            .O(N__6359),
            .I(N__6322));
    InMux I__1118 (
            .O(N__6358),
            .I(N__6322));
    LocalMux I__1117 (
            .O(N__6355),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1116 (
            .O(N__6352),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1115 (
            .O(N__6349),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1114 (
            .O(N__6346),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1113 (
            .O(N__6341),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1112 (
            .O(N__6336),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1111 (
            .O(N__6329),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1110 (
            .O(N__6322),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    InMux I__1109 (
            .O(N__6305),
            .I(N__6302));
    LocalMux I__1108 (
            .O(N__6302),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_0 ));
    InMux I__1107 (
            .O(N__6299),
            .I(N__6290));
    InMux I__1106 (
            .O(N__6298),
            .I(N__6287));
    InMux I__1105 (
            .O(N__6297),
            .I(N__6282));
    InMux I__1104 (
            .O(N__6296),
            .I(N__6282));
    InMux I__1103 (
            .O(N__6295),
            .I(N__6277));
    InMux I__1102 (
            .O(N__6294),
            .I(N__6277));
    CascadeMux I__1101 (
            .O(N__6293),
            .I(N__6273));
    LocalMux I__1100 (
            .O(N__6290),
            .I(N__6270));
    LocalMux I__1099 (
            .O(N__6287),
            .I(N__6259));
    LocalMux I__1098 (
            .O(N__6282),
            .I(N__6259));
    LocalMux I__1097 (
            .O(N__6277),
            .I(N__6259));
    InMux I__1096 (
            .O(N__6276),
            .I(N__6256));
    InMux I__1095 (
            .O(N__6273),
            .I(N__6253));
    Span4Mux_h I__1094 (
            .O(N__6270),
            .I(N__6250));
    InMux I__1093 (
            .O(N__6269),
            .I(N__6245));
    InMux I__1092 (
            .O(N__6268),
            .I(N__6245));
    InMux I__1091 (
            .O(N__6267),
            .I(N__6240));
    InMux I__1090 (
            .O(N__6266),
            .I(N__6240));
    Sp12to4 I__1089 (
            .O(N__6259),
            .I(N__6235));
    LocalMux I__1088 (
            .O(N__6256),
            .I(N__6235));
    LocalMux I__1087 (
            .O(N__6253),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1086 (
            .O(N__6250),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1085 (
            .O(N__6245),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1084 (
            .O(N__6240),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv12 I__1083 (
            .O(N__6235),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    InMux I__1082 (
            .O(N__6224),
            .I(N__6218));
    InMux I__1081 (
            .O(N__6223),
            .I(N__6215));
    CascadeMux I__1080 (
            .O(N__6222),
            .I(N__6208));
    InMux I__1079 (
            .O(N__6221),
            .I(N__6204));
    LocalMux I__1078 (
            .O(N__6218),
            .I(N__6197));
    LocalMux I__1077 (
            .O(N__6215),
            .I(N__6189));
    InMux I__1076 (
            .O(N__6214),
            .I(N__6184));
    InMux I__1075 (
            .O(N__6213),
            .I(N__6184));
    InMux I__1074 (
            .O(N__6212),
            .I(N__6181));
    InMux I__1073 (
            .O(N__6211),
            .I(N__6176));
    InMux I__1072 (
            .O(N__6208),
            .I(N__6176));
    InMux I__1071 (
            .O(N__6207),
            .I(N__6173));
    LocalMux I__1070 (
            .O(N__6204),
            .I(N__6170));
    InMux I__1069 (
            .O(N__6203),
            .I(N__6165));
    InMux I__1068 (
            .O(N__6202),
            .I(N__6165));
    InMux I__1067 (
            .O(N__6201),
            .I(N__6162));
    InMux I__1066 (
            .O(N__6200),
            .I(N__6157));
    Span4Mux_v I__1065 (
            .O(N__6197),
            .I(N__6154));
    InMux I__1064 (
            .O(N__6196),
            .I(N__6147));
    InMux I__1063 (
            .O(N__6195),
            .I(N__6147));
    InMux I__1062 (
            .O(N__6194),
            .I(N__6147));
    InMux I__1061 (
            .O(N__6193),
            .I(N__6142));
    InMux I__1060 (
            .O(N__6192),
            .I(N__6142));
    Span4Mux_v I__1059 (
            .O(N__6189),
            .I(N__6133));
    LocalMux I__1058 (
            .O(N__6184),
            .I(N__6133));
    LocalMux I__1057 (
            .O(N__6181),
            .I(N__6133));
    LocalMux I__1056 (
            .O(N__6176),
            .I(N__6133));
    LocalMux I__1055 (
            .O(N__6173),
            .I(N__6124));
    Span4Mux_h I__1054 (
            .O(N__6170),
            .I(N__6124));
    LocalMux I__1053 (
            .O(N__6165),
            .I(N__6124));
    LocalMux I__1052 (
            .O(N__6162),
            .I(N__6124));
    InMux I__1051 (
            .O(N__6161),
            .I(N__6121));
    InMux I__1050 (
            .O(N__6160),
            .I(N__6118));
    LocalMux I__1049 (
            .O(N__6157),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1048 (
            .O(N__6154),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1047 (
            .O(N__6147),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1046 (
            .O(N__6142),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1045 (
            .O(N__6133),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1044 (
            .O(N__6124),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1043 (
            .O(N__6121),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1042 (
            .O(N__6118),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    CascadeMux I__1041 (
            .O(N__6101),
            .I(N__6098));
    InMux I__1040 (
            .O(N__6098),
            .I(N__6090));
    InMux I__1039 (
            .O(N__6097),
            .I(N__6087));
    InMux I__1038 (
            .O(N__6096),
            .I(N__6084));
    CascadeMux I__1037 (
            .O(N__6095),
            .I(N__6081));
    CascadeMux I__1036 (
            .O(N__6094),
            .I(N__6078));
    InMux I__1035 (
            .O(N__6093),
            .I(N__6073));
    LocalMux I__1034 (
            .O(N__6090),
            .I(N__6070));
    LocalMux I__1033 (
            .O(N__6087),
            .I(N__6067));
    LocalMux I__1032 (
            .O(N__6084),
            .I(N__6064));
    InMux I__1031 (
            .O(N__6081),
            .I(N__6057));
    InMux I__1030 (
            .O(N__6078),
            .I(N__6057));
    InMux I__1029 (
            .O(N__6077),
            .I(N__6057));
    InMux I__1028 (
            .O(N__6076),
            .I(N__6054));
    LocalMux I__1027 (
            .O(N__6073),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    Odrv4 I__1026 (
            .O(N__6070),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    Odrv4 I__1025 (
            .O(N__6067),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    Odrv4 I__1024 (
            .O(N__6064),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    LocalMux I__1023 (
            .O(N__6057),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    LocalMux I__1022 (
            .O(N__6054),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    InMux I__1021 (
            .O(N__6041),
            .I(N__6038));
    LocalMux I__1020 (
            .O(N__6038),
            .I(\U712_CHIP_RAM.N_109_i ));
    InMux I__1019 (
            .O(N__6035),
            .I(N__6032));
    LocalMux I__1018 (
            .O(N__6032),
            .I(N__6029));
    Span12Mux_s11_v I__1017 (
            .O(N__6029),
            .I(N__6026));
    Span12Mux_h I__1016 (
            .O(N__6026),
            .I(N__6023));
    Odrv12 I__1015 (
            .O(N__6023),
            .I(A_c_10));
    InMux I__1014 (
            .O(N__6020),
            .I(N__6017));
    LocalMux I__1013 (
            .O(N__6017),
            .I(N__6014));
    Span12Mux_v I__1012 (
            .O(N__6014),
            .I(N__6011));
    Span12Mux_h I__1011 (
            .O(N__6011),
            .I(N__6008));
    Odrv12 I__1010 (
            .O(N__6008),
            .I(A_c_16));
    InMux I__1009 (
            .O(N__6005),
            .I(N__6002));
    LocalMux I__1008 (
            .O(N__6002),
            .I(N__5999));
    Span12Mux_v I__1007 (
            .O(N__5999),
            .I(N__5996));
    Span12Mux_h I__1006 (
            .O(N__5996),
            .I(N__5993));
    Odrv12 I__1005 (
            .O(N__5993),
            .I(A_c_18));
    InMux I__1004 (
            .O(N__5990),
            .I(N__5987));
    LocalMux I__1003 (
            .O(N__5987),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ));
    CascadeMux I__1002 (
            .O(N__5984),
            .I(\U712_CHIP_RAM.N_411_cascade_ ));
    InMux I__1001 (
            .O(N__5981),
            .I(N__5978));
    LocalMux I__1000 (
            .O(N__5978),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_1_0 ));
    CascadeMux I__999 (
            .O(N__5975),
            .I(N__5971));
    CascadeMux I__998 (
            .O(N__5974),
            .I(N__5967));
    InMux I__997 (
            .O(N__5971),
            .I(N__5960));
    InMux I__996 (
            .O(N__5970),
            .I(N__5960));
    InMux I__995 (
            .O(N__5967),
            .I(N__5960));
    LocalMux I__994 (
            .O(N__5960),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_o3_0_0 ));
    CascadeMux I__993 (
            .O(N__5957),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_1_0_cascade_ ));
    InMux I__992 (
            .O(N__5954),
            .I(N__5948));
    InMux I__991 (
            .O(N__5953),
            .I(N__5941));
    InMux I__990 (
            .O(N__5952),
            .I(N__5941));
    InMux I__989 (
            .O(N__5951),
            .I(N__5941));
    LocalMux I__988 (
            .O(N__5948),
            .I(\U712_CHIP_RAM.N_294 ));
    LocalMux I__987 (
            .O(N__5941),
            .I(\U712_CHIP_RAM.N_294 ));
    CEMux I__986 (
            .O(N__5936),
            .I(N__5932));
    CEMux I__985 (
            .O(N__5935),
            .I(N__5929));
    LocalMux I__984 (
            .O(N__5932),
            .I(N__5926));
    LocalMux I__983 (
            .O(N__5929),
            .I(N__5923));
    Span4Mux_v I__982 (
            .O(N__5926),
            .I(N__5920));
    Span4Mux_h I__981 (
            .O(N__5923),
            .I(N__5917));
    Odrv4 I__980 (
            .O(N__5920),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ));
    Odrv4 I__979 (
            .O(N__5917),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ));
    InMux I__978 (
            .O(N__5912),
            .I(N__5909));
    LocalMux I__977 (
            .O(N__5909),
            .I(N__5901));
    InMux I__976 (
            .O(N__5908),
            .I(N__5897));
    CascadeMux I__975 (
            .O(N__5907),
            .I(N__5894));
    InMux I__974 (
            .O(N__5906),
            .I(N__5888));
    InMux I__973 (
            .O(N__5905),
            .I(N__5885));
    InMux I__972 (
            .O(N__5904),
            .I(N__5882));
    Span4Mux_h I__971 (
            .O(N__5901),
            .I(N__5879));
    InMux I__970 (
            .O(N__5900),
            .I(N__5876));
    LocalMux I__969 (
            .O(N__5897),
            .I(N__5873));
    InMux I__968 (
            .O(N__5894),
            .I(N__5870));
    InMux I__967 (
            .O(N__5893),
            .I(N__5863));
    InMux I__966 (
            .O(N__5892),
            .I(N__5863));
    InMux I__965 (
            .O(N__5891),
            .I(N__5863));
    LocalMux I__964 (
            .O(N__5888),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__963 (
            .O(N__5885),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__962 (
            .O(N__5882),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    Odrv4 I__961 (
            .O(N__5879),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__960 (
            .O(N__5876),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    Odrv4 I__959 (
            .O(N__5873),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__958 (
            .O(N__5870),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__957 (
            .O(N__5863),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__956 (
            .O(N__5846),
            .I(N__5843));
    LocalMux I__955 (
            .O(N__5843),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_1_0_0 ));
    CascadeMux I__954 (
            .O(N__5840),
            .I(N__5836));
    CascadeMux I__953 (
            .O(N__5839),
            .I(N__5829));
    InMux I__952 (
            .O(N__5836),
            .I(N__5826));
    InMux I__951 (
            .O(N__5835),
            .I(N__5823));
    InMux I__950 (
            .O(N__5834),
            .I(N__5818));
    InMux I__949 (
            .O(N__5833),
            .I(N__5818));
    InMux I__948 (
            .O(N__5832),
            .I(N__5813));
    InMux I__947 (
            .O(N__5829),
            .I(N__5813));
    LocalMux I__946 (
            .O(N__5826),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__945 (
            .O(N__5823),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__944 (
            .O(N__5818),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__943 (
            .O(N__5813),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    CascadeMux I__942 (
            .O(N__5804),
            .I(N__5801));
    InMux I__941 (
            .O(N__5801),
            .I(N__5797));
    InMux I__940 (
            .O(N__5800),
            .I(N__5794));
    LocalMux I__939 (
            .O(N__5797),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    LocalMux I__938 (
            .O(N__5794),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    InMux I__937 (
            .O(N__5789),
            .I(N__5785));
    InMux I__936 (
            .O(N__5788),
            .I(N__5781));
    LocalMux I__935 (
            .O(N__5785),
            .I(N__5778));
    InMux I__934 (
            .O(N__5784),
            .I(N__5775));
    LocalMux I__933 (
            .O(N__5781),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    Odrv4 I__932 (
            .O(N__5778),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__931 (
            .O(N__5775),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    InMux I__930 (
            .O(N__5768),
            .I(N__5765));
    LocalMux I__929 (
            .O(N__5765),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_5 ));
    InMux I__928 (
            .O(N__5762),
            .I(N__5759));
    LocalMux I__927 (
            .O(N__5759),
            .I(N__5756));
    Span4Mux_v I__926 (
            .O(N__5756),
            .I(N__5752));
    InMux I__925 (
            .O(N__5755),
            .I(N__5749));
    Odrv4 I__924 (
            .O(N__5752),
            .I(LATCH_REG));
    LocalMux I__923 (
            .O(N__5749),
            .I(LATCH_REG));
    InMux I__922 (
            .O(N__5744),
            .I(N__5741));
    LocalMux I__921 (
            .O(N__5741),
            .I(N__5738));
    Span12Mux_v I__920 (
            .O(N__5738),
            .I(N__5734));
    InMux I__919 (
            .O(N__5737),
            .I(N__5731));
    Odrv12 I__918 (
            .O(N__5734),
            .I(REG_CPU_CYCLE));
    LocalMux I__917 (
            .O(N__5731),
            .I(REG_CPU_CYCLE));
    CascadeMux I__916 (
            .O(N__5726),
            .I(\U712_REG_SM.STATE_COUNTERc_0_cascade_ ));
    InMux I__915 (
            .O(N__5723),
            .I(N__5720));
    LocalMux I__914 (
            .O(N__5720),
            .I(\U712_REG_SM.REG_CPU_CYCLE_e_1 ));
    InMux I__913 (
            .O(N__5717),
            .I(N__5714));
    LocalMux I__912 (
            .O(N__5714),
            .I(N__5711));
    Span12Mux_v I__911 (
            .O(N__5711),
            .I(N__5708));
    Span12Mux_h I__910 (
            .O(N__5708),
            .I(N__5705));
    Span12Mux_v I__909 (
            .O(N__5705),
            .I(N__5702));
    Odrv12 I__908 (
            .O(N__5702),
            .I(A_c_3));
    InMux I__907 (
            .O(N__5699),
            .I(N__5693));
    InMux I__906 (
            .O(N__5698),
            .I(N__5693));
    LocalMux I__905 (
            .O(N__5693),
            .I(N__5690));
    Odrv4 I__904 (
            .O(N__5690),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_0_2 ));
    CascadeMux I__903 (
            .O(N__5687),
            .I(\U712_CHIP_RAM.N_421_cascade_ ));
    CEMux I__902 (
            .O(N__5684),
            .I(N__5681));
    LocalMux I__901 (
            .O(N__5681),
            .I(N__5677));
    CEMux I__900 (
            .O(N__5680),
            .I(N__5674));
    Span4Mux_h I__899 (
            .O(N__5677),
            .I(N__5671));
    LocalMux I__898 (
            .O(N__5674),
            .I(N__5668));
    Odrv4 I__897 (
            .O(N__5671),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    Odrv12 I__896 (
            .O(N__5668),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    InMux I__895 (
            .O(N__5663),
            .I(N__5659));
    InMux I__894 (
            .O(N__5662),
            .I(N__5656));
    LocalMux I__893 (
            .O(N__5659),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    LocalMux I__892 (
            .O(N__5656),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    InMux I__891 (
            .O(N__5651),
            .I(N__5648));
    LocalMux I__890 (
            .O(N__5648),
            .I(\U712_CHIP_RAM.N_18 ));
    CEMux I__889 (
            .O(N__5645),
            .I(N__5642));
    LocalMux I__888 (
            .O(N__5642),
            .I(\U712_CHIP_RAM.N_18_0 ));
    InMux I__887 (
            .O(N__5639),
            .I(N__5635));
    InMux I__886 (
            .O(N__5638),
            .I(N__5632));
    LocalMux I__885 (
            .O(N__5635),
            .I(N__5629));
    LocalMux I__884 (
            .O(N__5632),
            .I(N__5626));
    Span4Mux_h I__883 (
            .O(N__5629),
            .I(N__5623));
    Odrv4 I__882 (
            .O(N__5626),
            .I(\U712_CHIP_RAM.N_113 ));
    Odrv4 I__881 (
            .O(N__5623),
            .I(\U712_CHIP_RAM.N_113 ));
    CascadeMux I__880 (
            .O(N__5618),
            .I(N__5614));
    InMux I__879 (
            .O(N__5617),
            .I(N__5611));
    InMux I__878 (
            .O(N__5614),
            .I(N__5608));
    LocalMux I__877 (
            .O(N__5611),
            .I(N__5604));
    LocalMux I__876 (
            .O(N__5608),
            .I(N__5601));
    InMux I__875 (
            .O(N__5607),
            .I(N__5597));
    Span4Mux_v I__874 (
            .O(N__5604),
            .I(N__5592));
    Span4Mux_v I__873 (
            .O(N__5601),
            .I(N__5592));
    InMux I__872 (
            .O(N__5600),
            .I(N__5589));
    LocalMux I__871 (
            .O(N__5597),
            .I(\U712_CHIP_RAM.N_413 ));
    Odrv4 I__870 (
            .O(N__5592),
            .I(\U712_CHIP_RAM.N_413 ));
    LocalMux I__869 (
            .O(N__5589),
            .I(\U712_CHIP_RAM.N_413 ));
    IoInMux I__868 (
            .O(N__5582),
            .I(N__5579));
    LocalMux I__867 (
            .O(N__5579),
            .I(N__5576));
    IoSpan4Mux I__866 (
            .O(N__5576),
            .I(N__5573));
    Sp12to4 I__865 (
            .O(N__5573),
            .I(N__5570));
    Span12Mux_s7_h I__864 (
            .O(N__5570),
            .I(N__5567));
    Span12Mux_h I__863 (
            .O(N__5567),
            .I(N__5563));
    InMux I__862 (
            .O(N__5566),
            .I(N__5560));
    Odrv12 I__861 (
            .O(N__5563),
            .I(CLK_EN_c));
    LocalMux I__860 (
            .O(N__5560),
            .I(CLK_EN_c));
    InMux I__859 (
            .O(N__5555),
            .I(N__5552));
    LocalMux I__858 (
            .O(N__5552),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa ));
    CascadeMux I__857 (
            .O(N__5549),
            .I(N__5546));
    InMux I__856 (
            .O(N__5546),
            .I(N__5542));
    InMux I__855 (
            .O(N__5545),
            .I(N__5539));
    LocalMux I__854 (
            .O(N__5542),
            .I(\U712_CHIP_RAM.N_342 ));
    LocalMux I__853 (
            .O(N__5539),
            .I(\U712_CHIP_RAM.N_342 ));
    InMux I__852 (
            .O(N__5534),
            .I(N__5531));
    LocalMux I__851 (
            .O(N__5531),
            .I(N__5528));
    Odrv4 I__850 (
            .O(N__5528),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0 ));
    InMux I__849 (
            .O(N__5525),
            .I(N__5521));
    InMux I__848 (
            .O(N__5524),
            .I(N__5518));
    LocalMux I__847 (
            .O(N__5521),
            .I(N__5515));
    LocalMux I__846 (
            .O(N__5518),
            .I(N__5512));
    Span4Mux_v I__845 (
            .O(N__5515),
            .I(N__5509));
    Span4Mux_v I__844 (
            .O(N__5512),
            .I(N__5506));
    Sp12to4 I__843 (
            .O(N__5509),
            .I(N__5501));
    Sp12to4 I__842 (
            .O(N__5506),
            .I(N__5501));
    Span12Mux_h I__841 (
            .O(N__5501),
            .I(N__5498));
    Span12Mux_v I__840 (
            .O(N__5498),
            .I(N__5495));
    Odrv12 I__839 (
            .O(N__5495),
            .I(AWEn_c));
    IoInMux I__838 (
            .O(N__5492),
            .I(N__5489));
    LocalMux I__837 (
            .O(N__5489),
            .I(N__5486));
    Span4Mux_s3_v I__836 (
            .O(N__5486),
            .I(N__5483));
    Span4Mux_v I__835 (
            .O(N__5483),
            .I(N__5480));
    Span4Mux_v I__834 (
            .O(N__5480),
            .I(N__5477));
    Span4Mux_v I__833 (
            .O(N__5477),
            .I(N__5473));
    InMux I__832 (
            .O(N__5476),
            .I(N__5470));
    Odrv4 I__831 (
            .O(N__5473),
            .I(DBDIR_c));
    LocalMux I__830 (
            .O(N__5470),
            .I(DBDIR_c));
    InMux I__829 (
            .O(N__5465),
            .I(N__5462));
    LocalMux I__828 (
            .O(N__5462),
            .I(N__5458));
    InMux I__827 (
            .O(N__5461),
            .I(N__5455));
    Odrv4 I__826 (
            .O(N__5458),
            .I(DBRn_c_i));
    LocalMux I__825 (
            .O(N__5455),
            .I(DBRn_c_i));
    IoInMux I__824 (
            .O(N__5450),
            .I(N__5447));
    LocalMux I__823 (
            .O(N__5447),
            .I(N__5444));
    Span12Mux_s4_h I__822 (
            .O(N__5444),
            .I(N__5441));
    Odrv12 I__821 (
            .O(N__5441),
            .I(DBRn_c_i_0));
    InMux I__820 (
            .O(N__5438),
            .I(N__5435));
    LocalMux I__819 (
            .O(N__5435),
            .I(N__5432));
    Span4Mux_v I__818 (
            .O(N__5432),
            .I(N__5429));
    Sp12to4 I__817 (
            .O(N__5429),
            .I(N__5426));
    Odrv12 I__816 (
            .O(N__5426),
            .I(A_c_13));
    InMux I__815 (
            .O(N__5423),
            .I(N__5420));
    LocalMux I__814 (
            .O(N__5420),
            .I(N__5417));
    Span4Mux_v I__813 (
            .O(N__5417),
            .I(N__5414));
    Span4Mux_h I__812 (
            .O(N__5414),
            .I(N__5411));
    Sp12to4 I__811 (
            .O(N__5411),
            .I(N__5408));
    Odrv12 I__810 (
            .O(N__5408),
            .I(A_c_12));
    InMux I__809 (
            .O(N__5405),
            .I(N__5402));
    LocalMux I__808 (
            .O(N__5402),
            .I(N__5399));
    Span4Mux_v I__807 (
            .O(N__5399),
            .I(N__5396));
    Span4Mux_v I__806 (
            .O(N__5396),
            .I(N__5393));
    Sp12to4 I__805 (
            .O(N__5393),
            .I(N__5390));
    Odrv12 I__804 (
            .O(N__5390),
            .I(A_c_5));
    InMux I__803 (
            .O(N__5387),
            .I(N__5384));
    LocalMux I__802 (
            .O(N__5384),
            .I(N__5381));
    Span4Mux_v I__801 (
            .O(N__5381),
            .I(N__5378));
    Span4Mux_v I__800 (
            .O(N__5378),
            .I(N__5375));
    Sp12to4 I__799 (
            .O(N__5375),
            .I(N__5372));
    Odrv12 I__798 (
            .O(N__5372),
            .I(A_c_15));
    InMux I__797 (
            .O(N__5369),
            .I(N__5366));
    LocalMux I__796 (
            .O(N__5366),
            .I(N__5363));
    Span4Mux_h I__795 (
            .O(N__5363),
            .I(N__5360));
    Span4Mux_v I__794 (
            .O(N__5360),
            .I(N__5357));
    Sp12to4 I__793 (
            .O(N__5357),
            .I(N__5354));
    Odrv12 I__792 (
            .O(N__5354),
            .I(A_c_8));
    InMux I__791 (
            .O(N__5351),
            .I(N__5347));
    InMux I__790 (
            .O(N__5350),
            .I(N__5344));
    LocalMux I__789 (
            .O(N__5347),
            .I(N__5341));
    LocalMux I__788 (
            .O(N__5344),
            .I(N__5336));
    Span4Mux_v I__787 (
            .O(N__5341),
            .I(N__5333));
    InMux I__786 (
            .O(N__5340),
            .I(N__5330));
    InMux I__785 (
            .O(N__5339),
            .I(N__5327));
    Odrv4 I__784 (
            .O(N__5336),
            .I(\U712_CHIP_RAM.N_261 ));
    Odrv4 I__783 (
            .O(N__5333),
            .I(\U712_CHIP_RAM.N_261 ));
    LocalMux I__782 (
            .O(N__5330),
            .I(\U712_CHIP_RAM.N_261 ));
    LocalMux I__781 (
            .O(N__5327),
            .I(\U712_CHIP_RAM.N_261 ));
    InMux I__780 (
            .O(N__5318),
            .I(N__5315));
    LocalMux I__779 (
            .O(N__5315),
            .I(N__5312));
    Span4Mux_v I__778 (
            .O(N__5312),
            .I(N__5309));
    Sp12to4 I__777 (
            .O(N__5309),
            .I(N__5306));
    Odrv12 I__776 (
            .O(N__5306),
            .I(A_c_11));
    InMux I__775 (
            .O(N__5303),
            .I(N__5300));
    LocalMux I__774 (
            .O(N__5300),
            .I(N__5297));
    Sp12to4 I__773 (
            .O(N__5297),
            .I(N__5294));
    Span12Mux_v I__772 (
            .O(N__5294),
            .I(N__5291));
    Span12Mux_h I__771 (
            .O(N__5291),
            .I(N__5288));
    Odrv12 I__770 (
            .O(N__5288),
            .I(A_c_4));
    InMux I__769 (
            .O(N__5285),
            .I(N__5282));
    LocalMux I__768 (
            .O(N__5282),
            .I(\U712_CHIP_RAM.N_312 ));
    InMux I__767 (
            .O(N__5279),
            .I(N__5276));
    LocalMux I__766 (
            .O(N__5276),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_63_i_a2_0_i_0 ));
    CascadeMux I__765 (
            .O(N__5273),
            .I(N__5270));
    InMux I__764 (
            .O(N__5270),
            .I(N__5267));
    LocalMux I__763 (
            .O(N__5267),
            .I(N__5264));
    Span4Mux_h I__762 (
            .O(N__5264),
            .I(N__5261));
    Odrv4 I__761 (
            .O(N__5261),
            .I(\U712_CHIP_RAM.N_314 ));
    InMux I__760 (
            .O(N__5258),
            .I(N__5255));
    LocalMux I__759 (
            .O(N__5255),
            .I(N__5251));
    InMux I__758 (
            .O(N__5254),
            .I(N__5248));
    Span4Mux_h I__757 (
            .O(N__5251),
            .I(N__5245));
    LocalMux I__756 (
            .O(N__5248),
            .I(\U712_CHIP_RAM.N_459 ));
    Odrv4 I__755 (
            .O(N__5245),
            .I(\U712_CHIP_RAM.N_459 ));
    InMux I__754 (
            .O(N__5240),
            .I(N__5237));
    LocalMux I__753 (
            .O(N__5237),
            .I(N__5232));
    InMux I__752 (
            .O(N__5236),
            .I(N__5227));
    InMux I__751 (
            .O(N__5235),
            .I(N__5227));
    Span4Mux_h I__750 (
            .O(N__5232),
            .I(N__5224));
    LocalMux I__749 (
            .O(N__5227),
            .I(\U712_CHIP_RAM.N_449 ));
    Odrv4 I__748 (
            .O(N__5224),
            .I(\U712_CHIP_RAM.N_449 ));
    CascadeMux I__747 (
            .O(N__5219),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i_1_cascade_ ));
    InMux I__746 (
            .O(N__5216),
            .I(N__5211));
    CascadeMux I__745 (
            .O(N__5215),
            .I(N__5201));
    InMux I__744 (
            .O(N__5214),
            .I(N__5197));
    LocalMux I__743 (
            .O(N__5211),
            .I(N__5194));
    InMux I__742 (
            .O(N__5210),
            .I(N__5189));
    InMux I__741 (
            .O(N__5209),
            .I(N__5189));
    InMux I__740 (
            .O(N__5208),
            .I(N__5178));
    InMux I__739 (
            .O(N__5207),
            .I(N__5178));
    InMux I__738 (
            .O(N__5206),
            .I(N__5171));
    InMux I__737 (
            .O(N__5205),
            .I(N__5171));
    InMux I__736 (
            .O(N__5204),
            .I(N__5171));
    InMux I__735 (
            .O(N__5201),
            .I(N__5164));
    InMux I__734 (
            .O(N__5200),
            .I(N__5164));
    LocalMux I__733 (
            .O(N__5197),
            .I(N__5161));
    Span4Mux_h I__732 (
            .O(N__5194),
            .I(N__5156));
    LocalMux I__731 (
            .O(N__5189),
            .I(N__5156));
    InMux I__730 (
            .O(N__5188),
            .I(N__5153));
    InMux I__729 (
            .O(N__5187),
            .I(N__5144));
    InMux I__728 (
            .O(N__5186),
            .I(N__5144));
    InMux I__727 (
            .O(N__5185),
            .I(N__5144));
    InMux I__726 (
            .O(N__5184),
            .I(N__5144));
    InMux I__725 (
            .O(N__5183),
            .I(N__5141));
    LocalMux I__724 (
            .O(N__5178),
            .I(N__5138));
    LocalMux I__723 (
            .O(N__5171),
            .I(N__5135));
    InMux I__722 (
            .O(N__5170),
            .I(N__5130));
    InMux I__721 (
            .O(N__5169),
            .I(N__5130));
    LocalMux I__720 (
            .O(N__5164),
            .I(N__5126));
    Span4Mux_v I__719 (
            .O(N__5161),
            .I(N__5121));
    Span4Mux_v I__718 (
            .O(N__5156),
            .I(N__5121));
    LocalMux I__717 (
            .O(N__5153),
            .I(N__5114));
    LocalMux I__716 (
            .O(N__5144),
            .I(N__5114));
    LocalMux I__715 (
            .O(N__5141),
            .I(N__5114));
    Span4Mux_v I__714 (
            .O(N__5138),
            .I(N__5107));
    Span4Mux_v I__713 (
            .O(N__5135),
            .I(N__5107));
    LocalMux I__712 (
            .O(N__5130),
            .I(N__5107));
    InMux I__711 (
            .O(N__5129),
            .I(N__5104));
    Span12Mux_v I__710 (
            .O(N__5126),
            .I(N__5093));
    Sp12to4 I__709 (
            .O(N__5121),
            .I(N__5093));
    Span12Mux_v I__708 (
            .O(N__5114),
            .I(N__5093));
    Sp12to4 I__707 (
            .O(N__5107),
            .I(N__5093));
    LocalMux I__706 (
            .O(N__5104),
            .I(N__5093));
    Span12Mux_h I__705 (
            .O(N__5093),
            .I(N__5090));
    Odrv12 I__704 (
            .O(N__5090),
            .I(RESETn_c));
    InMux I__703 (
            .O(N__5087),
            .I(N__5078));
    InMux I__702 (
            .O(N__5086),
            .I(N__5078));
    InMux I__701 (
            .O(N__5085),
            .I(N__5078));
    LocalMux I__700 (
            .O(N__5078),
            .I(N__5074));
    InMux I__699 (
            .O(N__5077),
            .I(N__5071));
    Odrv4 I__698 (
            .O(N__5074),
            .I(\U712_CHIP_RAM.N_421 ));
    LocalMux I__697 (
            .O(N__5071),
            .I(\U712_CHIP_RAM.N_421 ));
    CascadeMux I__696 (
            .O(N__5066),
            .I(\U712_CYCLE_TERM.N_286_i_0_en_cascade_ ));
    IoInMux I__695 (
            .O(N__5063),
            .I(N__5060));
    LocalMux I__694 (
            .O(N__5060),
            .I(N__5057));
    Span12Mux_s1_v I__693 (
            .O(N__5057),
            .I(N__5054));
    Span12Mux_v I__692 (
            .O(N__5054),
            .I(N__5050));
    InMux I__691 (
            .O(N__5053),
            .I(N__5047));
    Odrv12 I__690 (
            .O(N__5050),
            .I(RESETn_c_i));
    LocalMux I__689 (
            .O(N__5047),
            .I(RESETn_c_i));
    CascadeMux I__688 (
            .O(N__5042),
            .I(N__5038));
    InMux I__687 (
            .O(N__5041),
            .I(N__5032));
    InMux I__686 (
            .O(N__5038),
            .I(N__5029));
    InMux I__685 (
            .O(N__5037),
            .I(N__5022));
    InMux I__684 (
            .O(N__5036),
            .I(N__5022));
    InMux I__683 (
            .O(N__5035),
            .I(N__5022));
    LocalMux I__682 (
            .O(N__5032),
            .I(N__5019));
    LocalMux I__681 (
            .O(N__5029),
            .I(N__5016));
    LocalMux I__680 (
            .O(N__5022),
            .I(N__5013));
    Odrv4 I__679 (
            .O(N__5019),
            .I(CPU_TACK));
    Odrv12 I__678 (
            .O(N__5016),
            .I(CPU_TACK));
    Odrv4 I__677 (
            .O(N__5013),
            .I(CPU_TACK));
    CEMux I__676 (
            .O(N__5006),
            .I(N__5003));
    LocalMux I__675 (
            .O(N__5003),
            .I(N__5000));
    Odrv4 I__674 (
            .O(N__5000),
            .I(\U712_CYCLE_TERM.N_286_i_0_en_0 ));
    InMux I__673 (
            .O(N__4997),
            .I(N__4993));
    InMux I__672 (
            .O(N__4996),
            .I(N__4989));
    LocalMux I__671 (
            .O(N__4993),
            .I(N__4986));
    InMux I__670 (
            .O(N__4992),
            .I(N__4983));
    LocalMux I__669 (
            .O(N__4989),
            .I(N__4980));
    Span4Mux_v I__668 (
            .O(N__4986),
            .I(N__4975));
    LocalMux I__667 (
            .O(N__4983),
            .I(N__4975));
    Span4Mux_v I__666 (
            .O(N__4980),
            .I(N__4972));
    Span4Mux_v I__665 (
            .O(N__4975),
            .I(N__4969));
    Span4Mux_h I__664 (
            .O(N__4972),
            .I(N__4966));
    Sp12to4 I__663 (
            .O(N__4969),
            .I(N__4963));
    Sp12to4 I__662 (
            .O(N__4966),
            .I(N__4958));
    Span12Mux_h I__661 (
            .O(N__4963),
            .I(N__4958));
    Odrv12 I__660 (
            .O(N__4958),
            .I(DBRn_c));
    InMux I__659 (
            .O(N__4955),
            .I(N__4952));
    LocalMux I__658 (
            .O(N__4952),
            .I(\U712_REG_SM.DBR_SYNCZ0Z_0 ));
    InMux I__657 (
            .O(N__4949),
            .I(N__4946));
    LocalMux I__656 (
            .O(N__4946),
            .I(N__4943));
    Odrv4 I__655 (
            .O(N__4943),
            .I(TACK_EN_i_ess));
    IoInMux I__654 (
            .O(N__4940),
            .I(N__4937));
    LocalMux I__653 (
            .O(N__4937),
            .I(N__4934));
    IoSpan4Mux I__652 (
            .O(N__4934),
            .I(N__4931));
    Span4Mux_s3_h I__651 (
            .O(N__4931),
            .I(N__4928));
    Span4Mux_h I__650 (
            .O(N__4928),
            .I(N__4925));
    Span4Mux_h I__649 (
            .O(N__4925),
            .I(N__4922));
    Odrv4 I__648 (
            .O(N__4922),
            .I(N_977_i));
    IoInMux I__647 (
            .O(N__4919),
            .I(N__4916));
    LocalMux I__646 (
            .O(N__4916),
            .I(N__4913));
    Span4Mux_s2_v I__645 (
            .O(N__4913),
            .I(N__4910));
    Span4Mux_v I__644 (
            .O(N__4910),
            .I(N__4907));
    Span4Mux_v I__643 (
            .O(N__4907),
            .I(N__4904));
    Odrv4 I__642 (
            .O(N__4904),
            .I(VBENn_c));
    IoInMux I__641 (
            .O(N__4901),
            .I(N__4898));
    LocalMux I__640 (
            .O(N__4898),
            .I(N__4895));
    Span4Mux_s2_v I__639 (
            .O(N__4895),
            .I(N__4892));
    Span4Mux_v I__638 (
            .O(N__4892),
            .I(N__4888));
    InMux I__637 (
            .O(N__4891),
            .I(N__4885));
    Span4Mux_v I__636 (
            .O(N__4888),
            .I(N__4882));
    LocalMux I__635 (
            .O(N__4885),
            .I(N__4879));
    Sp12to4 I__634 (
            .O(N__4882),
            .I(N__4876));
    Span4Mux_v I__633 (
            .O(N__4879),
            .I(N__4873));
    Odrv12 I__632 (
            .O(N__4876),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__631 (
            .O(N__4873),
            .I(CONSTANT_ONE_NET));
    InMux I__630 (
            .O(N__4868),
            .I(N__4865));
    LocalMux I__629 (
            .O(N__4865),
            .I(N__4862));
    Sp12to4 I__628 (
            .O(N__4862),
            .I(N__4859));
    Span12Mux_v I__627 (
            .O(N__4859),
            .I(N__4856));
    Span12Mux_h I__626 (
            .O(N__4856),
            .I(N__4853));
    Odrv12 I__625 (
            .O(N__4853),
            .I(A_c_6));
    InMux I__624 (
            .O(N__4850),
            .I(N__4847));
    LocalMux I__623 (
            .O(N__4847),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    InMux I__622 (
            .O(N__4844),
            .I(N__4841));
    LocalMux I__621 (
            .O(N__4841),
            .I(N__4838));
    Span4Mux_v I__620 (
            .O(N__4838),
            .I(N__4835));
    Odrv4 I__619 (
            .O(N__4835),
            .I(\U712_CHIP_RAM.DMA_CYCLE_START_RNOZ0Z_0 ));
    InMux I__618 (
            .O(N__4832),
            .I(N__4828));
    InMux I__617 (
            .O(N__4831),
            .I(N__4825));
    LocalMux I__616 (
            .O(N__4828),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    LocalMux I__615 (
            .O(N__4825),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    CascadeMux I__614 (
            .O(N__4820),
            .I(N__4817));
    InMux I__613 (
            .O(N__4817),
            .I(N__4814));
    LocalMux I__612 (
            .O(N__4814),
            .I(\U712_CYCLE_TERM.TACK_STATE_r_sx_1 ));
    InMux I__611 (
            .O(N__4811),
            .I(N__4806));
    InMux I__610 (
            .O(N__4810),
            .I(N__4801));
    InMux I__609 (
            .O(N__4809),
            .I(N__4801));
    LocalMux I__608 (
            .O(N__4806),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__607 (
            .O(N__4801),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    InMux I__606 (
            .O(N__4796),
            .I(N__4790));
    InMux I__605 (
            .O(N__4795),
            .I(N__4790));
    LocalMux I__604 (
            .O(N__4790),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    CascadeMux I__603 (
            .O(N__4787),
            .I(\U712_CYCLE_TERM.N_286_i_0_0_cascade_ ));
    InMux I__602 (
            .O(N__4784),
            .I(N__4781));
    LocalMux I__601 (
            .O(N__4781),
            .I(N__4777));
    InMux I__600 (
            .O(N__4780),
            .I(N__4773));
    Span4Mux_v I__599 (
            .O(N__4777),
            .I(N__4770));
    InMux I__598 (
            .O(N__4776),
            .I(N__4767));
    LocalMux I__597 (
            .O(N__4773),
            .I(\U712_CHIP_RAM.N_416 ));
    Odrv4 I__596 (
            .O(N__4770),
            .I(\U712_CHIP_RAM.N_416 ));
    LocalMux I__595 (
            .O(N__4767),
            .I(\U712_CHIP_RAM.N_416 ));
    InMux I__594 (
            .O(N__4760),
            .I(N__4757));
    LocalMux I__593 (
            .O(N__4757),
            .I(N__4754));
    Odrv12 I__592 (
            .O(N__4754),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_1 ));
    CascadeMux I__591 (
            .O(N__4751),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0_a2_0_a3_0_cascade_ ));
    InMux I__590 (
            .O(N__4748),
            .I(N__4745));
    LocalMux I__589 (
            .O(N__4745),
            .I(N__4742));
    Odrv12 I__588 (
            .O(N__4742),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    CascadeMux I__587 (
            .O(N__4739),
            .I(N__4736));
    InMux I__586 (
            .O(N__4736),
            .I(N__4733));
    LocalMux I__585 (
            .O(N__4733),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0_a2_0_a3_0 ));
    InMux I__584 (
            .O(N__4730),
            .I(N__4724));
    InMux I__583 (
            .O(N__4729),
            .I(N__4724));
    LocalMux I__582 (
            .O(N__4724),
            .I(N__4715));
    InMux I__581 (
            .O(N__4723),
            .I(N__4708));
    InMux I__580 (
            .O(N__4722),
            .I(N__4708));
    InMux I__579 (
            .O(N__4721),
            .I(N__4708));
    InMux I__578 (
            .O(N__4720),
            .I(N__4701));
    InMux I__577 (
            .O(N__4719),
            .I(N__4701));
    InMux I__576 (
            .O(N__4718),
            .I(N__4701));
    Odrv4 I__575 (
            .O(N__4715),
            .I(\U712_CHIP_RAM.N_45 ));
    LocalMux I__574 (
            .O(N__4708),
            .I(\U712_CHIP_RAM.N_45 ));
    LocalMux I__573 (
            .O(N__4701),
            .I(\U712_CHIP_RAM.N_45 ));
    CascadeMux I__572 (
            .O(N__4694),
            .I(\U712_CHIP_RAM.N_61_cascade_ ));
    CascadeMux I__571 (
            .O(N__4691),
            .I(N__4688));
    InMux I__570 (
            .O(N__4688),
            .I(N__4683));
    InMux I__569 (
            .O(N__4687),
            .I(N__4680));
    InMux I__568 (
            .O(N__4686),
            .I(N__4677));
    LocalMux I__567 (
            .O(N__4683),
            .I(N__4674));
    LocalMux I__566 (
            .O(N__4680),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__565 (
            .O(N__4677),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    Odrv12 I__564 (
            .O(N__4674),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    InMux I__563 (
            .O(N__4667),
            .I(N__4664));
    LocalMux I__562 (
            .O(N__4664),
            .I(\U712_CHIP_RAM.N_263 ));
    InMux I__561 (
            .O(N__4661),
            .I(N__4657));
    CascadeMux I__560 (
            .O(N__4660),
            .I(N__4653));
    LocalMux I__559 (
            .O(N__4657),
            .I(N__4650));
    InMux I__558 (
            .O(N__4656),
            .I(N__4647));
    InMux I__557 (
            .O(N__4653),
            .I(N__4644));
    Odrv4 I__556 (
            .O(N__4650),
            .I(\U712_CHIP_RAM.N_271 ));
    LocalMux I__555 (
            .O(N__4647),
            .I(\U712_CHIP_RAM.N_271 ));
    LocalMux I__554 (
            .O(N__4644),
            .I(\U712_CHIP_RAM.N_271 ));
    CascadeMux I__553 (
            .O(N__4637),
            .I(\U712_CHIP_RAM.N_341_cascade_ ));
    InMux I__552 (
            .O(N__4634),
            .I(N__4631));
    LocalMux I__551 (
            .O(N__4631),
            .I(\U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0 ));
    InMux I__550 (
            .O(N__4628),
            .I(N__4625));
    LocalMux I__549 (
            .O(N__4625),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_i_0_2 ));
    InMux I__548 (
            .O(N__4622),
            .I(N__4619));
    LocalMux I__547 (
            .O(N__4619),
            .I(N__4616));
    Span4Mux_v I__546 (
            .O(N__4616),
            .I(N__4613));
    Span4Mux_v I__545 (
            .O(N__4613),
            .I(N__4610));
    Sp12to4 I__544 (
            .O(N__4610),
            .I(N__4607));
    Span12Mux_h I__543 (
            .O(N__4607),
            .I(N__4604));
    Odrv12 I__542 (
            .O(N__4604),
            .I(A_c_20));
    CascadeMux I__541 (
            .O(N__4601),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_ ));
    InMux I__540 (
            .O(N__4598),
            .I(N__4595));
    LocalMux I__539 (
            .O(N__4595),
            .I(\U712_CHIP_RAM.N_362 ));
    InMux I__538 (
            .O(N__4592),
            .I(N__4588));
    InMux I__537 (
            .O(N__4591),
            .I(N__4585));
    LocalMux I__536 (
            .O(N__4588),
            .I(\U712_CHIP_RAM.N_470 ));
    LocalMux I__535 (
            .O(N__4585),
            .I(\U712_CHIP_RAM.N_470 ));
    CascadeMux I__534 (
            .O(N__4580),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_1_0_cascade_ ));
    InMux I__533 (
            .O(N__4577),
            .I(N__4574));
    LocalMux I__532 (
            .O(N__4574),
            .I(\U712_CHIP_RAM.N_344 ));
    InMux I__531 (
            .O(N__4571),
            .I(N__4568));
    LocalMux I__530 (
            .O(N__4568),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_i_i_a3_0_0 ));
    CascadeMux I__529 (
            .O(N__4565),
            .I(\U712_CHIP_RAM.N_344_cascade_ ));
    CascadeMux I__528 (
            .O(N__4562),
            .I(N__4558));
    InMux I__527 (
            .O(N__4561),
            .I(N__4554));
    InMux I__526 (
            .O(N__4558),
            .I(N__4551));
    InMux I__525 (
            .O(N__4557),
            .I(N__4548));
    LocalMux I__524 (
            .O(N__4554),
            .I(\U712_CHIP_RAM.N_267 ));
    LocalMux I__523 (
            .O(N__4551),
            .I(\U712_CHIP_RAM.N_267 ));
    LocalMux I__522 (
            .O(N__4548),
            .I(\U712_CHIP_RAM.N_267 ));
    InMux I__521 (
            .O(N__4541),
            .I(N__4538));
    LocalMux I__520 (
            .O(N__4538),
            .I(N__4535));
    Odrv4 I__519 (
            .O(N__4535),
            .I(\U712_CHIP_RAM.N_333 ));
    CascadeMux I__518 (
            .O(N__4532),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_0_cascade_ ));
    InMux I__517 (
            .O(N__4529),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    InMux I__516 (
            .O(N__4526),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    InMux I__515 (
            .O(N__4523),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__514 (
            .O(N__4520),
            .I(N__4516));
    InMux I__513 (
            .O(N__4519),
            .I(N__4513));
    LocalMux I__512 (
            .O(N__4516),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__511 (
            .O(N__4513),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    InMux I__510 (
            .O(N__4508),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__509 (
            .O(N__4505),
            .I(N__4501));
    InMux I__508 (
            .O(N__4504),
            .I(N__4498));
    LocalMux I__507 (
            .O(N__4501),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__506 (
            .O(N__4498),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__505 (
            .O(N__4493),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    InMux I__504 (
            .O(N__4490),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    InMux I__503 (
            .O(N__4487),
            .I(N__4483));
    InMux I__502 (
            .O(N__4486),
            .I(N__4480));
    LocalMux I__501 (
            .O(N__4483),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__500 (
            .O(N__4480),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    IoInMux I__499 (
            .O(N__4475),
            .I(N__4472));
    LocalMux I__498 (
            .O(N__4472),
            .I(N__4469));
    Span4Mux_s2_v I__497 (
            .O(N__4469),
            .I(N__4466));
    Sp12to4 I__496 (
            .O(N__4466),
            .I(N__4463));
    Span12Mux_h I__495 (
            .O(N__4463),
            .I(N__4460));
    Odrv12 I__494 (
            .O(N__4460),
            .I(BANK0_c));
    InMux I__493 (
            .O(N__4457),
            .I(N__4453));
    InMux I__492 (
            .O(N__4456),
            .I(N__4450));
    LocalMux I__491 (
            .O(N__4453),
            .I(\U712_CHIP_RAM.N_404 ));
    LocalMux I__490 (
            .O(N__4450),
            .I(\U712_CHIP_RAM.N_404 ));
    CascadeMux I__489 (
            .O(N__4445),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15_cascade_ ));
    InMux I__488 (
            .O(N__4442),
            .I(N__4438));
    CascadeMux I__487 (
            .O(N__4441),
            .I(N__4435));
    LocalMux I__486 (
            .O(N__4438),
            .I(N__4432));
    InMux I__485 (
            .O(N__4435),
            .I(N__4429));
    Odrv12 I__484 (
            .O(N__4432),
            .I(LATCH_RAM));
    LocalMux I__483 (
            .O(N__4429),
            .I(LATCH_RAM));
    IoInMux I__482 (
            .O(N__4424),
            .I(N__4421));
    LocalMux I__481 (
            .O(N__4421),
            .I(N__4418));
    Span12Mux_s11_v I__480 (
            .O(N__4418),
            .I(N__4415));
    Odrv12 I__479 (
            .O(N__4415),
            .I(LATCH_CLK_0_i));
    CascadeMux I__478 (
            .O(N__4412),
            .I(\U712_CHIP_RAM.N_296_cascade_ ));
    InMux I__477 (
            .O(N__4409),
            .I(N__4406));
    LocalMux I__476 (
            .O(N__4406),
            .I(\U712_CHIP_RAM.N_296 ));
    InMux I__475 (
            .O(N__4403),
            .I(N__4400));
    LocalMux I__474 (
            .O(N__4400),
            .I(N__4397));
    Span4Mux_v I__473 (
            .O(N__4397),
            .I(N__4394));
    Odrv4 I__472 (
            .O(N__4394),
            .I(\U712_CHIP_RAM.N_63 ));
    InMux I__471 (
            .O(N__4391),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__470 (
            .O(N__4388),
            .I(N__4383));
    InMux I__469 (
            .O(N__4387),
            .I(N__4378));
    InMux I__468 (
            .O(N__4386),
            .I(N__4378));
    LocalMux I__467 (
            .O(N__4383),
            .I(N__4375));
    LocalMux I__466 (
            .O(N__4378),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    Odrv4 I__465 (
            .O(N__4375),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    InMux I__464 (
            .O(N__4370),
            .I(N__4367));
    LocalMux I__463 (
            .O(N__4367),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0 ));
    IoInMux I__462 (
            .O(N__4364),
            .I(N__4361));
    LocalMux I__461 (
            .O(N__4361),
            .I(N__4358));
    IoSpan4Mux I__460 (
            .O(N__4358),
            .I(N__4355));
    Sp12to4 I__459 (
            .O(N__4355),
            .I(N__4352));
    Span12Mux_s6_h I__458 (
            .O(N__4352),
            .I(N__4349));
    Span12Mux_v I__457 (
            .O(N__4349),
            .I(N__4345));
    InMux I__456 (
            .O(N__4348),
            .I(N__4342));
    Odrv12 I__455 (
            .O(N__4345),
            .I(TACK_OUTn));
    LocalMux I__454 (
            .O(N__4342),
            .I(TACK_OUTn));
    InMux I__453 (
            .O(N__4337),
            .I(N__4334));
    LocalMux I__452 (
            .O(N__4334),
            .I(DBR_SYNCZ0Z_0));
    InMux I__451 (
            .O(N__4331),
            .I(N__4327));
    InMux I__450 (
            .O(N__4330),
            .I(N__4324));
    LocalMux I__449 (
            .O(N__4327),
            .I(N__4321));
    LocalMux I__448 (
            .O(N__4324),
            .I(DBR_SYNCZ0Z_1));
    Odrv12 I__447 (
            .O(N__4321),
            .I(DBR_SYNCZ0Z_1));
    InMux I__446 (
            .O(N__4316),
            .I(N__4311));
    InMux I__445 (
            .O(N__4315),
            .I(N__4308));
    IoInMux I__444 (
            .O(N__4314),
            .I(N__4305));
    LocalMux I__443 (
            .O(N__4311),
            .I(N__4300));
    LocalMux I__442 (
            .O(N__4308),
            .I(N__4300));
    LocalMux I__441 (
            .O(N__4305),
            .I(N__4297));
    Span4Mux_v I__440 (
            .O(N__4300),
            .I(N__4294));
    Span12Mux_s3_h I__439 (
            .O(N__4297),
            .I(N__4291));
    Sp12to4 I__438 (
            .O(N__4294),
            .I(N__4288));
    Span12Mux_v I__437 (
            .O(N__4291),
            .I(N__4285));
    Span12Mux_h I__436 (
            .O(N__4288),
            .I(N__4282));
    Span12Mux_h I__435 (
            .O(N__4285),
            .I(N__4279));
    Span12Mux_v I__434 (
            .O(N__4282),
            .I(N__4276));
    Odrv12 I__433 (
            .O(N__4279),
            .I(CLK40_PLL));
    Odrv12 I__432 (
            .O(N__4276),
            .I(CLK40_PLL));
    CascadeMux I__431 (
            .O(N__4271),
            .I(N__4268));
    InMux I__430 (
            .O(N__4268),
            .I(N__4265));
    LocalMux I__429 (
            .O(N__4265),
            .I(N__4262));
    Odrv12 I__428 (
            .O(N__4262),
            .I(\U712_BYTE_ENABLE.N_90 ));
    CascadeMux I__427 (
            .O(N__4259),
            .I(N__4255));
    InMux I__426 (
            .O(N__4258),
            .I(N__4250));
    InMux I__425 (
            .O(N__4255),
            .I(N__4250));
    LocalMux I__424 (
            .O(N__4250),
            .I(N__4240));
    ClkMux I__423 (
            .O(N__4249),
            .I(N__4223));
    ClkMux I__422 (
            .O(N__4248),
            .I(N__4223));
    ClkMux I__421 (
            .O(N__4247),
            .I(N__4223));
    ClkMux I__420 (
            .O(N__4246),
            .I(N__4223));
    ClkMux I__419 (
            .O(N__4245),
            .I(N__4223));
    ClkMux I__418 (
            .O(N__4244),
            .I(N__4223));
    ClkMux I__417 (
            .O(N__4243),
            .I(N__4223));
    Glb2LocalMux I__416 (
            .O(N__4240),
            .I(N__4223));
    GlobalMux I__415 (
            .O(N__4223),
            .I(N__4220));
    gio2CtrlBuf I__414 (
            .O(N__4220),
            .I(CLK40_PLL_g));
    IoInMux I__413 (
            .O(N__4217),
            .I(N__4213));
    IoInMux I__412 (
            .O(N__4216),
            .I(N__4210));
    LocalMux I__411 (
            .O(N__4213),
            .I(N__4205));
    LocalMux I__410 (
            .O(N__4210),
            .I(N__4205));
    IoSpan4Mux I__409 (
            .O(N__4205),
            .I(N__4201));
    IoInMux I__408 (
            .O(N__4204),
            .I(N__4198));
    Span4Mux_s2_v I__407 (
            .O(N__4201),
            .I(N__4195));
    LocalMux I__406 (
            .O(N__4198),
            .I(N__4192));
    Sp12to4 I__405 (
            .O(N__4195),
            .I(N__4189));
    IoSpan4Mux I__404 (
            .O(N__4192),
            .I(N__4186));
    Span12Mux_v I__403 (
            .O(N__4189),
            .I(N__4183));
    Span4Mux_s3_h I__402 (
            .O(N__4186),
            .I(N__4180));
    Span12Mux_h I__401 (
            .O(N__4183),
            .I(N__4177));
    Span4Mux_h I__400 (
            .O(N__4180),
            .I(N__4174));
    Odrv12 I__399 (
            .O(N__4177),
            .I(CLK40_PLL_iso_i));
    Odrv4 I__398 (
            .O(N__4174),
            .I(CLK40_PLL_iso_i));
    InMux I__397 (
            .O(N__4169),
            .I(N__4166));
    LocalMux I__396 (
            .O(N__4166),
            .I(\U712_CHIP_RAM.N_414 ));
    CascadeMux I__395 (
            .O(N__4163),
            .I(\U712_CHIP_RAM.N_415_cascade_ ));
    CascadeMux I__394 (
            .O(N__4160),
            .I(\U712_CHIP_RAM.N_373_cascade_ ));
    CascadeMux I__393 (
            .O(N__4157),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_cascade_ ));
    CEMux I__392 (
            .O(N__4154),
            .I(N__4151));
    LocalMux I__391 (
            .O(N__4151),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_0 ));
    InMux I__390 (
            .O(N__4148),
            .I(N__4145));
    LocalMux I__389 (
            .O(N__4145),
            .I(\U712_CHIP_RAM.N_373 ));
    IoInMux I__388 (
            .O(N__4142),
            .I(N__4139));
    LocalMux I__387 (
            .O(N__4139),
            .I(N__4136));
    IoSpan4Mux I__386 (
            .O(N__4136),
            .I(N__4133));
    Span4Mux_s2_v I__385 (
            .O(N__4133),
            .I(N__4130));
    Sp12to4 I__384 (
            .O(N__4130),
            .I(N__4127));
    Odrv12 I__383 (
            .O(N__4127),
            .I(N_48_i));
    InMux I__382 (
            .O(N__4124),
            .I(N__4121));
    LocalMux I__381 (
            .O(N__4121),
            .I(N__4118));
    Span12Mux_v I__380 (
            .O(N__4118),
            .I(N__4115));
    Odrv12 I__379 (
            .O(N__4115),
            .I(RAMSPACEn_c));
    CascadeMux I__378 (
            .O(N__4112),
            .I(\U712_CHIP_RAM.N_355_cascade_ ));
    CascadeMux I__377 (
            .O(N__4109),
            .I(\U712_CHIP_RAM.N_416_cascade_ ));
    InMux I__376 (
            .O(N__4106),
            .I(N__4103));
    LocalMux I__375 (
            .O(N__4103),
            .I(\U712_CHIP_RAM.N_448 ));
    CascadeMux I__374 (
            .O(N__4100),
            .I(\U712_CHIP_RAM.N_261_cascade_ ));
    CascadeMux I__373 (
            .O(N__4097),
            .I(\U712_CHIP_RAM.N_404_cascade_ ));
    CascadeMux I__372 (
            .O(N__4094),
            .I(\U712_CHIP_RAM.N_413_cascade_ ));
    IoInMux I__371 (
            .O(N__4091),
            .I(N__4088));
    LocalMux I__370 (
            .O(N__4088),
            .I(N__4085));
    Span4Mux_s2_v I__369 (
            .O(N__4085),
            .I(N__4082));
    Span4Mux_v I__368 (
            .O(N__4082),
            .I(N__4079));
    Odrv4 I__367 (
            .O(N__4079),
            .I(CLK80_PLL_i_i));
    CascadeMux I__366 (
            .O(N__4076),
            .I(\U712_CHIP_RAM.N_448_cascade_ ));
    CascadeMux I__365 (
            .O(N__4073),
            .I(\U712_CHIP_RAM.N_459_cascade_ ));
    CascadeMux I__364 (
            .O(N__4070),
            .I(\U712_CHIP_RAM.N_308_cascade_ ));
    InMux I__363 (
            .O(N__4067),
            .I(N__4064));
    LocalMux I__362 (
            .O(N__4064),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ));
    IoInMux I__361 (
            .O(N__4061),
            .I(N__4058));
    LocalMux I__360 (
            .O(N__4058),
            .I(N__4055));
    Span4Mux_s0_v I__359 (
            .O(N__4055),
            .I(N__4052));
    Span4Mux_v I__358 (
            .O(N__4052),
            .I(N__4049));
    Sp12to4 I__357 (
            .O(N__4049),
            .I(N__4046));
    Span12Mux_h I__356 (
            .O(N__4046),
            .I(N__4043));
    Span12Mux_v I__355 (
            .O(N__4043),
            .I(N__4040));
    Odrv12 I__354 (
            .O(N__4040),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .I(N__7673));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .I(N__7675));
    INV \INVU712_REG_SM.REG_CYCLE_STARTC  (
            .O(\INVU712_REG_SM.REG_CYCLE_STARTC_net ),
            .I(N__4244));
    INV \INVU712_REG_SM.UDSnC  (
            .O(\INVU712_REG_SM.UDSnC_net ),
            .I(N__4243));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .I(N__7676));
    INV \INVU712_REG_SM.C3_SYNC_0C  (
            .O(\INVU712_REG_SM.C3_SYNC_0C_net ),
            .I(N__4245));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .I(N__7677));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .I(N__7679));
    INV \INVU712_REG_SM.STATE_COUNTER_2C  (
            .O(\INVU712_REG_SM.STATE_COUNTER_2C_net ),
            .I(N__4248));
    INV \INVU712_REG_SM.REG_CYCLEC  (
            .O(\INVU712_REG_SM.REG_CYCLEC_net ),
            .I(N__4247));
    INV \INVU712_REG_SM.STATE_COUNTER_5C  (
            .O(\INVU712_REG_SM.STATE_COUNTER_5C_net ),
            .I(N__4246));
    INV \INVU712_CHIP_RAM.DMA_A20C  (
            .O(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .I(N__7678));
    INV \INVU712_REG_SM.DBR_SYNC_1C  (
            .O(\INVU712_REG_SM.DBR_SYNC_1C_net ),
            .I(N__4249));
    defparam IN_MUX_bfv_12_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_10_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_8_0_));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__7516),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    ICE_GB CLK40_PLL_derived_clock_RNIIOT (
            .USERSIGNALTOGLOBALBUFFER(N__4314),
            .GLOBALBUFFEROUTPUT(CLK40_PLL_g));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__5063),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB DBRn_c_i_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__5450),
            .GLOBALBUFFEROUTPUT(DBRn_c_i_0_g));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__7151),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_3_1_4.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_3_1_4.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_3_1_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLKRAM_obuf_RNO_LC_3_1_4 (
            .in0(N__9743),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBR_SYNC_0_LC_6_12_2.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_6_12_2.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_6_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_0_LC_6_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4996),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9737),
            .ce(),
            .sr(N__10992));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_7_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_7_7_6 .LUT_INIT=16'b0111101010110101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_7_7_6  (
            .in0(N__6473),
            .in1(N__6626),
            .in2(N__6406),
            .in3(N__6192),
            .lcout(\U712_CHIP_RAM.N_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_1_LC_7_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_1_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_1_LC_7_7_7 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_1_LC_7_7_7  (
            .in0(N__6193),
            .in1(N__4780),
            .in2(N__6293),
            .in3(N__6096),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8UIP2_4_LC_7_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8UIP2_4_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8UIP2_4_LC_7_8_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI8UIP2_4_LC_7_8_0  (
            .in0(N__6471),
            .in1(N__6687),
            .in2(N__5907),
            .in3(N__5339),
            .lcout(\U712_CHIP_RAM.N_448 ),
            .ltout(\U712_CHIP_RAM.N_448_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_7_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_7_8_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_7_8_1  (
            .in0(_gnd_net_),
            .in1(N__6617),
            .in2(N__4076),
            .in3(N__6388),
            .lcout(\U712_CHIP_RAM.N_459 ),
            .ltout(\U712_CHIP_RAM.N_459_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_7_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_7_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_7_8_2 .LUT_INIT=16'b1010101010100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_7_8_2  (
            .in0(N__5207),
            .in1(_gnd_net_),
            .in2(N__4073),
            .in3(N__6200),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9726),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_7_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_7_8_3 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_7_8_3  (
            .in0(N__6267),
            .in1(N__5525),
            .in2(_gnd_net_),
            .in3(N__7934),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_308_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_7_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_7_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_7_8_4 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_7_8_4  (
            .in0(N__5208),
            .in1(N__7410),
            .in2(N__4070),
            .in3(N__4067),
            .lcout(WRITE_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9726),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIEH9V_LC_7_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIEH9V_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIEH9V_LC_7_8_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIEH9V_LC_7_8_5  (
            .in0(N__4331),
            .in1(N__4686),
            .in2(_gnd_net_),
            .in3(N__4388),
            .lcout(\U712_CHIP_RAM.N_416 ),
            .ltout(\U712_CHIP_RAM.N_416_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_3_LC_7_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_3_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_3_LC_7_8_6 .LUT_INIT=16'b0000000011111100;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_RNO_3_LC_7_8_6  (
            .in0(_gnd_net_),
            .in1(N__6266),
            .in2(N__4109),
            .in3(N__4656),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_i_i_a3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISAAQ_4_LC_7_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISAAQ_4_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISAAQ_4_LC_7_9_0 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNISAAQ_4_LC_7_9_0  (
            .in0(_gnd_net_),
            .in1(N__5891),
            .in2(_gnd_net_),
            .in3(N__6160),
            .lcout(\U712_CHIP_RAM.N_271 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJIDU3_0_LC_7_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJIDU3_0_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJIDU3_0_LC_7_9_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIJIDU3_0_LC_7_9_1  (
            .in0(N__6360),
            .in1(N__4106),
            .in2(N__4562),
            .in3(N__10635),
            .lcout(\U712_CHIP_RAM.N_113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI94JE1_LC_7_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI94JE1_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI94JE1_LC_7_9_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNI94JE1_LC_7_9_2  (
            .in0(N__7000),
            .in1(N__6571),
            .in2(N__6719),
            .in3(N__5893),
            .lcout(\U712_CHIP_RAM.N_414 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_7_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_7_9_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_7_9_3  (
            .in0(N__4486),
            .in1(N__4504),
            .in2(_gnd_net_),
            .in3(N__4519),
            .lcout(\U712_CHIP_RAM.N_261 ),
            .ltout(\U712_CHIP_RAM.N_261_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI41LA2_1_LC_7_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI41LA2_1_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI41LA2_1_LC_7_9_4 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI41LA2_1_LC_7_9_4  (
            .in0(_gnd_net_),
            .in1(N__6445),
            .in2(N__4100),
            .in3(N__6358),
            .lcout(\U712_CHIP_RAM.N_404 ),
            .ltout(\U712_CHIP_RAM.N_404_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0CV43_4_LC_7_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0CV43_4_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0CV43_4_LC_7_9_5 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI0CV43_4_LC_7_9_5  (
            .in0(N__5892),
            .in1(_gnd_net_),
            .in2(N__4097),
            .in3(N__6161),
            .lcout(\U712_CHIP_RAM.N_449 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_1_LC_7_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_1_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_1_LC_7_9_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_1_LC_7_9_6  (
            .in0(N__6688),
            .in1(N__5340),
            .in2(N__4660),
            .in3(N__6446),
            .lcout(\U712_CHIP_RAM.N_413 ),
            .ltout(\U712_CHIP_RAM.N_413_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIPJCN3_LC_7_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIPJCN3_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIPJCN3_LC_7_9_7 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIPJCN3_LC_7_9_7  (
            .in0(N__6359),
            .in1(_gnd_net_),
            .in2(N__4094),
            .in3(N__7406),
            .lcout(\U712_CHIP_RAM.N_470 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIC9HD1_LC_7_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIC9HD1_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIC9HD1_LC_7_10_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIC9HD1_LC_7_10_0  (
            .in0(N__6720),
            .in1(N__6294),
            .in2(_gnd_net_),
            .in3(N__6581),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_415_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKV5I5_LC_7_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKV5I5_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKV5I5_LC_7_10_1 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKV5I5_LC_7_10_1  (
            .in0(N__6202),
            .in1(N__4169),
            .in2(N__4163),
            .in3(N__4457),
            .lcout(\U712_CHIP_RAM.N_373 ),
            .ltout(\U712_CHIP_RAM.N_373_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNICBGO9_2_LC_7_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNICBGO9_2_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNICBGO9_2_LC_7_10_2 .LUT_INIT=16'b1111001111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNICBGO9_2_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(N__6582),
            .in2(N__4160),
            .in3(N__4591),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_7_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_7_10_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_7_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4157),
            .in3(N__11029),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_7_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_7_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_7_10_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_LC_7_10_4  (
            .in0(N__6093),
            .in1(N__6203),
            .in2(_gnd_net_),
            .in3(N__6295),
            .lcout(DMA_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9730),
            .ce(N__4154),
            .sr(N__11000));
    defparam \U712_CHIP_RAM.LATCH_RAM_RNO_1_LC_7_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_RAM_RNO_1_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_RAM_RNO_1_LC_7_10_6 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \U712_CHIP_RAM.LATCH_RAM_RNO_1_LC_7_10_6  (
            .in0(N__4148),
            .in1(N__4561),
            .in2(N__6404),
            .in3(N__5607),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_48_i_LC_7_11_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_48_i_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_48_i_LC_7_11_0 .LUT_INIT=16'b0100110001011111;
    LogicCell40 \U712_BYTE_ENABLE.N_48_i_LC_7_11_0  (
            .in0(N__10646),
            .in1(N__10784),
            .in2(N__4271),
            .in3(N__6943),
            .lcout(N_48_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_7_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_7_11_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_7_11_3  (
            .in0(N__4387),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10645),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_355_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_7_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_7_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_7_11_4 .LUT_INIT=16'b1100000011000100;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_7_11_4  (
            .in0(N__4124),
            .in1(N__5169),
            .in2(N__4112),
            .in3(N__8011),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9732),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_7_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_7_11_6 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(N__4330),
            .in2(_gnd_net_),
            .in3(N__4386),
            .lcout(\U712_CHIP_RAM.N_263 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_RAM_LC_7_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_RAM_LC_7_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.LATCH_RAM_LC_7_11_7 .LUT_INIT=16'b0010001010100000;
    LogicCell40 \U712_CHIP_RAM.LATCH_RAM_LC_7_11_7  (
            .in0(N__5170),
            .in1(N__4403),
            .in2(N__4441),
            .in3(N__4370),
            .lcout(LATCH_RAM),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9732),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_7_12_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_7_12_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_7_12_0 .LUT_INIT=16'b1111111110001010;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_7_12_0  (
            .in0(N__4348),
            .in1(N__4315),
            .in2(N__5840),
            .in3(N__4811),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9735),
            .ce(),
            .sr(N__10987));
    defparam DBR_SYNC_1_LC_7_12_3.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_7_12_3.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_7_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_7_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4337),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9735),
            .ce(),
            .sr(N__10987));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_7_13_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_7_13_0 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_7_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__5205),
            .in2(_gnd_net_),
            .in3(N__4832),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9738),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_7_13_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_7_13_1 .LUT_INIT=16'b0101011101110111;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_7_13_1  (
            .in0(N__5206),
            .in1(N__5789),
            .in2(N__4259),
            .in3(N__5833),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_r_sx_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_7_13_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_7_13_3 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_7_13_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_7_13_3  (
            .in0(N__5204),
            .in1(N__4316),
            .in2(_gnd_net_),
            .in3(N__5834),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9738),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LLBE_i_o4_0_o3_LC_7_13_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LLBE_i_o4_0_o3_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LLBE_i_o4_0_o3_LC_7_13_6 .LUT_INIT=16'b1110110111100101;
    LogicCell40 \U712_BYTE_ENABLE.LLBE_i_o4_0_o3_LC_7_13_6  (
            .in0(N__10244),
            .in1(N__10319),
            .in2(N__10424),
            .in3(N__10141),
            .lcout(\U712_BYTE_ENABLE.N_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLK40_PLL_derived_clock_RNIIOT_0_LC_7_13_7.C_ON=1'b0;
    defparam CLK40_PLL_derived_clock_RNIIOT_0_LC_7_13_7.SEQ_MODE=4'b0000;
    defparam CLK40_PLL_derived_clock_RNIIOT_0_LC_7_13_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLK40_PLL_derived_clock_RNIIOT_0_LC_7_13_7 (
            .in0(N__4258),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK40_PLL_iso_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.LATCH_CLK_0_i_LC_7_15_0 .C_ON=1'b0;
    defparam \U712_BUFFERS.LATCH_CLK_0_i_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.LATCH_CLK_0_i_LC_7_15_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_BUFFERS.LATCH_CLK_0_i_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(N__5762),
            .in2(_gnd_net_),
            .in3(N__4442),
            .lcout(LATCH_CLK_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_8_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_8_7_0 .LUT_INIT=16'b1111000010110000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_8_7_0  (
            .in0(N__7697),
            .in1(N__7547),
            .in2(N__5215),
            .in3(N__6956),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9723),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_7_1 .LUT_INIT=16'b1100111010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_7_1  (
            .in0(N__6269),
            .in1(N__4844),
            .in2(N__7013),
            .in3(N__5200),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9723),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_7_2 .LUT_INIT=16'b0111001101100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_7_2  (
            .in0(N__6195),
            .in1(N__6475),
            .in2(N__6629),
            .in3(N__6739),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_63_i_a2_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIRILU_LC_8_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIRILU_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIRILU_LC_8_7_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIRILU_LC_8_7_4  (
            .in0(_gnd_net_),
            .in1(N__4687),
            .in2(_gnd_net_),
            .in3(N__6268),
            .lcout(\U712_CHIP_RAM.N_296 ),
            .ltout(\U712_CHIP_RAM.N_296_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_8_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_8_7_5 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_8_7_5  (
            .in0(N__6474),
            .in1(N__5904),
            .in2(N__4412),
            .in3(N__6196),
            .lcout(\U712_CHIP_RAM.N_312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_7_7 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_7_7  (
            .in0(N__4409),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6194),
            .lcout(\U712_CHIP_RAM.N_333 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_RAM_RNO_0_LC_8_8_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.LATCH_RAM_RNO_0_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_RAM_RNO_0_LC_8_8_0 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_CHIP_RAM.LATCH_RAM_RNO_0_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__6389),
            .in2(_gnd_net_),
            .in3(N__7001),
            .lcout(\U712_CHIP_RAM.N_63 ),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_1_LC_8_8_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_1_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_1_LC_8_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_1_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(N__6472),
            .in2(_gnd_net_),
            .in3(N__4391),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_8_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__6613),
            .in2(_gnd_net_),
            .in3(N__4529),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_8_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_8_3  (
            .in0(N__4718),
            .in1(N__6736),
            .in2(_gnd_net_),
            .in3(N__4526),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__9725),
            .ce(N__5680),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_8_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_8_4  (
            .in0(N__4729),
            .in1(N__5906),
            .in2(_gnd_net_),
            .in3(N__4523),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__9725),
            .ce(N__5680),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_8_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_8_5  (
            .in0(N__4719),
            .in1(N__4520),
            .in2(_gnd_net_),
            .in3(N__4508),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__9725),
            .ce(N__5680),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_8_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_8_6  (
            .in0(N__4730),
            .in1(N__4505),
            .in2(_gnd_net_),
            .in3(N__4493),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__9725),
            .ce(N__5680),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_8_7  (
            .in0(N__4720),
            .in1(N__4487),
            .in2(_gnd_net_),
            .in3(N__4490),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9725),
            .ce(N__5680),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_esr_LC_8_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_LC_8_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.BANK0_esr_LC_8_9_0 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_LC_8_9_0  (
            .in0(N__4598),
            .in1(N__6297),
            .in2(N__6095),
            .in3(N__5662),
            .lcout(BANK0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9727),
            .ce(N__5645),
            .sr(N__11001));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_3_LC_8_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_3_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_3_LC_8_9_1 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_3_LC_8_9_1  (
            .in0(N__6692),
            .in1(_gnd_net_),
            .in2(N__6606),
            .in3(N__4456),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER15 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIURFN4_LC_8_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIURFN4_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIURFN4_LC_8_9_2 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIURFN4_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__4776),
            .in2(N__4445),
            .in3(N__6296),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa ),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_8_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_8_9_3 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_8_9_3  (
            .in0(N__4622),
            .in1(_gnd_net_),
            .in2(N__4601),
            .in3(N__9971),
            .lcout(\U712_CHIP_RAM.N_362 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIP0AC7_3_LC_8_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIP0AC7_3_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIP0AC7_3_LC_8_9_4 .LUT_INIT=16'b0000101000000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIP0AC7_3_LC_8_9_4  (
            .in0(N__5214),
            .in1(N__5236),
            .in2(N__6094),
            .in3(N__6694),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIUMPVI_3_LC_8_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIUMPVI_3_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIUMPVI_3_LC_8_9_5 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIUMPVI_3_LC_8_9_5  (
            .in0(N__5254),
            .in1(N__4592),
            .in2(N__4580),
            .in3(N__4577),
            .lcout(\U712_CHIP_RAM.N_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8MK44_LC_8_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8MK44_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8MK44_LC_8_9_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8MK44_LC_8_9_6  (
            .in0(N__6987),
            .in1(N__6693),
            .in2(N__6627),
            .in3(N__5235),
            .lcout(\U712_CHIP_RAM.N_344 ),
            .ltout(\U712_CHIP_RAM.N_344_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_2_LC_8_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_2_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_2_LC_8_9_7 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_RNO_2_LC_8_9_7  (
            .in0(N__4571),
            .in1(N__5545),
            .in2(N__4565),
            .in3(N__6077),
            .lcout(\U712_CHIP_RAM.N_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_LC_8_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_LC_8_10_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_LC_8_10_0  (
            .in0(N__4557),
            .in1(N__6370),
            .in2(_gnd_net_),
            .in3(N__5600),
            .lcout(\U712_CHIP_RAM.N_342 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIO6DI_LC_8_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIO6DI_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIO6DI_LC_8_10_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIO6DI_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(N__7416),
            .in2(_gnd_net_),
            .in3(N__6567),
            .lcout(\U712_CHIP_RAM.N_267 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_8_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_8_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(N__4891),
            .in2(_gnd_net_),
            .in3(N__6371),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_s_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_10_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_10_3  (
            .in0(N__5087),
            .in1(N__4541),
            .in2(N__4532),
            .in3(N__4721),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9729),
            .ce(N__5684),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIMQBQ1_LC_8_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIMQBQ1_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIMQBQ1_LC_8_10_4 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIMQBQ1_LC_8_10_4  (
            .in0(N__4784),
            .in1(N__6298),
            .in2(_gnd_net_),
            .in3(N__6207),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0_a2_0_a3_0 ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0_a2_0_a3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_10_5 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_10_5  (
            .in0(N__5085),
            .in1(N__4760),
            .in2(N__4751),
            .in3(N__4722),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9729),
            .ce(N__5684),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_10_7 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_10_7  (
            .in0(N__5086),
            .in1(N__4748),
            .in2(N__4739),
            .in3(N__4723),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9729),
            .ce(N__5684),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_11_0 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_11_0  (
            .in0(N__7418),
            .in1(N__10573),
            .in2(N__6740),
            .in3(N__5638),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_61_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_11_1 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_8_11_1  (
            .in0(N__5041),
            .in1(N__5129),
            .in2(N__4694),
            .in3(N__4634),
            .lcout(CPU_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9731),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIMQBQ1_LC_8_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIMQBQ1_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIMQBQ1_LC_8_11_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIMQBQ1_LC_8_11_2  (
            .in0(N__6276),
            .in1(N__6201),
            .in2(N__4691),
            .in3(N__4667),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_11_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_11_3  (
            .in0(N__6730),
            .in1(N__7417),
            .in2(_gnd_net_),
            .in3(N__6373),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_341_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_11_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_11_4  (
            .in0(N__4628),
            .in1(N__4661),
            .in2(N__4637),
            .in3(N__5350),
            .lcout(\U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_11_6 .LUT_INIT=16'b1100111001111111;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_11_6  (
            .in0(N__6372),
            .in1(N__6599),
            .in2(N__6489),
            .in3(N__6729),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_i_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBRn_ibuf_RNIBAB_LC_8_12_1.C_ON=1'b0;
    defparam DBRn_ibuf_RNIBAB_LC_8_12_1.SEQ_MODE=4'b0000;
    defparam DBRn_ibuf_RNIBAB_LC_8_12_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 DBRn_ibuf_RNIBAB_LC_8_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4997),
            .lcout(DBRn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_8_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_8_12_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_8_12_6  (
            .in0(N__4796),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5183),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9733),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_8_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_8_12_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_8_12_7  (
            .in0(_gnd_net_),
            .in1(N__4850),
            .in2(_gnd_net_),
            .in3(N__4795),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_START_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_13_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_13_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_13_0  (
            .in0(N__4831),
            .in1(N__5036),
            .in2(N__5839),
            .in3(N__4809),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_8_13_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_8_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_8_13_1 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_8_13_1  (
            .in0(N__5037),
            .in1(N__6879),
            .in2(N__4820),
            .in3(N__5832),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9736),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_8_13_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_8_13_2 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_8_13_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__5187),
            .in2(_gnd_net_),
            .in3(N__4810),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9736),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_8_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_8_13_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_8_13_3 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_8_13_3  (
            .in0(N__5185),
            .in1(N__10783),
            .in2(_gnd_net_),
            .in3(N__10868),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9736),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_8_13_4.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_8_13_4.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_8_13_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_8_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5184),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_2_LC_8_13_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_2_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_2_LC_8_13_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_2_LC_8_13_5  (
            .in0(N__5186),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5784),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_286_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_13_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_13_6 .LUT_INIT=16'b1111101011101010;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_13_6  (
            .in0(N__5800),
            .in1(N__5035),
            .in2(N__4787),
            .in3(N__6878),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_286_i_0_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_13_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_13_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5066),
            .in3(N__5053),
            .lcout(\U712_CYCLE_TERM.N_286_i_0_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_14_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_14_5 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_14_5 .LUT_INIT=16'b0111011101111111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_14_5  (
            .in0(N__5188),
            .in1(N__5788),
            .in2(N__5042),
            .in3(N__6881),
            .lcout(TACK_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9739),
            .ce(N__5006),
            .sr(N__10979));
    defparam \U712_REG_SM.DBR_SYNC_1_LC_8_15_0 .C_ON=1'b0;
    defparam \U712_REG_SM.DBR_SYNC_1_LC_8_15_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DBR_SYNC_1_LC_8_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.DBR_SYNC_1_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4955),
            .lcout(\U712_REG_SM.DBR_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.DBR_SYNC_1C_net ),
            .ce(),
            .sr(N__10977));
    defparam \U712_REG_SM.DBR_SYNC_0_LC_8_15_6 .C_ON=1'b0;
    defparam \U712_REG_SM.DBR_SYNC_0_LC_8_15_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DBR_SYNC_0_LC_8_15_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.DBR_SYNC_0_LC_8_15_6  (
            .in0(N__4992),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.DBR_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.DBR_SYNC_1C_net ),
            .ce(),
            .sr(N__10977));
    defparam TACKn_obuft_RNO_LC_8_16_1.C_ON=1'b0;
    defparam TACKn_obuft_RNO_LC_8_16_1.SEQ_MODE=4'b0000;
    defparam TACKn_obuft_RNO_LC_8_16_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 TACKn_obuft_RNO_LC_8_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4949),
            .lcout(N_977_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_VBENn_LC_9_5_0 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_LC_9_5_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_VBENn_LC_9_5_0  (
            .in0(N__10690),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5744),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_9_5_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_9_5_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_9_5_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_9_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRUMR1_4_LC_9_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRUMR1_4_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRUMR1_4_LC_9_7_0 .LUT_INIT=16'b1111010001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIRUMR1_4_LC_9_7_0  (
            .in0(N__6622),
            .in1(N__6403),
            .in2(N__6497),
            .in3(N__5905),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_o3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_9_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_9_7_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_9_7_1  (
            .in0(N__4868),
            .in1(N__5438),
            .in2(_gnd_net_),
            .in3(N__9040),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_7_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_7_2  (
            .in0(N__9037),
            .in1(N__5423),
            .in2(_gnd_net_),
            .in3(N__5405),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_7_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_7_3  (
            .in0(N__5387),
            .in1(N__5369),
            .in2(_gnd_net_),
            .in3(N__9039),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVTLS1_7_LC_9_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVTLS1_7_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVTLS1_7_LC_9_7_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVTLS1_7_LC_9_7_6  (
            .in0(_gnd_net_),
            .in1(N__5216),
            .in2(_gnd_net_),
            .in3(N__5351),
            .lcout(\U712_CHIP_RAM.N_294 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_9_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_9_7_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_9_7_7  (
            .in0(N__5318),
            .in1(N__5303),
            .in2(_gnd_net_),
            .in3(N__9038),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_8_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_8_2  (
            .in0(N__5285),
            .in1(N__5279),
            .in2(N__5273),
            .in3(N__5954),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9724),
            .ce(N__5935),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6VAGA_2_LC_9_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6VAGA_2_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6VAGA_2_LC_9_8_3 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI6VAGA_2_LC_9_8_3  (
            .in0(N__5258),
            .in1(N__6618),
            .in2(N__5618),
            .in3(N__5240),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIBVVIG_2_LC_9_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIBVVIG_2_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIBVVIG_2_LC_9_8_4 .LUT_INIT=16'b0101000111110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIBVVIG_2_LC_9_8_4  (
            .in0(N__5699),
            .in1(N__5209),
            .in2(N__5219),
            .in3(N__5077),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_3_LC_9_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_3_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_3_LC_9_8_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_3_LC_9_8_5  (
            .in0(N__5210),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6076),
            .lcout(\U712_CHIP_RAM.N_421 ),
            .ltout(\U712_CHIP_RAM.N_421_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIB13D6_4_LC_9_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIB13D6_4_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIB13D6_4_LC_9_8_6 .LUT_INIT=16'b0101111100011111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIB13D6_4_LC_9_8_6  (
            .in0(N__5698),
            .in1(N__5900),
            .in2(N__5687),
            .in3(N__6212),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_A20_LC_9_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A20_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A20_LC_9_9_0 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_A20_LC_9_9_0  (
            .in0(N__9970),
            .in1(N__5465),
            .in2(N__9413),
            .in3(N__5663),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .ce(),
            .sr(N__10993));
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_9_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_9_9_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__11028),
            .in2(_gnd_net_),
            .in3(N__5651),
            .lcout(\U712_CHIP_RAM.N_18_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_LC_9_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_9_10_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_9_10_0 .LUT_INIT=16'b1100010111001100;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_9_10_0  (
            .in0(N__5639),
            .in1(N__5566),
            .in2(N__6405),
            .in3(N__5617),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9728),
            .ce(),
            .sr(N__10988));
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_9_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_9_10_4 .LUT_INIT=16'b1010111010101100;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_LC_9_10_4  (
            .in0(N__5555),
            .in1(N__10574),
            .in2(N__5549),
            .in3(N__6224),
            .lcout(CPU_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9728),
            .ce(),
            .sr(N__10988));
    defparam \U712_CHIP_RAM.DBENn_LC_9_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_9_10_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_9_10_5 .LUT_INIT=16'b0100111011101110;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_9_10_5  (
            .in0(N__5534),
            .in1(N__7031),
            .in2(N__6101),
            .in3(N__8501),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9728),
            .ce(),
            .sr(N__10988));
    defparam \U712_CHIP_RAM.DBDIR_LC_9_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_9_10_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_9_10_7 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_9_10_7  (
            .in0(N__5524),
            .in1(N__5476),
            .in2(_gnd_net_),
            .in3(N__6041),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9728),
            .ce(),
            .sr(N__10988));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_LC_9_11_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_LC_9_11_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_LC_9_11_2  (
            .in0(N__7032),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7012),
            .lcout(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_9_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_9_11_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_9_11_4  (
            .in0(N__11027),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5461),
            .lcout(DBRn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_9_13_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_9_13_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_9_13_0 .LUT_INIT=16'b0011000010111010;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_9_13_0  (
            .in0(N__5846),
            .in1(N__5835),
            .in2(N__5804),
            .in3(N__6880),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9734),
            .ce(),
            .sr(N__10980));
    defparam \U712_REG_SM.STATE_COUNTER_5_LC_9_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_5_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_5_LC_9_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_5_LC_9_14_1  (
            .in0(N__6800),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.STATE_COUNTER_5C_net ),
            .ce(),
            .sr(N__10978));
    defparam \U712_REG_SM.STATE_COUNTER_6_LC_9_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_6_LC_9_14_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_6_LC_9_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_6_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5768),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.STATE_COUNTER_5C_net ),
            .ce(),
            .sr(N__10978));
    defparam \U712_REG_SM.LATCH_REG_LC_9_14_3 .C_ON=1'b0;
    defparam \U712_REG_SM.LATCH_REG_LC_9_14_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.LATCH_REG_LC_9_14_3 .LUT_INIT=16'b1100000011001010;
    LogicCell40 \U712_REG_SM.LATCH_REG_LC_9_14_3  (
            .in0(N__5755),
            .in1(N__7880),
            .in2(N__6785),
            .in3(N__8087),
            .lcout(LATCH_REG),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.STATE_COUNTER_5C_net ),
            .ce(),
            .sr(N__10978));
    defparam \U712_REG_SM.REG_CPU_CYCLE_LC_9_14_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CPU_CYCLE_LC_9_14_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CPU_CYCLE_LC_9_14_5 .LUT_INIT=16'b0100111000000101;
    LogicCell40 \U712_REG_SM.REG_CPU_CYCLE_LC_9_14_5  (
            .in0(N__6799),
            .in1(N__5737),
            .in2(N__7214),
            .in3(N__5723),
            .lcout(REG_CPU_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.STATE_COUNTER_5C_net ),
            .ce(),
            .sr(N__10978));
    defparam \U712_REG_SM.DBR_SYNC_RNIVIGC1_1_LC_9_15_3 .C_ON=1'b0;
    defparam \U712_REG_SM.DBR_SYNC_RNIVIGC1_1_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DBR_SYNC_RNIVIGC1_1_LC_9_15_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_REG_SM.DBR_SYNC_RNIVIGC1_1_LC_9_15_3  (
            .in0(N__8376),
            .in1(N__6753),
            .in2(N__8332),
            .in3(N__8255),
            .lcout(\U712_REG_SM.STATE_COUNTERc_0 ),
            .ltout(\U712_REG_SM.STATE_COUNTERc_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CPU_CYCLE_RNO_0_LC_9_15_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CPU_CYCLE_RNO_0_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CPU_CYCLE_RNO_0_LC_9_15_4 .LUT_INIT=16'b0100010001000111;
    LogicCell40 \U712_REG_SM.REG_CPU_CYCLE_RNO_0_LC_9_15_4  (
            .in0(N__7875),
            .in1(N__6798),
            .in2(N__5726),
            .in3(N__8076),
            .lcout(\U712_REG_SM.REG_CPU_CYCLE_e_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_9_15_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_9_15_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_9_15_7  (
            .in0(N__8377),
            .in1(N__6834),
            .in2(_gnd_net_),
            .in3(N__7874),
            .lcout(\U712_REG_SM.N_297 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_5_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_5_0  (
            .in0(N__5717),
            .in1(N__6035),
            .in2(_gnd_net_),
            .in3(N__9075),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_10_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_10_6_0 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_10_6_0  (
            .in0(N__9171),
            .in1(N__8914),
            .in2(_gnd_net_),
            .in3(N__9067),
            .lcout(\U712_CHIP_RAM.CMA_5_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_6_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_6_6  (
            .in0(N__6020),
            .in1(N__6005),
            .in2(_gnd_net_),
            .in3(N__9066),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_10_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_10_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_10_6_7 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_10_6_7  (
            .in0(N__9068),
            .in1(N__5990),
            .in2(N__10674),
            .in3(N__7067),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_7_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_7_1  (
            .in0(N__6305),
            .in1(N__6641),
            .in2(N__5974),
            .in3(N__5951),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9719),
            .ce(N__5936),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_7_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_7_3  (
            .in0(N__6503),
            .in1(N__5981),
            .in2(N__5975),
            .in3(N__5953),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9719),
            .ce(N__5936),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIP0891_1_LC_10_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIP0891_1_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIP0891_1_LC_10_7_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIP0891_1_LC_10_7_5  (
            .in0(N__6737),
            .in1(N__6490),
            .in2(_gnd_net_),
            .in3(N__6221),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_411_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIPB1M2_4_LC_10_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIPB1M2_4_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIPB1M2_4_LC_10_7_6 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIPB1M2_4_LC_10_7_6  (
            .in0(N__5912),
            .in1(N__6628),
            .in2(N__5984),
            .in3(N__6738),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_1_0 ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_7_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_7_7  (
            .in0(N__5970),
            .in1(N__6635),
            .in2(N__5957),
            .in3(N__5952),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9719),
            .ce(N__5936),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_8_0 .LUT_INIT=16'b1100111111001010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_8_0  (
            .in0(N__6619),
            .in1(N__5908),
            .in2(N__6222),
            .in3(N__6734),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_316_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_8_1 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_8_1  (
            .in0(N__6735),
            .in1(N__6211),
            .in2(N__6644),
            .in3(N__6408),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_8_3 .LUT_INIT=16'b1110110110101000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_8_3  (
            .in0(N__6214),
            .in1(N__6496),
            .in2(N__6416),
            .in3(N__6621),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_101_i_a2_0_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_8_5 .LUT_INIT=16'b0110110100101000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_8_5  (
            .in0(N__6213),
            .in1(N__6495),
            .in2(N__6415),
            .in3(N__6620),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_8_7 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_8_7  (
            .in0(N__7419),
            .in1(N__6494),
            .in2(_gnd_net_),
            .in3(N__6407),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_10_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_10_9_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_10_9_6  (
            .in0(N__6299),
            .in1(N__6223),
            .in2(_gnd_net_),
            .in3(N__6097),
            .lcout(\U712_CHIP_RAM.N_109_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_10_14_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_10_14_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_1_LC_10_14_0  (
            .in0(N__6780),
            .in1(N__6835),
            .in2(_gnd_net_),
            .in3(N__7206),
            .lcout(\U712_REG_SM.un15_0_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNTER_RNIELLV_7_LC_10_14_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_RNIELLV_7_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNTER_RNIELLV_7_LC_10_14_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_RNIELLV_7_LC_10_14_3  (
            .in0(N__7205),
            .in1(N__8319),
            .in2(_gnd_net_),
            .in3(N__8251),
            .lcout(\U712_REG_SM.LATCH_REG_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_10_15_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_10_15_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_10_15_0 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_10_15_0  (
            .in0(N__8083),
            .in1(N__10879),
            .in2(_gnd_net_),
            .in3(N__6904),
            .lcout(REG_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.REG_CYCLEC_net ),
            .ce(),
            .sr(N__10976));
    defparam \U712_REG_SM.REG_TACK_LC_10_15_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_10_15_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_10_15_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_10_15_1  (
            .in0(N__6905),
            .in1(N__6896),
            .in2(N__6890),
            .in3(N__6865),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.REG_CYCLEC_net ),
            .ce(),
            .sr(N__10976));
    defparam \U712_REG_SM.C1_SYNC_1_LC_10_15_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_10_15_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.C1_SYNC_1_LC_10_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7481),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.REG_CYCLEC_net ),
            .ce(),
            .sr(N__10976));
    defparam \U712_REG_SM.STATE_COUNTER_7_LC_10_15_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_7_LC_10_15_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_7_LC_10_15_3 .LUT_INIT=16'b1111101011101010;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_7_LC_10_15_3  (
            .in0(N__6836),
            .in1(N__8326),
            .in2(N__7213),
            .in3(N__8259),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.REG_CYCLEC_net ),
            .ce(),
            .sr(N__10976));
    defparam \U712_REG_SM.C3_SYNC_1_LC_10_15_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_10_15_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.C3_SYNC_1_LC_10_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7109),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.REG_CYCLEC_net ),
            .ce(),
            .sr(N__10976));
    defparam \U712_REG_SM.REGENn_LC_10_15_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_LC_10_15_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_LC_10_15_5 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \U712_REG_SM.REGENn_LC_10_15_5  (
            .in0(N__6811),
            .in1(N__7957),
            .in2(_gnd_net_),
            .in3(N__8084),
            .lcout(REGENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.REG_CYCLEC_net ),
            .ce(),
            .sr(N__10976));
    defparam \U712_REG_SM.STATE_COUNTER_4_LC_10_15_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_4_LC_10_15_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_4_LC_10_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_4_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6784),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.REG_CYCLEC_net ),
            .ce(),
            .sr(N__10976));
    defparam \U712_REG_SM.STATE_COUNTER_3_LC_10_15_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_3_LC_10_15_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_3_LC_10_15_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_3_LC_10_15_7  (
            .in0(N__8378),
            .in1(N__8327),
            .in2(N__8261),
            .in3(N__6760),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.REG_CYCLEC_net ),
            .ce(),
            .sr(N__10976));
    defparam \U712_REG_SM.STATE_COUNTER_2_LC_10_16_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_2_LC_10_16_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_2_LC_10_16_4 .LUT_INIT=16'b1111111111010000;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_2_LC_10_16_4  (
            .in0(N__6764),
            .in1(N__7178),
            .in2(N__8392),
            .in3(N__7961),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.STATE_COUNTER_2C_net ),
            .ce(),
            .sr(N__10974));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_5_5 .LUT_INIT=16'b1101111111010101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_5_5  (
            .in0(N__8634),
            .in1(N__7097),
            .in2(N__10692),
            .in3(N__9569),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_5_6 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_5_6  (
            .in0(N__10686),
            .in1(N__7103),
            .in2(N__9137),
            .in3(N__8120),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_5_7 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_5_7  (
            .in0(N__8633),
            .in1(N__7096),
            .in2(N__10693),
            .in3(N__9568),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_6_2 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_6_2  (
            .in0(N__10639),
            .in1(N__7073),
            .in2(N__9136),
            .in3(N__7061),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_11_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_11_6_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_11_6_5  (
            .in0(_gnd_net_),
            .in1(N__9172),
            .in2(_gnd_net_),
            .in3(N__8915),
            .lcout(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_11_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_11_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_11_7_5  (
            .in0(N__9617),
            .in1(N__9554),
            .in2(_gnd_net_),
            .in3(N__9968),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .ce(N__9773),
            .sr(N__10994));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_11_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_11_8_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_11_8_1  (
            .in0(N__9969),
            .in1(N__9485),
            .in2(_gnd_net_),
            .in3(N__9406),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .ce(N__9770),
            .sr(N__10989));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0_LC_11_10_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0_LC_11_10_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0_LC_11_10_0  (
            .in0(N__7039),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7008),
            .lcout(\U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_10_1 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_10_1  (
            .in0(N__7768),
            .in1(N__7783),
            .in2(N__7754),
            .in3(N__7798),
            .lcout(\U712_CHIP_RAM.REFRESH5lt7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_49_i_LC_11_11_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_49_i_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_49_i_LC_11_11_3 .LUT_INIT=16'b0000110111011101;
    LogicCell40 \U712_BYTE_ENABLE.N_49_i_LC_11_11_3  (
            .in0(N__6944),
            .in1(N__10837),
            .in2(N__7250),
            .in3(N__10647),
            .lcout(N_49_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LMBE_i_o4_0_o3_LC_11_12_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LMBE_i_o4_0_o3_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LMBE_i_o4_0_o3_LC_11_12_4 .LUT_INIT=16'b1100111000111011;
    LogicCell40 \U712_BYTE_ENABLE.LMBE_i_o4_0_o3_LC_11_12_4  (
            .in0(N__10347),
            .in1(N__10251),
            .in2(N__10181),
            .in3(N__10407),
            .lcout(\U712_BYTE_ENABLE.N_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DRDDIR_0_m2_i_m2_LC_11_14_0 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_0_m2_i_m2_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_0_m2_i_m2_LC_11_14_0 .LUT_INIT=16'b0000100001111111;
    LogicCell40 \U712_BUFFERS.DRDDIR_0_m2_i_m2_LC_11_14_0  (
            .in0(N__10775),
            .in1(N__10864),
            .in2(N__7926),
            .in3(N__7426),
            .lcout(N_315),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_RNIGHT91_LC_11_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNIGHT91_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNIGHT91_LC_11_14_1 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNIGHT91_LC_11_14_1  (
            .in0(N__8480),
            .in1(N__8250),
            .in2(N__8282),
            .in3(N__7204),
            .lcout(\U712_REG_SM.N_278 ),
            .ltout(\U712_REG_SM.N_278_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNI5ITS1_1_LC_11_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI5ITS1_1_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI5ITS1_1_LC_11_14_2 .LUT_INIT=16'b1010101011111010;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI5ITS1_1_LC_11_14_2  (
            .in0(N__8398),
            .in1(_gnd_net_),
            .in2(N__7217),
            .in3(N__8318),
            .lcout(\U712_REG_SM.C1_SYNC_RNI5ITS1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.UDSn_RNO_1_LC_11_14_4 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_RNO_1_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDSn_RNO_1_LC_11_14_4 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \U712_REG_SM.UDSn_RNO_1_LC_11_14_4  (
            .in0(N__7174),
            .in1(N__7162),
            .in2(N__8399),
            .in3(N__8421),
            .lcout(\U712_REG_SM.UDSn_7_iv_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNTER_RNI5J3V_7_LC_11_14_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_RNI5J3V_7_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNTER_RNI5J3V_7_LC_11_14_5 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_RNI5J3V_7_LC_11_14_5  (
            .in0(N__8479),
            .in1(N__7919),
            .in2(_gnd_net_),
            .in3(N__7203),
            .lcout(\U712_REG_SM.N_309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_11_14_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_11_14_6 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_11_14_6  (
            .in0(N__8249),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8317),
            .lcout(\U712_REG_SM.N_272 ),
            .ltout(\U712_REG_SM.N_272_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDSn_RNO_1_LC_11_14_7 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_RNO_1_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDSn_RNO_1_LC_11_14_7 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \U712_REG_SM.LDSn_RNO_1_LC_11_14_7  (
            .in0(N__7163),
            .in1(N__8394),
            .in2(N__7154),
            .in3(N__7335),
            .lcout(\U712_REG_SM.LDSn_7_iv_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_0_LC_11_15_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_11_15_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.C3_SYNC_0_LC_11_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7132),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.C3_SYNC_0C_net ),
            .ce(),
            .sr(N__10975));
    defparam \U712_REG_SM.C1_SYNC_0_LC_11_15_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_11_15_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.C1_SYNC_0_LC_11_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7517),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.C3_SYNC_0C_net ),
            .ce(),
            .sr(N__10975));
    defparam \U712_REG_SM.LDSn_LC_11_15_3 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_LC_11_15_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.LDSn_LC_11_15_3 .LUT_INIT=16'b1111101011001100;
    LogicCell40 \U712_REG_SM.LDSn_LC_11_15_3  (
            .in0(N__7310),
            .in1(N__7336),
            .in2(N__7475),
            .in3(N__7634),
            .lcout(LDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.C3_SYNC_0C_net ),
            .ce(),
            .sr(N__10975));
    defparam \U712_REG_SM.ASn_LC_11_15_4 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_LC_11_15_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_LC_11_15_4 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \U712_REG_SM.ASn_LC_11_15_4  (
            .in0(N__7463),
            .in1(N__7441),
            .in2(N__8336),
            .in3(N__8085),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.C3_SYNC_0C_net ),
            .ce(),
            .sr(N__10975));
    defparam \U712_BUFFERS.DMA_LATCH_EN_i_LC_11_16_2 .C_ON=1'b0;
    defparam \U712_BUFFERS.DMA_LATCH_EN_i_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DMA_LATCH_EN_i_LC_11_16_2 .LUT_INIT=16'b1111111100000111;
    LogicCell40 \U712_BUFFERS.DMA_LATCH_EN_i_LC_11_16_2  (
            .in0(N__10857),
            .in1(N__10763),
            .in2(N__7430),
            .in3(N__7873),
            .lcout(N_259),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDSn_RNO_2_LC_11_16_3 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_RNO_2_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDSn_RNO_2_LC_11_16_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_REG_SM.LDSn_RNO_2_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(N__7334),
            .in2(_gnd_net_),
            .in3(N__8375),
            .lcout(),
            .ltout(\U712_REG_SM.N_467_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDSn_RNO_0_LC_11_16_4 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_11_16_4 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \U712_REG_SM.LDSn_RNO_0_LC_11_16_4  (
            .in0(N__10130),
            .in1(N__10259),
            .in2(N__7313),
            .in3(N__8491),
            .lcout(\U712_REG_SM.N_371 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_5_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_5_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_12_5_0  (
            .in0(N__7616),
            .in1(N__7622),
            .in2(_gnd_net_),
            .in3(N__7304),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9714),
            .ce(N__9647),
            .sr(N__10999));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_12_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_12_5_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_12_5_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_12_5_7  (
            .in0(N__7289),
            .in1(N__7283),
            .in2(_gnd_net_),
            .in3(N__7256),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9714),
            .ce(N__9647),
            .sr(N__10999));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_6_2 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_6_2  (
            .in0(N__8750),
            .in1(N__9118),
            .in2(_gnd_net_),
            .in3(N__7586),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_6_4 .LUT_INIT=16'b0000001011110000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_6_4  (
            .in0(N__8584),
            .in1(N__10641),
            .in2(N__8773),
            .in3(N__9117),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_6_6 .LUT_INIT=16'b0000111011111111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_6_6  (
            .in0(N__8585),
            .in1(N__10640),
            .in2(N__8774),
            .in3(N__9116),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_7_5 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_7_5  (
            .in0(N__7610),
            .in1(N__10655),
            .in2(N__9122),
            .in3(N__7535),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_12_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_12_7_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_12_7_6  (
            .in0(N__8919),
            .in1(N__9173),
            .in2(N__8972),
            .in3(N__9090),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_7_7 .LUT_INIT=16'b1011100010111000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_7_7  (
            .in0(N__7601),
            .in1(N__10654),
            .in2(N__8102),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_329 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_8_4  (
            .in0(N__7580),
            .in1(N__7562),
            .in2(_gnd_net_),
            .in3(N__9076),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_12_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_12_8_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_12_8_7  (
            .in0(_gnd_net_),
            .in1(N__7718),
            .in2(_gnd_net_),
            .in3(N__7736),
            .lcout(\U712_CHIP_RAM.REFRESH5lto7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_9_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_9_0  (
            .in0(N__9537),
            .in1(N__10076),
            .in2(_gnd_net_),
            .in3(N__9961),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__9771),
            .sr(N__10981));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_12_10_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_12_10_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_12_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(N__7526),
            .in2(_gnd_net_),
            .in3(N__7520),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_12_10_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__7674),
            .ce(),
            .sr(N__7652));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_12_10_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_12_10_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_12_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(N__7799),
            .in2(_gnd_net_),
            .in3(N__7787),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__7674),
            .ce(),
            .sr(N__7652));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_12_10_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_12_10_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_12_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(N__7784),
            .in2(_gnd_net_),
            .in3(N__7772),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__7674),
            .ce(),
            .sr(N__7652));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_12_10_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_12_10_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_12_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__7769),
            .in2(_gnd_net_),
            .in3(N__7757),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__7674),
            .ce(),
            .sr(N__7652));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_12_10_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_12_10_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_12_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(N__7753),
            .in2(_gnd_net_),
            .in3(N__7739),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__7674),
            .ce(),
            .sr(N__7652));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_12_10_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_12_10_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_12_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(N__7735),
            .in2(_gnd_net_),
            .in3(N__7721),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__7674),
            .ce(),
            .sr(N__7652));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_12_10_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_12_10_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_12_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_12_10_6  (
            .in0(_gnd_net_),
            .in1(N__7717),
            .in2(_gnd_net_),
            .in3(N__7703),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__7674),
            .ce(),
            .sr(N__7652));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_12_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_12_10_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_12_10_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(N__7693),
            .in2(_gnd_net_),
            .in3(N__7700),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7674),
            .ce(),
            .sr(N__7652));
    defparam \U712_REG_SM.UDSn_LC_12_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_LC_12_14_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.UDSn_LC_12_14_1 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \U712_REG_SM.UDSn_LC_12_14_1  (
            .in0(N__7640),
            .in1(N__8447),
            .in2(N__8428),
            .in3(N__7633),
            .lcout(UDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.UDSnC_net ),
            .ce(),
            .sr(N__10973));
    defparam \U712_REG_SM.STATE_COUNTER_0_LC_12_14_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_0_LC_12_14_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNTER_0_LC_12_14_6 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_0_LC_12_14_6  (
            .in0(N__8086),
            .in1(N__8216),
            .in2(_gnd_net_),
            .in3(N__8490),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.UDSnC_net ),
            .ce(),
            .sr(N__10973));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_12_15_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_12_15_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_12_15_0 .LUT_INIT=16'b0011011100000101;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_12_15_0  (
            .in0(N__8044),
            .in1(N__7970),
            .in2(N__8012),
            .in3(N__8281),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.REG_CYCLE_STARTC_net ),
            .ce(),
            .sr(N__10972));
    defparam \U712_REG_SM.CYCLE_RUN_LC_12_15_2 .C_ON=1'b0;
    defparam \U712_REG_SM.CYCLE_RUN_LC_12_15_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.CYCLE_RUN_LC_12_15_2 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \U712_REG_SM.CYCLE_RUN_LC_12_15_2  (
            .in0(N__8214),
            .in1(N__7969),
            .in2(N__8492),
            .in3(N__7950),
            .lcout(\U712_REG_SM.CYCLE_RUNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.REG_CYCLE_STARTC_net ),
            .ce(),
            .sr(N__10972));
    defparam \U712_REG_SM.STATE_COUNTER_1_LC_12_15_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_1_LC_12_15_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_1_LC_12_15_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_1_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(N__8213),
            .in2(_gnd_net_),
            .in3(N__8488),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.REG_CYCLE_STARTC_net ),
            .ce(),
            .sr(N__10972));
    defparam \U712_REG_SM.REG_WRITE_CYCLE_LC_12_15_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_WRITE_CYCLE_LC_12_15_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REG_WRITE_CYCLE_LC_12_15_7 .LUT_INIT=16'b1111000001110100;
    LogicCell40 \U712_REG_SM.REG_WRITE_CYCLE_LC_12_15_7  (
            .in0(N__7927),
            .in1(N__8489),
            .in2(N__7879),
            .in3(N__8215),
            .lcout(REG_WRITE_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.REG_CYCLE_STARTC_net ),
            .ce(),
            .sr(N__10972));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_13_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_13_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_13_5_0 .LUT_INIT=16'b0000011000000111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_13_5_0  (
            .in0(N__9183),
            .in1(N__9123),
            .in2(N__8980),
            .in3(N__8928),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_CMA28_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_13_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_13_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_13_5_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_13_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7844),
            .in3(N__11030),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_6_0 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_13_6_0  (
            .in0(N__8775),
            .in1(N__8594),
            .in2(N__8726),
            .in3(N__8144),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9716),
            .ce(N__9655),
            .sr(N__11002));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_13_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_13_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_13_6_4 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_13_6_4  (
            .in0(N__8776),
            .in1(N__9812),
            .in2(N__8727),
            .in3(N__7823),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9716),
            .ce(N__9655),
            .sr(N__11002));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_13_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_13_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_13_6_7 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_13_6_7  (
            .in0(N__8777),
            .in1(N__8718),
            .in2(N__9437),
            .in3(N__8180),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9716),
            .ce(N__9655),
            .sr(N__11002));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9_1_LC_13_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9_1_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9_1_LC_13_7_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9_1_LC_13_7_0  (
            .in0(_gnd_net_),
            .in1(N__9124),
            .in2(_gnd_net_),
            .in3(N__10670),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_7_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_7_3  (
            .in0(N__10671),
            .in1(N__8150),
            .in2(N__9138),
            .in3(N__8573),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_7_4 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_7_4  (
            .in0(N__8138),
            .in1(N__10673),
            .in2(N__9140),
            .in3(N__8093),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_13_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_13_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_13_7_7 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_13_7_7  (
            .in0(N__10672),
            .in1(N__8129),
            .in2(N__9139),
            .in3(N__8108),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_8_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_8_3  (
            .in0(N__10075),
            .in1(N__10023),
            .in2(_gnd_net_),
            .in3(N__9948),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__9775),
            .sr(N__10990));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_8_5  (
            .in0(N__9358),
            .in1(N__9611),
            .in2(_gnd_net_),
            .in3(N__9949),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__9775),
            .sr(N__10990));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_8_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_8_6  (
            .in0(N__9950),
            .in1(N__9359),
            .in2(_gnd_net_),
            .in3(N__9325),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__9775),
            .sr(N__10990));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_8_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_8_7  (
            .in0(N__9326),
            .in1(N__9484),
            .in2(_gnd_net_),
            .in3(N__9951),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__9775),
            .sr(N__10990));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_9_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_9_1  (
            .in0(N__9959),
            .in1(N__8528),
            .in2(_gnd_net_),
            .in3(N__8556),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9798),
            .ce(N__9774),
            .sr(N__10983));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_9_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_9_3  (
            .in0(N__9960),
            .in1(N__8557),
            .in2(_gnd_net_),
            .in3(N__10025),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9798),
            .ce(N__9774),
            .sr(N__10983));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_10_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_10_3  (
            .in0(N__8564),
            .in1(N__10019),
            .in2(_gnd_net_),
            .in3(N__9933),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__9772),
            .sr(N__10982));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_10_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_13_10_5  (
            .in0(N__8563),
            .in1(N__8521),
            .in2(_gnd_net_),
            .in3(N__9932),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__9772),
            .sr(N__10982));
    defparam \U712_REG_SM.UDSn_RNO_0_LC_13_14_0 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_RNO_0_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDSn_RNO_0_LC_13_14_0 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_REG_SM.UDSn_RNO_0_LC_13_14_0  (
            .in0(N__10281),
            .in1(N__8342),
            .in2(N__10187),
            .in3(N__8484),
            .lcout(\U712_REG_SM.N_369 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.UDSn_RNO_2_LC_13_14_7 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_RNO_2_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDSn_RNO_2_LC_13_14_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_REG_SM.UDSn_RNO_2_LC_13_14_7  (
            .in0(_gnd_net_),
            .in1(N__8420),
            .in2(_gnd_net_),
            .in3(N__8393),
            .lcout(\U712_REG_SM.N_465 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_RNIPBK41_LC_13_15_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNIPBK41_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNIPBK41_LC_13_15_5 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNIPBK41_LC_13_15_5  (
            .in0(N__8331),
            .in1(N__8280),
            .in2(_gnd_net_),
            .in3(N__8260),
            .lcout(\U712_REG_SM.N_288 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CASn_LC_14_2_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_14_2_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_14_2_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_14_2_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9135),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9713),
            .ce(),
            .sr(N__11014));
    defparam \U712_CHIP_RAM.WEn_LC_14_2_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_14_2_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_14_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_14_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8935),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9713),
            .ce(),
            .sr(N__11014));
    defparam \U712_CHIP_RAM.RASn_LC_14_2_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_14_2_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_14_2_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_14_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9191),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9713),
            .ce(),
            .sr(N__11014));
    defparam \U712_CHIP_RAM.CRCSn_LC_14_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_14_4_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_14_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_14_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8979),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9715),
            .ce(),
            .sr(N__11013));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_14_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_14_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_14_5_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_14_5_2  (
            .in0(N__9190),
            .in1(N__9134),
            .in2(N__8981),
            .in3(N__8936),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9717),
            .ce(N__9654),
            .sr(N__11012));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_14_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_14_5_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_14_5_7 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_14_5_7  (
            .in0(N__8645),
            .in1(N__8873),
            .in2(N__10697),
            .in3(N__9494),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9717),
            .ce(N__9654),
            .sr(N__11012));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_14_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_14_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_14_6_2 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_14_6_2  (
            .in0(N__8778),
            .in1(N__9503),
            .in2(N__8728),
            .in3(N__8831),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9718),
            .ce(N__9659),
            .sr(N__11007));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_14_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_14_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_14_6_3 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_14_6_3  (
            .in0(N__8780),
            .in1(N__8725),
            .in2(N__9281),
            .in3(N__8807),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9718),
            .ce(N__9659),
            .sr(N__11007));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_14_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_14_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_14_6_6 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_14_6_6  (
            .in0(N__8779),
            .in1(N__9623),
            .in2(N__8729),
            .in3(N__8693),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9718),
            .ce(N__9659),
            .sr(N__11007));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_6_7 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_14_6_7  (
            .in0(N__8666),
            .in1(N__8641),
            .in2(N__10691),
            .in3(N__9368),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9718),
            .ce(N__9659),
            .sr(N__11007));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_7_0  (
            .in0(N__9553),
            .in1(N__9612),
            .in2(_gnd_net_),
            .in3(N__9924),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9800),
            .ce(N__9778),
            .sr(N__11003));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_7_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_7_6  (
            .in0(N__9357),
            .in1(N__9613),
            .in2(_gnd_net_),
            .in3(N__9925),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9800),
            .ce(N__9778),
            .sr(N__11003));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_2  (
            .in0(N__10067),
            .in1(N__9546),
            .in2(_gnd_net_),
            .in3(N__9908),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9799),
            .ce(N__9777),
            .sr(N__10995));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_8_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_8_3  (
            .in0(N__9910),
            .in1(N__9477),
            .in2(_gnd_net_),
            .in3(N__9398),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9799),
            .ce(N__9777),
            .sr(N__10995));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_8_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_8_5  (
            .in0(N__9909),
            .in1(N__9324),
            .in2(_gnd_net_),
            .in3(N__9476),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9799),
            .ce(N__9777),
            .sr(N__10995));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_14_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_14_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_14_8_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_14_8_7  (
            .in0(N__9911),
            .in1(N__9425),
            .in2(_gnd_net_),
            .in3(N__9399),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9799),
            .ce(N__9777),
            .sr(N__10995));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_9_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_9_1  (
            .in0(N__9907),
            .in1(N__9351),
            .in2(_gnd_net_),
            .in3(N__9323),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9797),
            .ce(N__9776),
            .sr(N__10991));
    defparam \U712_BYTE_ENABLE.N_50_i_LC_14_11_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_50_i_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_50_i_LC_14_11_2 .LUT_INIT=16'b0101000111110011;
    LogicCell40 \U712_BYTE_ENABLE.N_50_i_LC_14_11_2  (
            .in0(N__10475),
            .in1(N__10516),
            .in2(N__10782),
            .in3(N__10678),
            .lcout(N_50_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UUBE_i_o4_0_o3_LC_14_12_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UUBE_i_o4_0_o3_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UUBE_i_o4_0_o3_LC_14_12_0 .LUT_INIT=16'b1100001111010111;
    LogicCell40 \U712_BYTE_ENABLE.UUBE_i_o4_0_o3_LC_14_12_0  (
            .in0(N__10186),
            .in1(N__10258),
            .in2(N__10423),
            .in3(N__10349),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_91_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_51_i_LC_14_12_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_51_i_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_51_i_LC_14_12_1 .LUT_INIT=16'b0101111100010011;
    LogicCell40 \U712_BYTE_ENABLE.N_51_i_LC_14_12_1  (
            .in0(N__10679),
            .in1(N__10517),
            .in2(N__10499),
            .in3(N__10836),
            .lcout(N_51_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UMBE_i_o4_0_o3_LC_14_12_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UMBE_i_o4_0_o3_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UMBE_i_o4_0_o3_LC_14_12_5 .LUT_INIT=16'b1101011111000111;
    LogicCell40 \U712_BYTE_ENABLE.UMBE_i_o4_0_o3_LC_14_12_5  (
            .in0(N__10348),
            .in1(N__10416),
            .in2(N__10272),
            .in3(N__10185),
            .lcout(\U712_BYTE_ENABLE.N_89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_90_i_LC_14_20_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_90_i_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_90_i_LC_14_20_2 .LUT_INIT=16'b0001000101001100;
    LogicCell40 \U712_BYTE_ENABLE.N_90_i_LC_14_20_2  (
            .in0(N__10336),
            .in1(N__10276),
            .in2(N__10179),
            .in3(N__10404),
            .lcout(N_90_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_92_i_LC_14_20_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_92_i_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_92_i_LC_14_20_3 .LUT_INIT=16'b0101101000010010;
    LogicCell40 \U712_BYTE_ENABLE.N_92_i_LC_14_20_3  (
            .in0(N__10406),
            .in1(N__10338),
            .in2(N__10283),
            .in3(N__10167),
            .lcout(N_92_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_91_i_LC_14_20_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_91_i_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_91_i_LC_14_20_6 .LUT_INIT=16'b0011001011001000;
    LogicCell40 \U712_BYTE_ENABLE.N_91_i_LC_14_20_6  (
            .in0(N__10337),
            .in1(N__10277),
            .in2(N__10180),
            .in3(N__10405),
            .lcout(N_91_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_89_i_LC_14_20_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_89_i_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_89_i_LC_14_20_7 .LUT_INIT=16'b0100100001011000;
    LogicCell40 \U712_BYTE_ENABLE.N_89_i_LC_14_20_7  (
            .in0(N__10403),
            .in1(N__10335),
            .in2(N__10282),
            .in3(N__10160),
            .lcout(N_89_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_16_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_16_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_16_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_16_8_4  (
            .in0(N__10068),
            .in1(N__10024),
            .in2(_gnd_net_),
            .in3(N__9955),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9796),
            .ce(N__9779),
            .sr(N__11008));
    defparam \U712_BUFFERS.un1_DRDENn_LC_24_19_4 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_DRDENn_LC_24_19_4 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_DRDENn_LC_24_19_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_BUFFERS.un1_DRDENn_LC_24_19_4  (
            .in0(N__10895),
            .in1(N__10832),
            .in2(_gnd_net_),
            .in3(N__10740),
            .lcout(DRDENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U712_TOP

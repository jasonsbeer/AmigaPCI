-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Apr 8 2025 19:54:41

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DA : out std_logic_vector(2 downto 0);
    A : in std_logic_vector(20 downto 0);
    DBRn : in std_logic;
    RAMENn : out std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    TCIn : out std_logic;
    TBIn : out std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__12194\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12067\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11967\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11770\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10380\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7972\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4084\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \U712_CYCLE_TERM_TBIn_0_i\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_13\ : std_logic;
signal \A_c_14\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.N_543_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_322_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_a2_0_0\ : std_logic;
signal \U712_CHIP_RAM.CLK_EN_6_0_a3_0_a2_1\ : std_logic;
signal \U712_CHIP_RAM.N_599_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CLK_EN_6_0\ : std_logic;
signal \U712_CHIP_RAM.N_504_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_404\ : std_logic;
signal \U712_CHIP_RAM.N_404_cascade_\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U712_CHIP_RAM.N_591\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \A_c_8\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U712_CHIP_RAM.N_578_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_545\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER18_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_552\ : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.N_554_cascade_\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \U712_CHIP_RAM.N_588\ : std_logic;
signal \U712_CHIP_RAM.N_553_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_437_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_414\ : std_logic;
signal \U712_CHIP_RAM.N_507\ : std_logic;
signal \U712_CHIP_RAM.N_507_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_506\ : std_logic;
signal \U712_CHIP_RAM.N_696\ : std_logic;
signal \U712_CHIP_RAM.N_534\ : std_logic;
signal \U712_CHIP_RAM.N_442_cascade_\ : std_logic;
signal \U712_CHIP_RAM.BANK0_RNOZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_\ : std_logic;
signal \U712_CHIP_RAM.BANK0_RNOZ0Z_1\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.BANK0_RNOZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_605_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_605\ : std_logic;
signal \U712_CHIP_RAM.N_697_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_539\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.N_697\ : std_logic;
signal \U712_CHIP_RAM.N_551\ : std_logic;
signal \U712_CHIP_RAM.N_580\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \U712_CHIP_RAM.N_505\ : std_logic;
signal \U712_CHIP_RAM.N_437\ : std_logic;
signal \U712_CHIP_RAM.N_587\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.N_70\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_REG_SM.N_513_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_589\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\ : std_logic;
signal \U712_REG_SM.N_694_cascade_\ : std_logic;
signal \U712_REG_SM.N_522_cascade_\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_START_RNOZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5\ : std_logic;
signal \U712_REG_SM.N_429_cascade_\ : std_logic;
signal \U712_REG_SM.N_511_cascade_\ : std_logic;
signal \U712_REG_SM.N_694\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_0\ : std_logic;
signal \U712_CHIP_RAM.N_700\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_0_a2_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_578\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.N_405\ : std_logic;
signal \U712_CHIP_RAM.N_699\ : std_logic;
signal \U712_CHIP_RAM.N_597_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_\ : std_logic;
signal \LATCH_CLK_c\ : std_logic;
signal \U712_CHIP_RAM.N_528\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_482_cascade_\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \U712_CHIP_RAM.N_527\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_553\ : std_logic;
signal \U712_CHIP_RAM.BANK0_0_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_597\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_537\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_703\ : std_logic;
signal \U712_CHIP_RAM.N_530_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_600\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.BANK0_0_sqmuxa_1\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0\ : std_logic;
signal \U712_CHIP_RAM.DBENn_8_0\ : std_logic;
signal \U712_REG_SM.START_RSTZ0\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_srsts_i_i_i_a2_0_0_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_2\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_0\ : std_logic;
signal \U712_REG_SM.START_RST_0_sqmuxa\ : std_logic;
signal \U712_REG_SM.un1_STATE_COUNT_4_i_i_0_0\ : std_logic;
signal \U712_REG_SM.DS_EN_RNOZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_515\ : std_logic;
signal \U712_REG_SM.N_443\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \N_549\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \bfn_11_5_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_9\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST_cascade_\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_595\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN_RNOZ0Z_0_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.N_598_cascade_\ : std_logic;
signal \U712_REG_SM.N_422\ : std_logic;
signal \U712_REG_SM.N_514\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.N_571_cascade_\ : std_logic;
signal \U712_REG_SM.N_480\ : std_logic;
signal \U712_REG_SM.REG_TACK_RNOZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_407\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \RnW_c\ : std_logic;
signal \WRITE_CYCLEm\ : std_logic;
signal \N_483\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i\ : std_logic;
signal \U712_CHIP_RAM.N_412_cascade_\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U712_CHIP_RAM.N_478\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0_cascade_\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \CLK40_PLL_i\ : std_logic;
signal \CLK40_PLL_i_i\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.N_598\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ1Z_2\ : std_logic;
signal \U712_CYCLE_TERM.N_440\ : std_logic;
signal \U712_CYCLE_TERM.un13_0\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U712_CYCLE_TERM.N_566\ : std_logic;
signal \U712_CYCLE_TERM.un13_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_93\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.N_455\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U712_CYCLE_TERM.RAM_CYCLEZ0\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \U712_CYCLE_TERM_TCIn_0_i\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U712_BYTE_ENABLE.N_563_cascade_\ : std_logic;
signal \N_56_i\ : std_logic;
signal \WEn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_i_0_8\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z20\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A20C_net\ : std_logic;
signal \N_58_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_410\ : std_logic;
signal \U712_BYTE_ENABLE.N_559\ : std_logic;
signal \N_129_i\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \RASn_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\ : std_logic;
signal \U712_CHIP_RAM.N_412\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4_cascade_\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\ : std_logic;
signal \un1_UDSn_i_0_0\ : std_logic;
signal \DS_ENm\ : std_logic;
signal \un1_LDSn_i_0_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \N_57_i\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \N_59_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_557\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \U712_BYTE_ENABLE.N_561\ : std_logic;
signal \U712_BYTE_ENABLE.N_397_i\ : std_logic;
signal \N_130_i\ : std_logic;
signal \N_127_i\ : std_logic;
signal \A_c_0\ : std_logic;
signal \A_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \N_128_i\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \DA_wire\ : std_logic_vector(2 downto 0);
signal \C3_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    TCIn <= \TCIn_wire\;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    ASn <= \ASn_wire\;
    DA <= \DA_wire\;
    \C3_wire\ <= C3;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    TBIn <= \TBIn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL_i\,
            REFERENCECLK => \N__4102\,
            RESETB => \N__7546\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12194\,
            DIN => \N__12193\,
            DOUT => \N__12192\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12194\,
            PADOUT => \N__12193\,
            PADIN => \N__12192\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9849\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12185\,
            DIN => \N__12184\,
            DOUT => \N__12183\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12185\,
            PADOUT => \N__12184\,
            PADIN => \N__12183\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12176\,
            DIN => \N__12175\,
            DOUT => \N__12174\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12176\,
            PADOUT => \N__12175\,
            PADIN => \N__12174\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9187\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12167\,
            DIN => \N__12166\,
            DOUT => \N__12165\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12167\,
            PADOUT => \N__12166\,
            PADIN => \N__12165\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7099\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12158\,
            DIN => \N__12157\,
            DOUT => \N__12156\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12158\,
            PADOUT => \N__12157\,
            PADIN => \N__12156\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12149\,
            DIN => \N__12148\,
            DOUT => \N__12147\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12149\,
            PADOUT => \N__12148\,
            PADIN => \N__12147\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12140\,
            DIN => \N__12139\,
            DOUT => \N__12138\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12140\,
            PADOUT => \N__12139\,
            PADIN => \N__12138\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12131\,
            DIN => \N__12130\,
            DOUT => \N__12129\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12131\,
            PADOUT => \N__12130\,
            PADIN => \N__12129\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12122\,
            DIN => \N__12121\,
            DOUT => \N__12120\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12122\,
            PADOUT => \N__12121\,
            PADIN => \N__12120\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12113\,
            DIN => \N__12112\,
            DOUT => \N__12111\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12113\,
            PADOUT => \N__12112\,
            PADIN => \N__12111\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12104\,
            DIN => \N__12103\,
            DOUT => \N__12102\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12104\,
            PADOUT => \N__12103\,
            PADIN => \N__12102\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8542\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12095\,
            DIN => \N__12094\,
            DOUT => \N__12093\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12095\,
            PADOUT => \N__12094\,
            PADIN => \N__12093\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9202\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12086\,
            DIN => \N__12085\,
            DOUT => \N__12084\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12086\,
            PADOUT => \N__12085\,
            PADIN => \N__12084\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12077\,
            DIN => \N__12076\,
            DOUT => \N__12075\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12077\,
            PADOUT => \N__12076\,
            PADIN => \N__12075\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5607\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12068\,
            DIN => \N__12067\,
            DOUT => \N__12066\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12068\,
            PADOUT => \N__12067\,
            PADIN => \N__12066\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12059\,
            DIN => \N__12058\,
            DOUT => \N__12057\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12059\,
            PADOUT => \N__12058\,
            PADIN => \N__12057\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12050\,
            DIN => \N__12049\,
            DOUT => \N__12048\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12050\,
            PADOUT => \N__12049\,
            PADIN => \N__12048\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4348\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12041\,
            DIN => \N__12040\,
            DOUT => \N__12039\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12041\,
            PADOUT => \N__12040\,
            PADIN => \N__12039\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12032\,
            DIN => \N__12031\,
            DOUT => \N__12030\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12032\,
            PADOUT => \N__12031\,
            PADIN => \N__12030\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12023\,
            DIN => \N__12022\,
            DOUT => \N__12021\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12023\,
            PADOUT => \N__12022\,
            PADIN => \N__12021\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7465\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12014\,
            DIN => \N__12013\,
            DOUT => \N__12012\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12014\,
            PADOUT => \N__12013\,
            PADIN => \N__12012\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12005\,
            DIN => \N__12004\,
            DOUT => \N__12003\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12005\,
            PADOUT => \N__12004\,
            PADIN => \N__12003\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8320\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11996\,
            DIN => \N__11995\,
            DOUT => \N__11994\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11996\,
            PADOUT => \N__11995\,
            PADIN => \N__11994\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11987\,
            DIN => \N__11986\,
            DOUT => \N__11985\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11987\,
            PADOUT => \N__11986\,
            PADIN => \N__11985\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10798\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11978\,
            DIN => \N__11977\,
            DOUT => \N__11976\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11978\,
            PADOUT => \N__11977\,
            PADIN => \N__11976\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11969\,
            DIN => \N__11968\,
            DOUT => \N__11967\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11969\,
            PADOUT => \N__11968\,
            PADIN => \N__11967\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11960\,
            DIN => \N__11959\,
            DOUT => \N__11958\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11960\,
            PADOUT => \N__11959\,
            PADIN => \N__11958\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11951\,
            DIN => \N__11950\,
            DOUT => \N__11949\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11951\,
            PADOUT => \N__11950\,
            PADIN => \N__11949\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11942\,
            DIN => \N__11941\,
            DOUT => \N__11940\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11942\,
            PADOUT => \N__11941\,
            PADIN => \N__11940\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11933\,
            DIN => \N__11932\,
            DOUT => \N__11931\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11933\,
            PADOUT => \N__11932\,
            PADIN => \N__11931\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6391\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11924\,
            DIN => \N__11923\,
            DOUT => \N__11922\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11924\,
            PADOUT => \N__11923\,
            PADIN => \N__11922\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11915\,
            DIN => \N__11914\,
            DOUT => \N__11913\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11915\,
            PADOUT => \N__11914\,
            PADIN => \N__11913\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11906\,
            DIN => \N__11905\,
            DOUT => \N__11904\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11906\,
            PADOUT => \N__11905\,
            PADIN => \N__11904\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11897\,
            DIN => \N__11896\,
            DOUT => \N__11895\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11897\,
            PADOUT => \N__11896\,
            PADIN => \N__11895\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11888\,
            DIN => \N__11887\,
            DOUT => \N__11886\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11888\,
            PADOUT => \N__11887\,
            PADIN => \N__11886\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7567\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11879\,
            DIN => \N__11878\,
            DOUT => \N__11877\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11879\,
            PADOUT => \N__11878\,
            PADIN => \N__11877\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11870\,
            DIN => \N__11869\,
            DOUT => \N__11868\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11870\,
            PADOUT => \N__11869\,
            PADIN => \N__11868\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9118\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11861\,
            DIN => \N__11860\,
            DOUT => \N__11859\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11861\,
            PADOUT => \N__11860\,
            PADIN => \N__11859\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4612\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11852\,
            DIN => \N__11851\,
            DOUT => \N__11850\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11852\,
            PADOUT => \N__11851\,
            PADIN => \N__11850\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11843\,
            DIN => \N__11842\,
            DOUT => \N__11841\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11843\,
            PADOUT => \N__11842\,
            PADIN => \N__11841\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6463\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11834\,
            DIN => \N__11833\,
            DOUT => \N__11832\,
            PACKAGEPIN => \DA_wire\(0)
        );

    \DA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11834\,
            PADOUT => \N__11833\,
            PADIN => \N__11832\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6814\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11825\,
            DIN => \N__11824\,
            DOUT => \N__11823\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11825\,
            PADOUT => \N__11824\,
            PADIN => \N__11823\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8464\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11816\,
            DIN => \N__11815\,
            DOUT => \N__11814\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11816\,
            PADOUT => \N__11815\,
            PADIN => \N__11814\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11807\,
            DIN => \N__11806\,
            DOUT => \N__11805\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11807\,
            PADOUT => \N__11806\,
            PADIN => \N__11805\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11798\,
            DIN => \N__11797\,
            DOUT => \N__11796\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11798\,
            PADOUT => \N__11797\,
            PADIN => \N__11796\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11789\,
            DIN => \N__11788\,
            DOUT => \N__11787\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11789\,
            PADOUT => \N__11788\,
            PADIN => \N__11787\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11780\,
            DIN => \N__11779\,
            DOUT => \N__11778\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11780\,
            PADOUT => \N__11779\,
            PADIN => \N__11778\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7075\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11771\,
            DIN => \N__11770\,
            DOUT => \N__11769\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11771\,
            PADOUT => \N__11770\,
            PADIN => \N__11769\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11762\,
            DIN => \N__11761\,
            DOUT => \N__11760\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11762\,
            PADOUT => \N__11761\,
            PADIN => \N__11760\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8141\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11753\,
            DIN => \N__11752\,
            DOUT => \N__11751\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11753\,
            PADOUT => \N__11752\,
            PADIN => \N__11751\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8824\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11744\,
            DIN => \N__11743\,
            DOUT => \N__11742\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11744\,
            PADOUT => \N__11743\,
            PADIN => \N__11742\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11179\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11735\,
            DIN => \N__11734\,
            DOUT => \N__11733\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11735\,
            PADOUT => \N__11734\,
            PADIN => \N__11733\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8404\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11726\,
            DIN => \N__11725\,
            DOUT => \N__11724\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11726\,
            PADOUT => \N__11725\,
            PADIN => \N__11724\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8491\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11717\,
            DIN => \N__11716\,
            DOUT => \N__11715\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11717\,
            PADOUT => \N__11716\,
            PADIN => \N__11715\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6462\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11708\,
            DIN => \N__11707\,
            DOUT => \N__11706\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11708\,
            PADOUT => \N__11707\,
            PADIN => \N__11706\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11699\,
            DIN => \N__11698\,
            DOUT => \N__11697\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11699\,
            PADOUT => \N__11698\,
            PADIN => \N__11697\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11690\,
            DIN => \N__11689\,
            DOUT => \N__11688\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11690\,
            PADOUT => \N__11689\,
            PADIN => \N__11688\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9868\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11681\,
            DIN => \N__11680\,
            DOUT => \N__11679\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11681\,
            PADOUT => \N__11680\,
            PADIN => \N__11679\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8383\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11672\,
            DIN => \N__11671\,
            DOUT => \N__11670\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11672\,
            PADOUT => \N__11671\,
            PADIN => \N__11670\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5743\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11663\,
            DIN => \N__11662\,
            DOUT => \N__11661\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11663\,
            PADOUT => \N__11662\,
            PADIN => \N__11661\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9256\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11654\,
            DIN => \N__11653\,
            DOUT => \N__11652\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11654\,
            PADOUT => \N__11653\,
            PADIN => \N__11652\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11645\,
            DIN => \N__11644\,
            DOUT => \N__11643\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11645\,
            PADOUT => \N__11644\,
            PADIN => \N__11643\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11636\,
            DIN => \N__11635\,
            DOUT => \N__11634\,
            PACKAGEPIN => \DA_wire\(2)
        );

    \DA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11636\,
            PADOUT => \N__11635\,
            PADIN => \N__11634\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7414\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11627\,
            DIN => \N__11626\,
            DOUT => \N__11625\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11627\,
            PADOUT => \N__11626\,
            PADIN => \N__11625\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11618\,
            DIN => \N__11617\,
            DOUT => \N__11616\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11618\,
            PADOUT => \N__11617\,
            PADIN => \N__11616\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11609\,
            DIN => \N__11608\,
            DOUT => \N__11607\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11609\,
            PADOUT => \N__11608\,
            PADIN => \N__11607\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7063\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11600\,
            DIN => \N__11599\,
            DOUT => \N__11598\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11600\,
            PADOUT => \N__11599\,
            PADIN => \N__11598\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11122\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11591\,
            DIN => \N__11590\,
            DOUT => \N__11589\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11591\,
            PADOUT => \N__11590\,
            PADIN => \N__11589\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11582\,
            DIN => \N__11581\,
            DOUT => \N__11580\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11582\,
            PADOUT => \N__11581\,
            PADIN => \N__11580\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9694\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11573\,
            DIN => \N__11572\,
            DOUT => \N__11571\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11573\,
            PADOUT => \N__11572\,
            PADIN => \N__11571\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7609\,
            DIN0 => OPEN,
            DOUT0 => \N__7666\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11564\,
            DIN => \N__11563\,
            DOUT => \N__11562\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11564\,
            PADOUT => \N__11563\,
            PADIN => \N__11562\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7453\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11555\,
            DIN => \N__11554\,
            DOUT => \N__11553\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11555\,
            PADOUT => \N__11554\,
            PADIN => \N__11553\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11546\,
            DIN => \N__11545\,
            DOUT => \N__11544\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11546\,
            PADOUT => \N__11545\,
            PADIN => \N__11544\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11537\,
            DIN => \N__11536\,
            DOUT => \N__11535\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11537\,
            PADOUT => \N__11536\,
            PADIN => \N__11535\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8569\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11528\,
            DIN => \N__11527\,
            DOUT => \N__11526\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11528\,
            PADOUT => \N__11527\,
            PADIN => \N__11526\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4273\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11519\,
            DIN => \N__11518\,
            DOUT => \N__11517\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11519\,
            PADOUT => \N__11518\,
            PADIN => \N__11517\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11510\,
            DIN => \N__11509\,
            DOUT => \N__11508\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11510\,
            PADOUT => \N__11509\,
            PADIN => \N__11508\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11501\,
            DIN => \N__11500\,
            DOUT => \N__11499\,
            PACKAGEPIN => \DA_wire\(1)
        );

    \DA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11501\,
            PADOUT => \N__11500\,
            PADIN => \N__11499\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7717\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11492\,
            DIN => \N__11491\,
            DOUT => \N__11490\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11492\,
            PADOUT => \N__11491\,
            PADIN => \N__11490\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11483\,
            DIN => \N__11482\,
            DOUT => \N__11481\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11483\,
            PADOUT => \N__11482\,
            PADIN => \N__11481\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11474\,
            DIN => \N__11473\,
            DOUT => \N__11472\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11474\,
            PADOUT => \N__11473\,
            PADIN => \N__11472\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8215\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11465\,
            DIN => \N__11464\,
            DOUT => \N__11463\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11465\,
            PADOUT => \N__11464\,
            PADIN => \N__11463\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9358\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11456\,
            DIN => \N__11455\,
            DOUT => \N__11454\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11456\,
            PADOUT => \N__11455\,
            PADIN => \N__11454\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11107\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11447\,
            DIN => \N__11446\,
            DOUT => \N__11445\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11447\,
            PADOUT => \N__11446\,
            PADIN => \N__11445\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4216\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11438\,
            DIN => \N__11437\,
            DOUT => \N__11436\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11438\,
            PADOUT => \N__11437\,
            PADIN => \N__11436\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11429\,
            DIN => \N__11428\,
            DOUT => \N__11427\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11429\,
            PADOUT => \N__11428\,
            PADIN => \N__11427\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11420\,
            DIN => \N__11419\,
            DOUT => \N__11418\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11420\,
            PADOUT => \N__11419\,
            PADIN => \N__11418\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8611\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11411\,
            DIN => \N__11410\,
            DOUT => \N__11409\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11411\,
            PADOUT => \N__11410\,
            PADIN => \N__11409\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11402\,
            DIN => \N__11401\,
            DOUT => \N__11400\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11402\,
            PADOUT => \N__11401\,
            PADIN => \N__11400\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11393\,
            DIN => \N__11392\,
            DOUT => \N__11391\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11393\,
            PADOUT => \N__11392\,
            PADIN => \N__11391\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5692\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11384\,
            DIN => \N__11383\,
            DOUT => \N__11382\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11384\,
            PADOUT => \N__11383\,
            PADIN => \N__11382\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9313\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11375\,
            DIN => \N__11374\,
            DOUT => \N__11373\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11375\,
            PADOUT => \N__11374\,
            PADIN => \N__11373\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8149\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11366\,
            DIN => \N__11365\,
            DOUT => \N__11364\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11366\,
            PADOUT => \N__11365\,
            PADIN => \N__11364\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11357\,
            DIN => \N__11356\,
            DOUT => \N__11355\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11357\,
            PADOUT => \N__11356\,
            PADIN => \N__11355\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8148\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11348\,
            DIN => \N__11347\,
            DOUT => \N__11346\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11348\,
            PADOUT => \N__11347\,
            PADIN => \N__11346\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4252\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2768\ : InMux
    port map (
            O => \N__11329\,
            I => \N__11326\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__11326\,
            I => \N__11321\
        );

    \I__2766\ : InMux
    port map (
            O => \N__11325\,
            I => \N__11317\
        );

    \I__2765\ : InMux
    port map (
            O => \N__11324\,
            I => \N__11313\
        );

    \I__2764\ : Span4Mux_v
    port map (
            O => \N__11321\,
            I => \N__11310\
        );

    \I__2763\ : InMux
    port map (
            O => \N__11320\,
            I => \N__11307\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__11317\,
            I => \N__11304\
        );

    \I__2761\ : InMux
    port map (
            O => \N__11316\,
            I => \N__11301\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__11313\,
            I => \N__11297\
        );

    \I__2759\ : Span4Mux_v
    port map (
            O => \N__11310\,
            I => \N__11294\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__11307\,
            I => \N__11289\
        );

    \I__2757\ : Sp12to4
    port map (
            O => \N__11304\,
            I => \N__11289\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__11301\,
            I => \N__11286\
        );

    \I__2755\ : InMux
    port map (
            O => \N__11300\,
            I => \N__11283\
        );

    \I__2754\ : Span12Mux_h
    port map (
            O => \N__11297\,
            I => \N__11280\
        );

    \I__2753\ : Sp12to4
    port map (
            O => \N__11294\,
            I => \N__11275\
        );

    \I__2752\ : Span12Mux_v
    port map (
            O => \N__11289\,
            I => \N__11275\
        );

    \I__2751\ : Span12Mux_h
    port map (
            O => \N__11286\,
            I => \N__11270\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__11283\,
            I => \N__11270\
        );

    \I__2749\ : Span12Mux_v
    port map (
            O => \N__11280\,
            I => \N__11267\
        );

    \I__2748\ : Span12Mux_h
    port map (
            O => \N__11275\,
            I => \N__11262\
        );

    \I__2747\ : Span12Mux_v
    port map (
            O => \N__11270\,
            I => \N__11262\
        );

    \I__2746\ : Odrv12
    port map (
            O => \N__11267\,
            I => \CASLn_c\
        );

    \I__2745\ : Odrv12
    port map (
            O => \N__11262\,
            I => \CASLn_c\
        );

    \I__2744\ : InMux
    port map (
            O => \N__11257\,
            I => \N__11252\
        );

    \I__2743\ : InMux
    port map (
            O => \N__11256\,
            I => \N__11249\
        );

    \I__2742\ : InMux
    port map (
            O => \N__11255\,
            I => \N__11246\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__11252\,
            I => \N__11242\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__11249\,
            I => \N__11237\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__11246\,
            I => \N__11237\
        );

    \I__2738\ : InMux
    port map (
            O => \N__11245\,
            I => \N__11234\
        );

    \I__2737\ : Span4Mux_v
    port map (
            O => \N__11242\,
            I => \N__11231\
        );

    \I__2736\ : Span4Mux_h
    port map (
            O => \N__11237\,
            I => \N__11228\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__11234\,
            I => \N__11225\
        );

    \I__2734\ : Span4Mux_v
    port map (
            O => \N__11231\,
            I => \N__11219\
        );

    \I__2733\ : Span4Mux_h
    port map (
            O => \N__11228\,
            I => \N__11219\
        );

    \I__2732\ : Span4Mux_v
    port map (
            O => \N__11225\,
            I => \N__11215\
        );

    \I__2731\ : InMux
    port map (
            O => \N__11224\,
            I => \N__11212\
        );

    \I__2730\ : Span4Mux_h
    port map (
            O => \N__11219\,
            I => \N__11209\
        );

    \I__2729\ : InMux
    port map (
            O => \N__11218\,
            I => \N__11206\
        );

    \I__2728\ : Sp12to4
    port map (
            O => \N__11215\,
            I => \N__11201\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__11212\,
            I => \N__11201\
        );

    \I__2726\ : Span4Mux_h
    port map (
            O => \N__11209\,
            I => \N__11196\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__11206\,
            I => \N__11196\
        );

    \I__2724\ : Span12Mux_h
    port map (
            O => \N__11201\,
            I => \N__11193\
        );

    \I__2723\ : Span4Mux_h
    port map (
            O => \N__11196\,
            I => \N__11190\
        );

    \I__2722\ : Span12Mux_v
    port map (
            O => \N__11193\,
            I => \N__11187\
        );

    \I__2721\ : Span4Mux_v
    port map (
            O => \N__11190\,
            I => \N__11184\
        );

    \I__2720\ : Odrv12
    port map (
            O => \N__11187\,
            I => \CASUn_c\
        );

    \I__2719\ : Odrv4
    port map (
            O => \N__11184\,
            I => \CASUn_c\
        );

    \I__2718\ : IoInMux
    port map (
            O => \N__11179\,
            I => \N__11176\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__11176\,
            I => \N__11173\
        );

    \I__2716\ : Span12Mux_s7_v
    port map (
            O => \N__11173\,
            I => \N__11170\
        );

    \I__2715\ : Odrv12
    port map (
            O => \N__11170\,
            I => \DRDENn_c\
        );

    \I__2714\ : InMux
    port map (
            O => \N__11167\,
            I => \N__11164\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__11164\,
            I => \N__11161\
        );

    \I__2712\ : Odrv4
    port map (
            O => \N__11161\,
            I => \U712_BYTE_ENABLE.N_561\
        );

    \I__2711\ : InMux
    port map (
            O => \N__11158\,
            I => \N__11152\
        );

    \I__2710\ : InMux
    port map (
            O => \N__11157\,
            I => \N__11149\
        );

    \I__2709\ : CascadeMux
    port map (
            O => \N__11156\,
            I => \N__11146\
        );

    \I__2708\ : CascadeMux
    port map (
            O => \N__11155\,
            I => \N__11143\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__11152\,
            I => \N__11138\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__11149\,
            I => \N__11138\
        );

    \I__2705\ : InMux
    port map (
            O => \N__11146\,
            I => \N__11133\
        );

    \I__2704\ : InMux
    port map (
            O => \N__11143\,
            I => \N__11133\
        );

    \I__2703\ : Span4Mux_v
    port map (
            O => \N__11138\,
            I => \N__11130\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__11133\,
            I => \N__11127\
        );

    \I__2701\ : Odrv4
    port map (
            O => \N__11130\,
            I => \U712_BYTE_ENABLE.N_397_i\
        );

    \I__2700\ : Odrv4
    port map (
            O => \N__11127\,
            I => \U712_BYTE_ENABLE.N_397_i\
        );

    \I__2699\ : IoInMux
    port map (
            O => \N__11122\,
            I => \N__11119\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__11119\,
            I => \N__11116\
        );

    \I__2697\ : Span4Mux_s0_v
    port map (
            O => \N__11116\,
            I => \N__11113\
        );

    \I__2696\ : Span4Mux_v
    port map (
            O => \N__11113\,
            I => \N__11110\
        );

    \I__2695\ : Odrv4
    port map (
            O => \N__11110\,
            I => \N_130_i\
        );

    \I__2694\ : IoInMux
    port map (
            O => \N__11107\,
            I => \N__11104\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__11104\,
            I => \N__11101\
        );

    \I__2692\ : IoSpan4Mux
    port map (
            O => \N__11101\,
            I => \N__11098\
        );

    \I__2691\ : Span4Mux_s2_v
    port map (
            O => \N__11098\,
            I => \N__11095\
        );

    \I__2690\ : Span4Mux_v
    port map (
            O => \N__11095\,
            I => \N__11092\
        );

    \I__2689\ : Odrv4
    port map (
            O => \N__11092\,
            I => \N_127_i\
        );

    \I__2688\ : InMux
    port map (
            O => \N__11089\,
            I => \N__11076\
        );

    \I__2687\ : InMux
    port map (
            O => \N__11088\,
            I => \N__11076\
        );

    \I__2686\ : InMux
    port map (
            O => \N__11087\,
            I => \N__11076\
        );

    \I__2685\ : InMux
    port map (
            O => \N__11086\,
            I => \N__11071\
        );

    \I__2684\ : InMux
    port map (
            O => \N__11085\,
            I => \N__11071\
        );

    \I__2683\ : InMux
    port map (
            O => \N__11084\,
            I => \N__11066\
        );

    \I__2682\ : InMux
    port map (
            O => \N__11083\,
            I => \N__11066\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__11076\,
            I => \N__11060\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__11071\,
            I => \N__11060\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__11066\,
            I => \N__11057\
        );

    \I__2678\ : InMux
    port map (
            O => \N__11065\,
            I => \N__11054\
        );

    \I__2677\ : Span4Mux_v
    port map (
            O => \N__11060\,
            I => \N__11048\
        );

    \I__2676\ : Span4Mux_v
    port map (
            O => \N__11057\,
            I => \N__11048\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__11054\,
            I => \N__11045\
        );

    \I__2674\ : InMux
    port map (
            O => \N__11053\,
            I => \N__11042\
        );

    \I__2673\ : Span4Mux_h
    port map (
            O => \N__11048\,
            I => \N__11039\
        );

    \I__2672\ : Span4Mux_v
    port map (
            O => \N__11045\,
            I => \N__11036\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__11042\,
            I => \N__11033\
        );

    \I__2670\ : Sp12to4
    port map (
            O => \N__11039\,
            I => \N__11026\
        );

    \I__2669\ : Sp12to4
    port map (
            O => \N__11036\,
            I => \N__11026\
        );

    \I__2668\ : Span12Mux_v
    port map (
            O => \N__11033\,
            I => \N__11026\
        );

    \I__2667\ : Span12Mux_h
    port map (
            O => \N__11026\,
            I => \N__11023\
        );

    \I__2666\ : Odrv12
    port map (
            O => \N__11023\,
            I => \A_c_0\
        );

    \I__2665\ : InMux
    port map (
            O => \N__11020\,
            I => \N__11013\
        );

    \I__2664\ : InMux
    port map (
            O => \N__11019\,
            I => \N__11013\
        );

    \I__2663\ : InMux
    port map (
            O => \N__11018\,
            I => \N__11007\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__11013\,
            I => \N__11002\
        );

    \I__2661\ : InMux
    port map (
            O => \N__11012\,
            I => \N__10995\
        );

    \I__2660\ : InMux
    port map (
            O => \N__11011\,
            I => \N__10995\
        );

    \I__2659\ : InMux
    port map (
            O => \N__11010\,
            I => \N__10995\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__11007\,
            I => \N__10992\
        );

    \I__2657\ : InMux
    port map (
            O => \N__11006\,
            I => \N__10989\
        );

    \I__2656\ : InMux
    port map (
            O => \N__11005\,
            I => \N__10986\
        );

    \I__2655\ : Span4Mux_v
    port map (
            O => \N__11002\,
            I => \N__10983\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__10995\,
            I => \N__10980\
        );

    \I__2653\ : Span4Mux_v
    port map (
            O => \N__10992\,
            I => \N__10977\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__10989\,
            I => \N__10974\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__10986\,
            I => \N__10971\
        );

    \I__2650\ : Span4Mux_v
    port map (
            O => \N__10983\,
            I => \N__10966\
        );

    \I__2649\ : Span4Mux_v
    port map (
            O => \N__10980\,
            I => \N__10966\
        );

    \I__2648\ : Span4Mux_v
    port map (
            O => \N__10977\,
            I => \N__10961\
        );

    \I__2647\ : Span4Mux_v
    port map (
            O => \N__10974\,
            I => \N__10961\
        );

    \I__2646\ : Span12Mux_v
    port map (
            O => \N__10971\,
            I => \N__10958\
        );

    \I__2645\ : Sp12to4
    port map (
            O => \N__10966\,
            I => \N__10953\
        );

    \I__2644\ : Sp12to4
    port map (
            O => \N__10961\,
            I => \N__10953\
        );

    \I__2643\ : Span12Mux_h
    port map (
            O => \N__10958\,
            I => \N__10950\
        );

    \I__2642\ : Span12Mux_h
    port map (
            O => \N__10953\,
            I => \N__10947\
        );

    \I__2641\ : Odrv12
    port map (
            O => \N__10950\,
            I => \A_c_1\
        );

    \I__2640\ : Odrv12
    port map (
            O => \N__10947\,
            I => \A_c_1\
        );

    \I__2639\ : InMux
    port map (
            O => \N__10942\,
            I => \N__10937\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__10941\,
            I => \N__10933\
        );

    \I__2637\ : CascadeMux
    port map (
            O => \N__10940\,
            I => \N__10930\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__10937\,
            I => \N__10924\
        );

    \I__2635\ : InMux
    port map (
            O => \N__10936\,
            I => \N__10917\
        );

    \I__2634\ : InMux
    port map (
            O => \N__10933\,
            I => \N__10917\
        );

    \I__2633\ : InMux
    port map (
            O => \N__10930\,
            I => \N__10917\
        );

    \I__2632\ : CascadeMux
    port map (
            O => \N__10929\,
            I => \N__10914\
        );

    \I__2631\ : CascadeMux
    port map (
            O => \N__10928\,
            I => \N__10911\
        );

    \I__2630\ : CascadeMux
    port map (
            O => \N__10927\,
            I => \N__10908\
        );

    \I__2629\ : Span4Mux_h
    port map (
            O => \N__10924\,
            I => \N__10905\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__10917\,
            I => \N__10902\
        );

    \I__2627\ : InMux
    port map (
            O => \N__10914\,
            I => \N__10897\
        );

    \I__2626\ : InMux
    port map (
            O => \N__10911\,
            I => \N__10897\
        );

    \I__2625\ : InMux
    port map (
            O => \N__10908\,
            I => \N__10894\
        );

    \I__2624\ : Span4Mux_v
    port map (
            O => \N__10905\,
            I => \N__10885\
        );

    \I__2623\ : Span4Mux_h
    port map (
            O => \N__10902\,
            I => \N__10885\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__10897\,
            I => \N__10885\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__10894\,
            I => \N__10885\
        );

    \I__2620\ : Span4Mux_h
    port map (
            O => \N__10885\,
            I => \N__10882\
        );

    \I__2619\ : Span4Mux_v
    port map (
            O => \N__10882\,
            I => \N__10879\
        );

    \I__2618\ : Sp12to4
    port map (
            O => \N__10879\,
            I => \N__10876\
        );

    \I__2617\ : Span12Mux_h
    port map (
            O => \N__10876\,
            I => \N__10873\
        );

    \I__2616\ : Odrv12
    port map (
            O => \N__10873\,
            I => \SIZ_c_0\
        );

    \I__2615\ : InMux
    port map (
            O => \N__10870\,
            I => \N__10865\
        );

    \I__2614\ : InMux
    port map (
            O => \N__10869\,
            I => \N__10862\
        );

    \I__2613\ : CascadeMux
    port map (
            O => \N__10868\,
            I => \N__10859\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__10865\,
            I => \N__10854\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__10862\,
            I => \N__10851\
        );

    \I__2610\ : InMux
    port map (
            O => \N__10859\,
            I => \N__10844\
        );

    \I__2609\ : InMux
    port map (
            O => \N__10858\,
            I => \N__10844\
        );

    \I__2608\ : InMux
    port map (
            O => \N__10857\,
            I => \N__10844\
        );

    \I__2607\ : Span4Mux_h
    port map (
            O => \N__10854\,
            I => \N__10836\
        );

    \I__2606\ : Span4Mux_v
    port map (
            O => \N__10851\,
            I => \N__10836\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__10844\,
            I => \N__10833\
        );

    \I__2604\ : InMux
    port map (
            O => \N__10843\,
            I => \N__10828\
        );

    \I__2603\ : InMux
    port map (
            O => \N__10842\,
            I => \N__10828\
        );

    \I__2602\ : InMux
    port map (
            O => \N__10841\,
            I => \N__10825\
        );

    \I__2601\ : Span4Mux_v
    port map (
            O => \N__10836\,
            I => \N__10822\
        );

    \I__2600\ : Span4Mux_h
    port map (
            O => \N__10833\,
            I => \N__10815\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__10828\,
            I => \N__10815\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__10825\,
            I => \N__10815\
        );

    \I__2597\ : Span4Mux_v
    port map (
            O => \N__10822\,
            I => \N__10812\
        );

    \I__2596\ : Sp12to4
    port map (
            O => \N__10815\,
            I => \N__10809\
        );

    \I__2595\ : Sp12to4
    port map (
            O => \N__10812\,
            I => \N__10804\
        );

    \I__2594\ : Span12Mux_v
    port map (
            O => \N__10809\,
            I => \N__10804\
        );

    \I__2593\ : Span12Mux_h
    port map (
            O => \N__10804\,
            I => \N__10801\
        );

    \I__2592\ : Odrv12
    port map (
            O => \N__10801\,
            I => \SIZ_c_1\
        );

    \I__2591\ : IoInMux
    port map (
            O => \N__10798\,
            I => \N__10795\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__10795\,
            I => \N__10792\
        );

    \I__2589\ : Span4Mux_s3_v
    port map (
            O => \N__10792\,
            I => \N__10789\
        );

    \I__2588\ : Odrv4
    port map (
            O => \N__10789\,
            I => \N_128_i\
        );

    \I__2587\ : InMux
    port map (
            O => \N__10786\,
            I => \N__10782\
        );

    \I__2586\ : InMux
    port map (
            O => \N__10785\,
            I => \N__10779\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__10782\,
            I => \N__10773\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__10779\,
            I => \N__10773\
        );

    \I__2583\ : InMux
    port map (
            O => \N__10778\,
            I => \N__10770\
        );

    \I__2582\ : Span4Mux_h
    port map (
            O => \N__10773\,
            I => \N__10764\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__10770\,
            I => \N__10764\
        );

    \I__2580\ : InMux
    port map (
            O => \N__10769\,
            I => \N__10761\
        );

    \I__2579\ : Span4Mux_v
    port map (
            O => \N__10764\,
            I => \N__10758\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__10761\,
            I => \N__10755\
        );

    \I__2577\ : Span4Mux_v
    port map (
            O => \N__10758\,
            I => \N__10752\
        );

    \I__2576\ : Span4Mux_h
    port map (
            O => \N__10755\,
            I => \N__10749\
        );

    \I__2575\ : Span4Mux_h
    port map (
            O => \N__10752\,
            I => \N__10746\
        );

    \I__2574\ : Sp12to4
    port map (
            O => \N__10749\,
            I => \N__10743\
        );

    \I__2573\ : Sp12to4
    port map (
            O => \N__10746\,
            I => \N__10738\
        );

    \I__2572\ : Span12Mux_v
    port map (
            O => \N__10743\,
            I => \N__10738\
        );

    \I__2571\ : Odrv12
    port map (
            O => \N__10738\,
            I => \DRA_c_6\
        );

    \I__2570\ : InMux
    port map (
            O => \N__10735\,
            I => \N__10732\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__10732\,
            I => \N__10727\
        );

    \I__2568\ : InMux
    port map (
            O => \N__10731\,
            I => \N__10724\
        );

    \I__2567\ : InMux
    port map (
            O => \N__10730\,
            I => \N__10721\
        );

    \I__2566\ : Span4Mux_h
    port map (
            O => \N__10727\,
            I => \N__10715\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__10724\,
            I => \N__10715\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__10721\,
            I => \N__10712\
        );

    \I__2563\ : InMux
    port map (
            O => \N__10720\,
            I => \N__10709\
        );

    \I__2562\ : Span4Mux_v
    port map (
            O => \N__10715\,
            I => \N__10706\
        );

    \I__2561\ : Sp12to4
    port map (
            O => \N__10712\,
            I => \N__10701\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__10709\,
            I => \N__10701\
        );

    \I__2559\ : Sp12to4
    port map (
            O => \N__10706\,
            I => \N__10698\
        );

    \I__2558\ : Span12Mux_v
    port map (
            O => \N__10701\,
            I => \N__10695\
        );

    \I__2557\ : Span12Mux_h
    port map (
            O => \N__10698\,
            I => \N__10692\
        );

    \I__2556\ : Span12Mux_h
    port map (
            O => \N__10695\,
            I => \N__10689\
        );

    \I__2555\ : Odrv12
    port map (
            O => \N__10692\,
            I => \DRA_c_7\
        );

    \I__2554\ : Odrv12
    port map (
            O => \N__10689\,
            I => \DRA_c_7\
        );

    \I__2553\ : InMux
    port map (
            O => \N__10684\,
            I => \N__10681\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__10681\,
            I => \N__10678\
        );

    \I__2551\ : Odrv4
    port map (
            O => \N__10678\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2550\ : InMux
    port map (
            O => \N__10675\,
            I => \N__10668\
        );

    \I__2549\ : InMux
    port map (
            O => \N__10674\,
            I => \N__10668\
        );

    \I__2548\ : InMux
    port map (
            O => \N__10673\,
            I => \N__10664\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__10668\,
            I => \N__10661\
        );

    \I__2546\ : InMux
    port map (
            O => \N__10667\,
            I => \N__10658\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__10664\,
            I => \N__10655\
        );

    \I__2544\ : Span4Mux_v
    port map (
            O => \N__10661\,
            I => \N__10652\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__10658\,
            I => \N__10649\
        );

    \I__2542\ : Span12Mux_v
    port map (
            O => \N__10655\,
            I => \N__10646\
        );

    \I__2541\ : Span4Mux_h
    port map (
            O => \N__10652\,
            I => \N__10641\
        );

    \I__2540\ : Span4Mux_v
    port map (
            O => \N__10649\,
            I => \N__10641\
        );

    \I__2539\ : Span12Mux_h
    port map (
            O => \N__10646\,
            I => \N__10638\
        );

    \I__2538\ : Sp12to4
    port map (
            O => \N__10641\,
            I => \N__10635\
        );

    \I__2537\ : Odrv12
    port map (
            O => \N__10638\,
            I => \DRA_c_8\
        );

    \I__2536\ : Odrv12
    port map (
            O => \N__10635\,
            I => \DRA_c_8\
        );

    \I__2535\ : InMux
    port map (
            O => \N__10630\,
            I => \N__10627\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__10627\,
            I => \N__10624\
        );

    \I__2533\ : Span4Mux_v
    port map (
            O => \N__10624\,
            I => \N__10621\
        );

    \I__2532\ : Odrv4
    port map (
            O => \N__10621\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__2531\ : InMux
    port map (
            O => \N__10618\,
            I => \N__10606\
        );

    \I__2530\ : InMux
    port map (
            O => \N__10617\,
            I => \N__10606\
        );

    \I__2529\ : InMux
    port map (
            O => \N__10616\,
            I => \N__10606\
        );

    \I__2528\ : InMux
    port map (
            O => \N__10615\,
            I => \N__10603\
        );

    \I__2527\ : InMux
    port map (
            O => \N__10614\,
            I => \N__10600\
        );

    \I__2526\ : InMux
    port map (
            O => \N__10613\,
            I => \N__10588\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__10606\,
            I => \N__10584\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__10603\,
            I => \N__10579\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__10600\,
            I => \N__10579\
        );

    \I__2522\ : InMux
    port map (
            O => \N__10599\,
            I => \N__10576\
        );

    \I__2521\ : InMux
    port map (
            O => \N__10598\,
            I => \N__10573\
        );

    \I__2520\ : InMux
    port map (
            O => \N__10597\,
            I => \N__10570\
        );

    \I__2519\ : InMux
    port map (
            O => \N__10596\,
            I => \N__10562\
        );

    \I__2518\ : InMux
    port map (
            O => \N__10595\,
            I => \N__10562\
        );

    \I__2517\ : InMux
    port map (
            O => \N__10594\,
            I => \N__10562\
        );

    \I__2516\ : InMux
    port map (
            O => \N__10593\,
            I => \N__10559\
        );

    \I__2515\ : InMux
    port map (
            O => \N__10592\,
            I => \N__10556\
        );

    \I__2514\ : CascadeMux
    port map (
            O => \N__10591\,
            I => \N__10552\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__10588\,
            I => \N__10549\
        );

    \I__2512\ : InMux
    port map (
            O => \N__10587\,
            I => \N__10546\
        );

    \I__2511\ : Span4Mux_v
    port map (
            O => \N__10584\,
            I => \N__10535\
        );

    \I__2510\ : Span4Mux_v
    port map (
            O => \N__10579\,
            I => \N__10535\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__10576\,
            I => \N__10535\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__10573\,
            I => \N__10535\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__10570\,
            I => \N__10535\
        );

    \I__2506\ : InMux
    port map (
            O => \N__10569\,
            I => \N__10532\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__10562\,
            I => \N__10527\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__10559\,
            I => \N__10522\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__10556\,
            I => \N__10522\
        );

    \I__2502\ : InMux
    port map (
            O => \N__10555\,
            I => \N__10518\
        );

    \I__2501\ : InMux
    port map (
            O => \N__10552\,
            I => \N__10515\
        );

    \I__2500\ : Span4Mux_v
    port map (
            O => \N__10549\,
            I => \N__10512\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__10546\,
            I => \N__10509\
        );

    \I__2498\ : Span4Mux_v
    port map (
            O => \N__10535\,
            I => \N__10506\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__10532\,
            I => \N__10503\
        );

    \I__2496\ : InMux
    port map (
            O => \N__10531\,
            I => \N__10498\
        );

    \I__2495\ : InMux
    port map (
            O => \N__10530\,
            I => \N__10498\
        );

    \I__2494\ : Span4Mux_h
    port map (
            O => \N__10527\,
            I => \N__10493\
        );

    \I__2493\ : Span4Mux_v
    port map (
            O => \N__10522\,
            I => \N__10493\
        );

    \I__2492\ : InMux
    port map (
            O => \N__10521\,
            I => \N__10490\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__10518\,
            I => \N__10485\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__10515\,
            I => \N__10485\
        );

    \I__2489\ : Span4Mux_h
    port map (
            O => \N__10512\,
            I => \N__10480\
        );

    \I__2488\ : Span4Mux_v
    port map (
            O => \N__10509\,
            I => \N__10480\
        );

    \I__2487\ : Span4Mux_h
    port map (
            O => \N__10506\,
            I => \N__10475\
        );

    \I__2486\ : Span4Mux_v
    port map (
            O => \N__10503\,
            I => \N__10475\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__10498\,
            I => \N__10468\
        );

    \I__2484\ : Sp12to4
    port map (
            O => \N__10493\,
            I => \N__10468\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__10490\,
            I => \N__10468\
        );

    \I__2482\ : Sp12to4
    port map (
            O => \N__10485\,
            I => \N__10465\
        );

    \I__2481\ : Sp12to4
    port map (
            O => \N__10480\,
            I => \N__10460\
        );

    \I__2480\ : Sp12to4
    port map (
            O => \N__10475\,
            I => \N__10460\
        );

    \I__2479\ : Span12Mux_h
    port map (
            O => \N__10468\,
            I => \N__10457\
        );

    \I__2478\ : Span12Mux_v
    port map (
            O => \N__10465\,
            I => \N__10454\
        );

    \I__2477\ : Span12Mux_h
    port map (
            O => \N__10460\,
            I => \N__10451\
        );

    \I__2476\ : Span12Mux_v
    port map (
            O => \N__10457\,
            I => \N__10446\
        );

    \I__2475\ : Span12Mux_h
    port map (
            O => \N__10454\,
            I => \N__10446\
        );

    \I__2474\ : Span12Mux_v
    port map (
            O => \N__10451\,
            I => \N__10443\
        );

    \I__2473\ : Odrv12
    port map (
            O => \N__10446\,
            I => \AGNUS_REV_c\
        );

    \I__2472\ : Odrv12
    port map (
            O => \N__10443\,
            I => \AGNUS_REV_c\
        );

    \I__2471\ : InMux
    port map (
            O => \N__10438\,
            I => \N__10435\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__10435\,
            I => \N__10432\
        );

    \I__2469\ : Odrv12
    port map (
            O => \N__10432\,
            I => \RAS0n_c\
        );

    \I__2468\ : InMux
    port map (
            O => \N__10429\,
            I => \N__10425\
        );

    \I__2467\ : InMux
    port map (
            O => \N__10428\,
            I => \N__10422\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__10425\,
            I => \N__10418\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__10422\,
            I => \N__10415\
        );

    \I__2464\ : InMux
    port map (
            O => \N__10421\,
            I => \N__10412\
        );

    \I__2463\ : Span4Mux_v
    port map (
            O => \N__10418\,
            I => \N__10409\
        );

    \I__2462\ : Span4Mux_v
    port map (
            O => \N__10415\,
            I => \N__10404\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__10412\,
            I => \N__10404\
        );

    \I__2460\ : Span4Mux_v
    port map (
            O => \N__10409\,
            I => \N__10398\
        );

    \I__2459\ : Span4Mux_v
    port map (
            O => \N__10404\,
            I => \N__10398\
        );

    \I__2458\ : InMux
    port map (
            O => \N__10403\,
            I => \N__10395\
        );

    \I__2457\ : Sp12to4
    port map (
            O => \N__10398\,
            I => \N__10392\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__10395\,
            I => \N__10389\
        );

    \I__2455\ : Span12Mux_h
    port map (
            O => \N__10392\,
            I => \N__10386\
        );

    \I__2454\ : Span12Mux_v
    port map (
            O => \N__10389\,
            I => \N__10383\
        );

    \I__2453\ : Span12Mux_v
    port map (
            O => \N__10386\,
            I => \N__10380\
        );

    \I__2452\ : Span12Mux_v
    port map (
            O => \N__10383\,
            I => \N__10377\
        );

    \I__2451\ : Odrv12
    port map (
            O => \N__10380\,
            I => \DRA_c_9\
        );

    \I__2450\ : Odrv12
    port map (
            O => \N__10377\,
            I => \DRA_c_9\
        );

    \I__2449\ : InMux
    port map (
            O => \N__10372\,
            I => \N__10369\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__10369\,
            I => \N__10366\
        );

    \I__2447\ : Span4Mux_h
    port map (
            O => \N__10366\,
            I => \N__10363\
        );

    \I__2446\ : Span4Mux_h
    port map (
            O => \N__10363\,
            I => \N__10360\
        );

    \I__2445\ : Odrv4
    port map (
            O => \N__10360\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2444\ : ClkMux
    port map (
            O => \N__10357\,
            I => \N__10333\
        );

    \I__2443\ : ClkMux
    port map (
            O => \N__10356\,
            I => \N__10333\
        );

    \I__2442\ : ClkMux
    port map (
            O => \N__10355\,
            I => \N__10333\
        );

    \I__2441\ : ClkMux
    port map (
            O => \N__10354\,
            I => \N__10333\
        );

    \I__2440\ : ClkMux
    port map (
            O => \N__10353\,
            I => \N__10333\
        );

    \I__2439\ : ClkMux
    port map (
            O => \N__10352\,
            I => \N__10333\
        );

    \I__2438\ : ClkMux
    port map (
            O => \N__10351\,
            I => \N__10333\
        );

    \I__2437\ : ClkMux
    port map (
            O => \N__10350\,
            I => \N__10333\
        );

    \I__2436\ : GlobalMux
    port map (
            O => \N__10333\,
            I => \N__10330\
        );

    \I__2435\ : gio2CtrlBuf
    port map (
            O => \N__10330\,
            I => \C3_c_g\
        );

    \I__2434\ : CEMux
    port map (
            O => \N__10327\,
            I => \N__10285\
        );

    \I__2433\ : CEMux
    port map (
            O => \N__10326\,
            I => \N__10285\
        );

    \I__2432\ : CEMux
    port map (
            O => \N__10325\,
            I => \N__10285\
        );

    \I__2431\ : CEMux
    port map (
            O => \N__10324\,
            I => \N__10285\
        );

    \I__2430\ : CEMux
    port map (
            O => \N__10323\,
            I => \N__10285\
        );

    \I__2429\ : CEMux
    port map (
            O => \N__10322\,
            I => \N__10285\
        );

    \I__2428\ : CEMux
    port map (
            O => \N__10321\,
            I => \N__10285\
        );

    \I__2427\ : CEMux
    port map (
            O => \N__10320\,
            I => \N__10285\
        );

    \I__2426\ : CEMux
    port map (
            O => \N__10319\,
            I => \N__10285\
        );

    \I__2425\ : CEMux
    port map (
            O => \N__10318\,
            I => \N__10285\
        );

    \I__2424\ : CEMux
    port map (
            O => \N__10317\,
            I => \N__10285\
        );

    \I__2423\ : CEMux
    port map (
            O => \N__10316\,
            I => \N__10285\
        );

    \I__2422\ : CEMux
    port map (
            O => \N__10315\,
            I => \N__10285\
        );

    \I__2421\ : CEMux
    port map (
            O => \N__10314\,
            I => \N__10285\
        );

    \I__2420\ : GlobalMux
    port map (
            O => \N__10285\,
            I => \N__10282\
        );

    \I__2419\ : gio2CtrlBuf
    port map (
            O => \N__10282\,
            I => \DBRn_c_i_0_g\
        );

    \I__2418\ : InMux
    port map (
            O => \N__10279\,
            I => \N__10272\
        );

    \I__2417\ : InMux
    port map (
            O => \N__10278\,
            I => \N__10269\
        );

    \I__2416\ : InMux
    port map (
            O => \N__10277\,
            I => \N__10266\
        );

    \I__2415\ : InMux
    port map (
            O => \N__10276\,
            I => \N__10261\
        );

    \I__2414\ : InMux
    port map (
            O => \N__10275\,
            I => \N__10261\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__10272\,
            I => \N__10247\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__10269\,
            I => \N__10240\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__10266\,
            I => \N__10229\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__10261\,
            I => \N__10226\
        );

    \I__2409\ : SRMux
    port map (
            O => \N__10260\,
            I => \N__10132\
        );

    \I__2408\ : SRMux
    port map (
            O => \N__10259\,
            I => \N__10132\
        );

    \I__2407\ : SRMux
    port map (
            O => \N__10258\,
            I => \N__10132\
        );

    \I__2406\ : SRMux
    port map (
            O => \N__10257\,
            I => \N__10132\
        );

    \I__2405\ : SRMux
    port map (
            O => \N__10256\,
            I => \N__10132\
        );

    \I__2404\ : SRMux
    port map (
            O => \N__10255\,
            I => \N__10132\
        );

    \I__2403\ : SRMux
    port map (
            O => \N__10254\,
            I => \N__10132\
        );

    \I__2402\ : SRMux
    port map (
            O => \N__10253\,
            I => \N__10132\
        );

    \I__2401\ : SRMux
    port map (
            O => \N__10252\,
            I => \N__10132\
        );

    \I__2400\ : SRMux
    port map (
            O => \N__10251\,
            I => \N__10132\
        );

    \I__2399\ : SRMux
    port map (
            O => \N__10250\,
            I => \N__10132\
        );

    \I__2398\ : Glb2LocalMux
    port map (
            O => \N__10247\,
            I => \N__10132\
        );

    \I__2397\ : SRMux
    port map (
            O => \N__10246\,
            I => \N__10132\
        );

    \I__2396\ : SRMux
    port map (
            O => \N__10245\,
            I => \N__10132\
        );

    \I__2395\ : SRMux
    port map (
            O => \N__10244\,
            I => \N__10132\
        );

    \I__2394\ : SRMux
    port map (
            O => \N__10243\,
            I => \N__10132\
        );

    \I__2393\ : Glb2LocalMux
    port map (
            O => \N__10240\,
            I => \N__10132\
        );

    \I__2392\ : SRMux
    port map (
            O => \N__10239\,
            I => \N__10132\
        );

    \I__2391\ : SRMux
    port map (
            O => \N__10238\,
            I => \N__10132\
        );

    \I__2390\ : SRMux
    port map (
            O => \N__10237\,
            I => \N__10132\
        );

    \I__2389\ : SRMux
    port map (
            O => \N__10236\,
            I => \N__10132\
        );

    \I__2388\ : SRMux
    port map (
            O => \N__10235\,
            I => \N__10132\
        );

    \I__2387\ : SRMux
    port map (
            O => \N__10234\,
            I => \N__10132\
        );

    \I__2386\ : SRMux
    port map (
            O => \N__10233\,
            I => \N__10132\
        );

    \I__2385\ : SRMux
    port map (
            O => \N__10232\,
            I => \N__10132\
        );

    \I__2384\ : Glb2LocalMux
    port map (
            O => \N__10229\,
            I => \N__10132\
        );

    \I__2383\ : Glb2LocalMux
    port map (
            O => \N__10226\,
            I => \N__10132\
        );

    \I__2382\ : SRMux
    port map (
            O => \N__10225\,
            I => \N__10132\
        );

    \I__2381\ : SRMux
    port map (
            O => \N__10224\,
            I => \N__10132\
        );

    \I__2380\ : SRMux
    port map (
            O => \N__10223\,
            I => \N__10132\
        );

    \I__2379\ : SRMux
    port map (
            O => \N__10222\,
            I => \N__10132\
        );

    \I__2378\ : SRMux
    port map (
            O => \N__10221\,
            I => \N__10132\
        );

    \I__2377\ : SRMux
    port map (
            O => \N__10220\,
            I => \N__10132\
        );

    \I__2376\ : SRMux
    port map (
            O => \N__10219\,
            I => \N__10132\
        );

    \I__2375\ : SRMux
    port map (
            O => \N__10218\,
            I => \N__10132\
        );

    \I__2374\ : SRMux
    port map (
            O => \N__10217\,
            I => \N__10132\
        );

    \I__2373\ : SRMux
    port map (
            O => \N__10216\,
            I => \N__10132\
        );

    \I__2372\ : SRMux
    port map (
            O => \N__10215\,
            I => \N__10132\
        );

    \I__2371\ : SRMux
    port map (
            O => \N__10214\,
            I => \N__10132\
        );

    \I__2370\ : SRMux
    port map (
            O => \N__10213\,
            I => \N__10132\
        );

    \I__2369\ : GlobalMux
    port map (
            O => \N__10132\,
            I => \N__10129\
        );

    \I__2368\ : gio2CtrlBuf
    port map (
            O => \N__10129\,
            I => \RESETn_c_i_g\
        );

    \I__2367\ : InMux
    port map (
            O => \N__10126\,
            I => \N__10123\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__10123\,
            I => \N__10120\
        );

    \I__2365\ : Sp12to4
    port map (
            O => \N__10120\,
            I => \N__10116\
        );

    \I__2364\ : InMux
    port map (
            O => \N__10119\,
            I => \N__10113\
        );

    \I__2363\ : Span12Mux_v
    port map (
            O => \N__10116\,
            I => \N__10110\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__10113\,
            I => \N__10107\
        );

    \I__2361\ : Span12Mux_h
    port map (
            O => \N__10110\,
            I => \N__10103\
        );

    \I__2360\ : Span4Mux_v
    port map (
            O => \N__10107\,
            I => \N__10100\
        );

    \I__2359\ : InMux
    port map (
            O => \N__10106\,
            I => \N__10097\
        );

    \I__2358\ : Odrv12
    port map (
            O => \N__10103\,
            I => \REG_CYCLEm\
        );

    \I__2357\ : Odrv4
    port map (
            O => \N__10100\,
            I => \REG_CYCLEm\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__10097\,
            I => \REG_CYCLEm\
        );

    \I__2355\ : InMux
    port map (
            O => \N__10090\,
            I => \N__10087\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__10087\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__2353\ : InMux
    port map (
            O => \N__10084\,
            I => \N__10081\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__10081\,
            I => \N__10077\
        );

    \I__2351\ : InMux
    port map (
            O => \N__10080\,
            I => \N__10074\
        );

    \I__2350\ : Span4Mux_h
    port map (
            O => \N__10077\,
            I => \N__10069\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__10074\,
            I => \N__10069\
        );

    \I__2348\ : Span4Mux_v
    port map (
            O => \N__10069\,
            I => \N__10064\
        );

    \I__2347\ : InMux
    port map (
            O => \N__10068\,
            I => \N__10061\
        );

    \I__2346\ : InMux
    port map (
            O => \N__10067\,
            I => \N__10058\
        );

    \I__2345\ : Span4Mux_v
    port map (
            O => \N__10064\,
            I => \N__10055\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__10061\,
            I => \N__10050\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__10058\,
            I => \N__10050\
        );

    \I__2342\ : Sp12to4
    port map (
            O => \N__10055\,
            I => \N__10045\
        );

    \I__2341\ : Span12Mux_v
    port map (
            O => \N__10050\,
            I => \N__10045\
        );

    \I__2340\ : Span12Mux_h
    port map (
            O => \N__10045\,
            I => \N__10042\
        );

    \I__2339\ : Odrv12
    port map (
            O => \N__10042\,
            I => \DRA_c_5\
        );

    \I__2338\ : InMux
    port map (
            O => \N__10039\,
            I => \N__10033\
        );

    \I__2337\ : InMux
    port map (
            O => \N__10038\,
            I => \N__10033\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__10033\,
            I => \N__10030\
        );

    \I__2335\ : Span4Mux_v
    port map (
            O => \N__10030\,
            I => \N__10027\
        );

    \I__2334\ : Odrv4
    port map (
            O => \N__10027\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__2333\ : CascadeMux
    port map (
            O => \N__10024\,
            I => \N__10021\
        );

    \I__2332\ : InMux
    port map (
            O => \N__10021\,
            I => \N__10013\
        );

    \I__2331\ : InMux
    port map (
            O => \N__10020\,
            I => \N__10013\
        );

    \I__2330\ : InMux
    port map (
            O => \N__10019\,
            I => \N__10010\
        );

    \I__2329\ : InMux
    port map (
            O => \N__10018\,
            I => \N__10007\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__10013\,
            I => \N__10002\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__10010\,
            I => \N__10002\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__10007\,
            I => \N__9999\
        );

    \I__2325\ : Span4Mux_v
    port map (
            O => \N__10002\,
            I => \N__9996\
        );

    \I__2324\ : Sp12to4
    port map (
            O => \N__9999\,
            I => \N__9993\
        );

    \I__2323\ : Sp12to4
    port map (
            O => \N__9996\,
            I => \N__9990\
        );

    \I__2322\ : Span12Mux_v
    port map (
            O => \N__9993\,
            I => \N__9987\
        );

    \I__2321\ : Span12Mux_h
    port map (
            O => \N__9990\,
            I => \N__9984\
        );

    \I__2320\ : Span12Mux_h
    port map (
            O => \N__9987\,
            I => \N__9979\
        );

    \I__2319\ : Span12Mux_v
    port map (
            O => \N__9984\,
            I => \N__9979\
        );

    \I__2318\ : Odrv12
    port map (
            O => \N__9979\,
            I => \DRA_c_2\
        );

    \I__2317\ : InMux
    port map (
            O => \N__9976\,
            I => \N__9973\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__9973\,
            I => \N__9970\
        );

    \I__2315\ : Odrv4
    port map (
            O => \N__9970\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__2314\ : InMux
    port map (
            O => \N__9967\,
            I => \N__9964\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__9964\,
            I => \N__9961\
        );

    \I__2312\ : Span4Mux_h
    port map (
            O => \N__9961\,
            I => \N__9958\
        );

    \I__2311\ : Odrv4
    port map (
            O => \N__9958\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__2310\ : InMux
    port map (
            O => \N__9955\,
            I => \N__9950\
        );

    \I__2309\ : InMux
    port map (
            O => \N__9954\,
            I => \N__9947\
        );

    \I__2308\ : InMux
    port map (
            O => \N__9953\,
            I => \N__9943\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__9950\,
            I => \N__9938\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__9947\,
            I => \N__9938\
        );

    \I__2305\ : InMux
    port map (
            O => \N__9946\,
            I => \N__9935\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__9943\,
            I => \N__9932\
        );

    \I__2303\ : Span4Mux_v
    port map (
            O => \N__9938\,
            I => \N__9925\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__9935\,
            I => \N__9925\
        );

    \I__2301\ : Span4Mux_v
    port map (
            O => \N__9932\,
            I => \N__9925\
        );

    \I__2300\ : Sp12to4
    port map (
            O => \N__9925\,
            I => \N__9922\
        );

    \I__2299\ : Span12Mux_h
    port map (
            O => \N__9922\,
            I => \N__9919\
        );

    \I__2298\ : Span12Mux_v
    port map (
            O => \N__9919\,
            I => \N__9916\
        );

    \I__2297\ : Odrv12
    port map (
            O => \N__9916\,
            I => \DRA_c_1\
        );

    \I__2296\ : InMux
    port map (
            O => \N__9913\,
            I => \N__9910\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__9910\,
            I => \N__9906\
        );

    \I__2294\ : InMux
    port map (
            O => \N__9909\,
            I => \N__9903\
        );

    \I__2293\ : Sp12to4
    port map (
            O => \N__9906\,
            I => \N__9900\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__9903\,
            I => \N__9897\
        );

    \I__2291\ : Span12Mux_v
    port map (
            O => \N__9900\,
            I => \N__9894\
        );

    \I__2290\ : Span12Mux_h
    port map (
            O => \N__9897\,
            I => \N__9891\
        );

    \I__2289\ : Span12Mux_h
    port map (
            O => \N__9894\,
            I => \N__9888\
        );

    \I__2288\ : Span12Mux_v
    port map (
            O => \N__9891\,
            I => \N__9885\
        );

    \I__2287\ : Odrv12
    port map (
            O => \N__9888\,
            I => \DRA_c_0\
        );

    \I__2286\ : Odrv12
    port map (
            O => \N__9885\,
            I => \DRA_c_0\
        );

    \I__2285\ : InMux
    port map (
            O => \N__9880\,
            I => \N__9877\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__9877\,
            I => \N__9874\
        );

    \I__2283\ : Span4Mux_h
    port map (
            O => \N__9874\,
            I => \N__9871\
        );

    \I__2282\ : Odrv4
    port map (
            O => \N__9871\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2281\ : IoInMux
    port map (
            O => \N__9868\,
            I => \N__9865\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__9865\,
            I => \N__9862\
        );

    \I__2279\ : Sp12to4
    port map (
            O => \N__9862\,
            I => \N__9859\
        );

    \I__2278\ : Span12Mux_h
    port map (
            O => \N__9859\,
            I => \N__9856\
        );

    \I__2277\ : Span12Mux_v
    port map (
            O => \N__9856\,
            I => \N__9853\
        );

    \I__2276\ : Odrv12
    port map (
            O => \N__9853\,
            I => \N_57_i\
        );

    \I__2275\ : CascadeMux
    port map (
            O => \N__9850\,
            I => \N__9846\
        );

    \I__2274\ : IoInMux
    port map (
            O => \N__9849\,
            I => \N__9842\
        );

    \I__2273\ : InMux
    port map (
            O => \N__9846\,
            I => \N__9839\
        );

    \I__2272\ : InMux
    port map (
            O => \N__9845\,
            I => \N__9836\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__9842\,
            I => \N__9831\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__9839\,
            I => \N__9826\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__9836\,
            I => \N__9826\
        );

    \I__2268\ : InMux
    port map (
            O => \N__9835\,
            I => \N__9823\
        );

    \I__2267\ : InMux
    port map (
            O => \N__9834\,
            I => \N__9820\
        );

    \I__2266\ : Span12Mux_s2_v
    port map (
            O => \N__9831\,
            I => \N__9817\
        );

    \I__2265\ : Span4Mux_v
    port map (
            O => \N__9826\,
            I => \N__9814\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__9823\,
            I => \N__9809\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__9820\,
            I => \N__9809\
        );

    \I__2262\ : Span12Mux_v
    port map (
            O => \N__9817\,
            I => \N__9805\
        );

    \I__2261\ : Span4Mux_h
    port map (
            O => \N__9814\,
            I => \N__9802\
        );

    \I__2260\ : Span4Mux_v
    port map (
            O => \N__9809\,
            I => \N__9799\
        );

    \I__2259\ : InMux
    port map (
            O => \N__9808\,
            I => \N__9796\
        );

    \I__2258\ : Odrv12
    port map (
            O => \N__9805\,
            I => \DBENn_c\
        );

    \I__2257\ : Odrv4
    port map (
            O => \N__9802\,
            I => \DBENn_c\
        );

    \I__2256\ : Odrv4
    port map (
            O => \N__9799\,
            I => \DBENn_c\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__9796\,
            I => \DBENn_c\
        );

    \I__2254\ : CascadeMux
    port map (
            O => \N__9787\,
            I => \N__9784\
        );

    \I__2253\ : InMux
    port map (
            O => \N__9784\,
            I => \N__9778\
        );

    \I__2252\ : InMux
    port map (
            O => \N__9783\,
            I => \N__9775\
        );

    \I__2251\ : InMux
    port map (
            O => \N__9782\,
            I => \N__9771\
        );

    \I__2250\ : InMux
    port map (
            O => \N__9781\,
            I => \N__9767\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__9778\,
            I => \N__9764\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__9775\,
            I => \N__9761\
        );

    \I__2247\ : InMux
    port map (
            O => \N__9774\,
            I => \N__9758\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__9771\,
            I => \N__9754\
        );

    \I__2245\ : InMux
    port map (
            O => \N__9770\,
            I => \N__9751\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__9767\,
            I => \N__9748\
        );

    \I__2243\ : Span4Mux_h
    port map (
            O => \N__9764\,
            I => \N__9743\
        );

    \I__2242\ : Span4Mux_v
    port map (
            O => \N__9761\,
            I => \N__9743\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__9758\,
            I => \N__9740\
        );

    \I__2240\ : InMux
    port map (
            O => \N__9757\,
            I => \N__9735\
        );

    \I__2239\ : Span4Mux_v
    port map (
            O => \N__9754\,
            I => \N__9732\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__9751\,
            I => \N__9729\
        );

    \I__2237\ : Span4Mux_v
    port map (
            O => \N__9748\,
            I => \N__9726\
        );

    \I__2236\ : Span4Mux_v
    port map (
            O => \N__9743\,
            I => \N__9721\
        );

    \I__2235\ : Span4Mux_v
    port map (
            O => \N__9740\,
            I => \N__9721\
        );

    \I__2234\ : InMux
    port map (
            O => \N__9739\,
            I => \N__9718\
        );

    \I__2233\ : InMux
    port map (
            O => \N__9738\,
            I => \N__9715\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__9735\,
            I => \N__9712\
        );

    \I__2231\ : Span4Mux_h
    port map (
            O => \N__9732\,
            I => \N__9707\
        );

    \I__2230\ : Span4Mux_h
    port map (
            O => \N__9729\,
            I => \N__9707\
        );

    \I__2229\ : Odrv4
    port map (
            O => \N__9726\,
            I => \DMA_CYCLEm\
        );

    \I__2228\ : Odrv4
    port map (
            O => \N__9721\,
            I => \DMA_CYCLEm\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__9718\,
            I => \DMA_CYCLEm\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__9715\,
            I => \DMA_CYCLEm\
        );

    \I__2225\ : Odrv12
    port map (
            O => \N__9712\,
            I => \DMA_CYCLEm\
        );

    \I__2224\ : Odrv4
    port map (
            O => \N__9707\,
            I => \DMA_CYCLEm\
        );

    \I__2223\ : IoInMux
    port map (
            O => \N__9694\,
            I => \N__9691\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__9691\,
            I => \N__9688\
        );

    \I__2221\ : Span4Mux_s2_h
    port map (
            O => \N__9688\,
            I => \N__9685\
        );

    \I__2220\ : Span4Mux_v
    port map (
            O => \N__9685\,
            I => \N__9682\
        );

    \I__2219\ : Span4Mux_v
    port map (
            O => \N__9682\,
            I => \N__9679\
        );

    \I__2218\ : Sp12to4
    port map (
            O => \N__9679\,
            I => \N__9676\
        );

    \I__2217\ : Odrv12
    port map (
            O => \N__9676\,
            I => \N_59_i\
        );

    \I__2216\ : InMux
    port map (
            O => \N__9673\,
            I => \N__9670\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__9670\,
            I => \U712_BYTE_ENABLE.N_557\
        );

    \I__2214\ : CascadeMux
    port map (
            O => \N__9667\,
            I => \N__9660\
        );

    \I__2213\ : InMux
    port map (
            O => \N__9666\,
            I => \N__9655\
        );

    \I__2212\ : CascadeMux
    port map (
            O => \N__9665\,
            I => \N__9652\
        );

    \I__2211\ : CascadeMux
    port map (
            O => \N__9664\,
            I => \N__9649\
        );

    \I__2210\ : CascadeMux
    port map (
            O => \N__9663\,
            I => \N__9645\
        );

    \I__2209\ : InMux
    port map (
            O => \N__9660\,
            I => \N__9640\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__9659\,
            I => \N__9637\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__9658\,
            I => \N__9630\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__9655\,
            I => \N__9625\
        );

    \I__2205\ : InMux
    port map (
            O => \N__9652\,
            I => \N__9622\
        );

    \I__2204\ : InMux
    port map (
            O => \N__9649\,
            I => \N__9617\
        );

    \I__2203\ : InMux
    port map (
            O => \N__9648\,
            I => \N__9613\
        );

    \I__2202\ : InMux
    port map (
            O => \N__9645\,
            I => \N__9606\
        );

    \I__2201\ : InMux
    port map (
            O => \N__9644\,
            I => \N__9606\
        );

    \I__2200\ : InMux
    port map (
            O => \N__9643\,
            I => \N__9606\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__9640\,
            I => \N__9603\
        );

    \I__2198\ : InMux
    port map (
            O => \N__9637\,
            I => \N__9600\
        );

    \I__2197\ : InMux
    port map (
            O => \N__9636\,
            I => \N__9597\
        );

    \I__2196\ : InMux
    port map (
            O => \N__9635\,
            I => \N__9592\
        );

    \I__2195\ : InMux
    port map (
            O => \N__9634\,
            I => \N__9592\
        );

    \I__2194\ : InMux
    port map (
            O => \N__9633\,
            I => \N__9589\
        );

    \I__2193\ : InMux
    port map (
            O => \N__9630\,
            I => \N__9586\
        );

    \I__2192\ : InMux
    port map (
            O => \N__9629\,
            I => \N__9580\
        );

    \I__2191\ : InMux
    port map (
            O => \N__9628\,
            I => \N__9580\
        );

    \I__2190\ : Span4Mux_v
    port map (
            O => \N__9625\,
            I => \N__9572\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__9622\,
            I => \N__9572\
        );

    \I__2188\ : InMux
    port map (
            O => \N__9621\,
            I => \N__9567\
        );

    \I__2187\ : InMux
    port map (
            O => \N__9620\,
            I => \N__9567\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__9617\,
            I => \N__9564\
        );

    \I__2185\ : InMux
    port map (
            O => \N__9616\,
            I => \N__9561\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__9613\,
            I => \N__9556\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__9606\,
            I => \N__9556\
        );

    \I__2182\ : Span4Mux_v
    port map (
            O => \N__9603\,
            I => \N__9547\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__9600\,
            I => \N__9547\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__9597\,
            I => \N__9547\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__9592\,
            I => \N__9547\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__9589\,
            I => \N__9544\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__9586\,
            I => \N__9541\
        );

    \I__2176\ : InMux
    port map (
            O => \N__9585\,
            I => \N__9538\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__9580\,
            I => \N__9535\
        );

    \I__2174\ : InMux
    port map (
            O => \N__9579\,
            I => \N__9532\
        );

    \I__2173\ : InMux
    port map (
            O => \N__9578\,
            I => \N__9527\
        );

    \I__2172\ : InMux
    port map (
            O => \N__9577\,
            I => \N__9527\
        );

    \I__2171\ : Span4Mux_v
    port map (
            O => \N__9572\,
            I => \N__9520\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__9567\,
            I => \N__9520\
        );

    \I__2169\ : Span4Mux_v
    port map (
            O => \N__9564\,
            I => \N__9520\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__9561\,
            I => \N__9513\
        );

    \I__2167\ : Span4Mux_h
    port map (
            O => \N__9556\,
            I => \N__9513\
        );

    \I__2166\ : Span4Mux_v
    port map (
            O => \N__9547\,
            I => \N__9513\
        );

    \I__2165\ : Span4Mux_v
    port map (
            O => \N__9544\,
            I => \N__9506\
        );

    \I__2164\ : Span4Mux_h
    port map (
            O => \N__9541\,
            I => \N__9506\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__9538\,
            I => \N__9506\
        );

    \I__2162\ : Span12Mux_h
    port map (
            O => \N__9535\,
            I => \N__9501\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__9532\,
            I => \N__9501\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__9527\,
            I => \CPU_CYCLEm\
        );

    \I__2159\ : Odrv4
    port map (
            O => \N__9520\,
            I => \CPU_CYCLEm\
        );

    \I__2158\ : Odrv4
    port map (
            O => \N__9513\,
            I => \CPU_CYCLEm\
        );

    \I__2157\ : Odrv4
    port map (
            O => \N__9506\,
            I => \CPU_CYCLEm\
        );

    \I__2156\ : Odrv12
    port map (
            O => \N__9501\,
            I => \CPU_CYCLEm\
        );

    \I__2155\ : InMux
    port map (
            O => \N__9490\,
            I => \N__9487\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__9487\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2153\ : InMux
    port map (
            O => \N__9484\,
            I => \N__9481\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__9481\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__2151\ : InMux
    port map (
            O => \N__9478\,
            I => \N__9475\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__9475\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2149\ : InMux
    port map (
            O => \N__9472\,
            I => \N__9469\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__9469\,
            I => \N__9466\
        );

    \I__2147\ : Span4Mux_h
    port map (
            O => \N__9466\,
            I => \N__9463\
        );

    \I__2146\ : Odrv4
    port map (
            O => \N__9463\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__2145\ : InMux
    port map (
            O => \N__9460\,
            I => \N__9457\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__9457\,
            I => \N__9452\
        );

    \I__2143\ : InMux
    port map (
            O => \N__9456\,
            I => \N__9449\
        );

    \I__2142\ : InMux
    port map (
            O => \N__9455\,
            I => \N__9445\
        );

    \I__2141\ : Span4Mux_h
    port map (
            O => \N__9452\,
            I => \N__9440\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__9449\,
            I => \N__9440\
        );

    \I__2139\ : InMux
    port map (
            O => \N__9448\,
            I => \N__9437\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__9445\,
            I => \N__9430\
        );

    \I__2137\ : Sp12to4
    port map (
            O => \N__9440\,
            I => \N__9430\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9437\,
            I => \N__9430\
        );

    \I__2135\ : Span12Mux_v
    port map (
            O => \N__9430\,
            I => \N__9427\
        );

    \I__2134\ : Span12Mux_h
    port map (
            O => \N__9427\,
            I => \N__9424\
        );

    \I__2133\ : Odrv12
    port map (
            O => \N__9424\,
            I => \DRA_c_3\
        );

    \I__2132\ : InMux
    port map (
            O => \N__9421\,
            I => \N__9418\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__9418\,
            I => \N__9415\
        );

    \I__2130\ : Span4Mux_h
    port map (
            O => \N__9415\,
            I => \N__9412\
        );

    \I__2129\ : Odrv4
    port map (
            O => \N__9412\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__2128\ : InMux
    port map (
            O => \N__9409\,
            I => \N__9402\
        );

    \I__2127\ : InMux
    port map (
            O => \N__9408\,
            I => \N__9402\
        );

    \I__2126\ : InMux
    port map (
            O => \N__9407\,
            I => \N__9399\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__9402\,
            I => \N__9395\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__9399\,
            I => \N__9392\
        );

    \I__2123\ : InMux
    port map (
            O => \N__9398\,
            I => \N__9389\
        );

    \I__2122\ : Span4Mux_v
    port map (
            O => \N__9395\,
            I => \N__9382\
        );

    \I__2121\ : Span4Mux_h
    port map (
            O => \N__9392\,
            I => \N__9382\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__9389\,
            I => \N__9382\
        );

    \I__2119\ : Span4Mux_v
    port map (
            O => \N__9382\,
            I => \N__9379\
        );

    \I__2118\ : Span4Mux_v
    port map (
            O => \N__9379\,
            I => \N__9376\
        );

    \I__2117\ : Sp12to4
    port map (
            O => \N__9376\,
            I => \N__9373\
        );

    \I__2116\ : Span12Mux_h
    port map (
            O => \N__9373\,
            I => \N__9370\
        );

    \I__2115\ : Odrv12
    port map (
            O => \N__9370\,
            I => \DRA_c_4\
        );

    \I__2114\ : InMux
    port map (
            O => \N__9367\,
            I => \N__9364\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__9364\,
            I => \N__9361\
        );

    \I__2112\ : Odrv4
    port map (
            O => \N__9361\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__2111\ : IoInMux
    port map (
            O => \N__9358\,
            I => \N__9355\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__9355\,
            I => \N__9352\
        );

    \I__2109\ : Span4Mux_s2_v
    port map (
            O => \N__9352\,
            I => \N__9349\
        );

    \I__2108\ : Span4Mux_v
    port map (
            O => \N__9349\,
            I => \N__9346\
        );

    \I__2107\ : Sp12to4
    port map (
            O => \N__9346\,
            I => \N__9343\
        );

    \I__2106\ : Odrv12
    port map (
            O => \N__9343\,
            I => \un1_UDSn_i_0_0\
        );

    \I__2105\ : InMux
    port map (
            O => \N__9340\,
            I => \N__9334\
        );

    \I__2104\ : InMux
    port map (
            O => \N__9339\,
            I => \N__9334\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__9334\,
            I => \N__9331\
        );

    \I__2102\ : Span4Mux_v
    port map (
            O => \N__9331\,
            I => \N__9328\
        );

    \I__2101\ : Span4Mux_h
    port map (
            O => \N__9328\,
            I => \N__9325\
        );

    \I__2100\ : Span4Mux_v
    port map (
            O => \N__9325\,
            I => \N__9321\
        );

    \I__2099\ : InMux
    port map (
            O => \N__9324\,
            I => \N__9318\
        );

    \I__2098\ : Odrv4
    port map (
            O => \N__9321\,
            I => \DS_ENm\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__9318\,
            I => \DS_ENm\
        );

    \I__2096\ : IoInMux
    port map (
            O => \N__9313\,
            I => \N__9310\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__9310\,
            I => \N__9307\
        );

    \I__2094\ : Span12Mux_s6_v
    port map (
            O => \N__9307\,
            I => \N__9304\
        );

    \I__2093\ : Odrv12
    port map (
            O => \N__9304\,
            I => \un1_LDSn_i_0_0\
        );

    \I__2092\ : CascadeMux
    port map (
            O => \N__9301\,
            I => \N__9298\
        );

    \I__2091\ : InMux
    port map (
            O => \N__9298\,
            I => \N__9295\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__9295\,
            I => \N__9292\
        );

    \I__2089\ : Odrv12
    port map (
            O => \N__9292\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__2088\ : InMux
    port map (
            O => \N__9289\,
            I => \N__9286\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__9286\,
            I => \N__9282\
        );

    \I__2086\ : InMux
    port map (
            O => \N__9285\,
            I => \N__9279\
        );

    \I__2085\ : Odrv12
    port map (
            O => \N__9282\,
            I => \DBRn_c_i\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__9279\,
            I => \DBRn_c_i\
        );

    \I__2083\ : InMux
    port map (
            O => \N__9274\,
            I => \N__9271\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__9271\,
            I => \N__9267\
        );

    \I__2081\ : InMux
    port map (
            O => \N__9270\,
            I => \N__9264\
        );

    \I__2080\ : Span4Mux_h
    port map (
            O => \N__9267\,
            I => \N__9261\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__9264\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__9261\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__2077\ : IoInMux
    port map (
            O => \N__9256\,
            I => \N__9253\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__9253\,
            I => \N__9250\
        );

    \I__2075\ : IoSpan4Mux
    port map (
            O => \N__9250\,
            I => \N__9247\
        );

    \I__2074\ : Span4Mux_s1_h
    port map (
            O => \N__9247\,
            I => \N__9244\
        );

    \I__2073\ : Sp12to4
    port map (
            O => \N__9244\,
            I => \N__9241\
        );

    \I__2072\ : Span12Mux_h
    port map (
            O => \N__9241\,
            I => \N__9238\
        );

    \I__2071\ : Span12Mux_v
    port map (
            O => \N__9238\,
            I => \N__9235\
        );

    \I__2070\ : Odrv12
    port map (
            O => \N__9235\,
            I => \N_58_i\
        );

    \I__2069\ : CascadeMux
    port map (
            O => \N__9232\,
            I => \N__9229\
        );

    \I__2068\ : InMux
    port map (
            O => \N__9229\,
            I => \N__9225\
        );

    \I__2067\ : InMux
    port map (
            O => \N__9228\,
            I => \N__9222\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__9225\,
            I => \N__9219\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__9222\,
            I => \N__9216\
        );

    \I__2064\ : Odrv4
    port map (
            O => \N__9219\,
            I => \U712_BYTE_ENABLE.N_410\
        );

    \I__2063\ : Odrv4
    port map (
            O => \N__9216\,
            I => \U712_BYTE_ENABLE.N_410\
        );

    \I__2062\ : CascadeMux
    port map (
            O => \N__9211\,
            I => \N__9208\
        );

    \I__2061\ : InMux
    port map (
            O => \N__9208\,
            I => \N__9205\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__9205\,
            I => \U712_BYTE_ENABLE.N_559\
        );

    \I__2059\ : IoInMux
    port map (
            O => \N__9202\,
            I => \N__9199\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__9199\,
            I => \N__9196\
        );

    \I__2057\ : IoSpan4Mux
    port map (
            O => \N__9196\,
            I => \N__9193\
        );

    \I__2056\ : Span4Mux_s3_v
    port map (
            O => \N__9193\,
            I => \N__9190\
        );

    \I__2055\ : Odrv4
    port map (
            O => \N__9190\,
            I => \N_129_i\
        );

    \I__2054\ : IoInMux
    port map (
            O => \N__9187\,
            I => \N__9184\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__9184\,
            I => \N__9181\
        );

    \I__2052\ : IoSpan4Mux
    port map (
            O => \N__9181\,
            I => \N__9178\
        );

    \I__2051\ : Sp12to4
    port map (
            O => \N__9178\,
            I => \N__9175\
        );

    \I__2050\ : Span12Mux_s7_v
    port map (
            O => \N__9175\,
            I => \N__9172\
        );

    \I__2049\ : Odrv12
    port map (
            O => \N__9172\,
            I => \CASn_c\
        );

    \I__2048\ : InMux
    port map (
            O => \N__9169\,
            I => \N__9165\
        );

    \I__2047\ : InMux
    port map (
            O => \N__9168\,
            I => \N__9162\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__9165\,
            I => \N__9155\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__9162\,
            I => \N__9155\
        );

    \I__2044\ : CascadeMux
    port map (
            O => \N__9161\,
            I => \N__9152\
        );

    \I__2043\ : InMux
    port map (
            O => \N__9160\,
            I => \N__9149\
        );

    \I__2042\ : Span4Mux_h
    port map (
            O => \N__9155\,
            I => \N__9144\
        );

    \I__2041\ : InMux
    port map (
            O => \N__9152\,
            I => \N__9141\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__9149\,
            I => \N__9138\
        );

    \I__2039\ : InMux
    port map (
            O => \N__9148\,
            I => \N__9133\
        );

    \I__2038\ : InMux
    port map (
            O => \N__9147\,
            I => \N__9133\
        );

    \I__2037\ : Span4Mux_h
    port map (
            O => \N__9144\,
            I => \N__9130\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__9141\,
            I => \N__9123\
        );

    \I__2035\ : Span4Mux_v
    port map (
            O => \N__9138\,
            I => \N__9123\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__9133\,
            I => \N__9123\
        );

    \I__2033\ : Odrv4
    port map (
            O => \N__9130\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2032\ : Odrv4
    port map (
            O => \N__9123\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2031\ : IoInMux
    port map (
            O => \N__9118\,
            I => \N__9115\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__9115\,
            I => \N__9112\
        );

    \I__2029\ : IoSpan4Mux
    port map (
            O => \N__9112\,
            I => \N__9109\
        );

    \I__2028\ : Sp12to4
    port map (
            O => \N__9109\,
            I => \N__9106\
        );

    \I__2027\ : Span12Mux_s9_v
    port map (
            O => \N__9106\,
            I => \N__9103\
        );

    \I__2026\ : Odrv12
    port map (
            O => \N__9103\,
            I => \RASn_c\
        );

    \I__2025\ : InMux
    port map (
            O => \N__9100\,
            I => \N__9097\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__9097\,
            I => \N__9094\
        );

    \I__2023\ : Span12Mux_h
    port map (
            O => \N__9094\,
            I => \N__9091\
        );

    \I__2022\ : Odrv12
    port map (
            O => \N__9091\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\
        );

    \I__2021\ : InMux
    port map (
            O => \N__9088\,
            I => \N__9083\
        );

    \I__2020\ : CascadeMux
    port map (
            O => \N__9087\,
            I => \N__9080\
        );

    \I__2019\ : CascadeMux
    port map (
            O => \N__9086\,
            I => \N__9077\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__9083\,
            I => \N__9065\
        );

    \I__2017\ : InMux
    port map (
            O => \N__9080\,
            I => \N__9062\
        );

    \I__2016\ : InMux
    port map (
            O => \N__9077\,
            I => \N__9059\
        );

    \I__2015\ : InMux
    port map (
            O => \N__9076\,
            I => \N__9052\
        );

    \I__2014\ : InMux
    port map (
            O => \N__9075\,
            I => \N__9052\
        );

    \I__2013\ : InMux
    port map (
            O => \N__9074\,
            I => \N__9052\
        );

    \I__2012\ : InMux
    port map (
            O => \N__9073\,
            I => \N__9047\
        );

    \I__2011\ : InMux
    port map (
            O => \N__9072\,
            I => \N__9044\
        );

    \I__2010\ : InMux
    port map (
            O => \N__9071\,
            I => \N__9039\
        );

    \I__2009\ : InMux
    port map (
            O => \N__9070\,
            I => \N__9039\
        );

    \I__2008\ : InMux
    port map (
            O => \N__9069\,
            I => \N__9036\
        );

    \I__2007\ : InMux
    port map (
            O => \N__9068\,
            I => \N__9032\
        );

    \I__2006\ : Span4Mux_v
    port map (
            O => \N__9065\,
            I => \N__9023\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__9062\,
            I => \N__9023\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__9059\,
            I => \N__9023\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__9052\,
            I => \N__9023\
        );

    \I__2002\ : InMux
    port map (
            O => \N__9051\,
            I => \N__9016\
        );

    \I__2001\ : InMux
    port map (
            O => \N__9050\,
            I => \N__9016\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__9047\,
            I => \N__9011\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__9044\,
            I => \N__9011\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__9039\,
            I => \N__9006\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__9036\,
            I => \N__9006\
        );

    \I__1996\ : InMux
    port map (
            O => \N__9035\,
            I => \N__8998\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__9032\,
            I => \N__8991\
        );

    \I__1994\ : Span4Mux_h
    port map (
            O => \N__9023\,
            I => \N__8991\
        );

    \I__1993\ : InMux
    port map (
            O => \N__9022\,
            I => \N__8988\
        );

    \I__1992\ : InMux
    port map (
            O => \N__9021\,
            I => \N__8985\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__9016\,
            I => \N__8982\
        );

    \I__1990\ : Span4Mux_v
    port map (
            O => \N__9011\,
            I => \N__8977\
        );

    \I__1989\ : Span4Mux_v
    port map (
            O => \N__9006\,
            I => \N__8977\
        );

    \I__1988\ : InMux
    port map (
            O => \N__9005\,
            I => \N__8970\
        );

    \I__1987\ : InMux
    port map (
            O => \N__9004\,
            I => \N__8970\
        );

    \I__1986\ : InMux
    port map (
            O => \N__9003\,
            I => \N__8970\
        );

    \I__1985\ : InMux
    port map (
            O => \N__9002\,
            I => \N__8967\
        );

    \I__1984\ : InMux
    port map (
            O => \N__9001\,
            I => \N__8964\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__8998\,
            I => \N__8961\
        );

    \I__1982\ : InMux
    port map (
            O => \N__8997\,
            I => \N__8956\
        );

    \I__1981\ : InMux
    port map (
            O => \N__8996\,
            I => \N__8956\
        );

    \I__1980\ : Span4Mux_h
    port map (
            O => \N__8991\,
            I => \N__8951\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__8988\,
            I => \N__8951\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__8985\,
            I => \N__8942\
        );

    \I__1977\ : Span12Mux_s11_v
    port map (
            O => \N__8982\,
            I => \N__8942\
        );

    \I__1976\ : Sp12to4
    port map (
            O => \N__8977\,
            I => \N__8942\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__8970\,
            I => \N__8942\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__8967\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__8964\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1972\ : Odrv4
    port map (
            O => \N__8961\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__8956\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1970\ : Odrv4
    port map (
            O => \N__8951\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1969\ : Odrv12
    port map (
            O => \N__8942\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1968\ : InMux
    port map (
            O => \N__8929\,
            I => \N__8923\
        );

    \I__1967\ : InMux
    port map (
            O => \N__8928\,
            I => \N__8916\
        );

    \I__1966\ : InMux
    port map (
            O => \N__8927\,
            I => \N__8916\
        );

    \I__1965\ : InMux
    port map (
            O => \N__8926\,
            I => \N__8913\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__8923\,
            I => \N__8910\
        );

    \I__1963\ : InMux
    port map (
            O => \N__8922\,
            I => \N__8905\
        );

    \I__1962\ : InMux
    port map (
            O => \N__8921\,
            I => \N__8905\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__8916\,
            I => \N__8902\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__8913\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__1959\ : Odrv4
    port map (
            O => \N__8910\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__8905\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__8902\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__1956\ : CascadeMux
    port map (
            O => \N__8893\,
            I => \N__8885\
        );

    \I__1955\ : CascadeMux
    port map (
            O => \N__8892\,
            I => \N__8882\
        );

    \I__1954\ : CascadeMux
    port map (
            O => \N__8891\,
            I => \N__8879\
        );

    \I__1953\ : CascadeMux
    port map (
            O => \N__8890\,
            I => \N__8876\
        );

    \I__1952\ : InMux
    port map (
            O => \N__8889\,
            I => \N__8871\
        );

    \I__1951\ : InMux
    port map (
            O => \N__8888\,
            I => \N__8868\
        );

    \I__1950\ : InMux
    port map (
            O => \N__8885\,
            I => \N__8864\
        );

    \I__1949\ : InMux
    port map (
            O => \N__8882\,
            I => \N__8861\
        );

    \I__1948\ : InMux
    port map (
            O => \N__8879\,
            I => \N__8856\
        );

    \I__1947\ : InMux
    port map (
            O => \N__8876\,
            I => \N__8856\
        );

    \I__1946\ : InMux
    port map (
            O => \N__8875\,
            I => \N__8851\
        );

    \I__1945\ : InMux
    port map (
            O => \N__8874\,
            I => \N__8851\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__8871\,
            I => \N__8848\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__8868\,
            I => \N__8845\
        );

    \I__1942\ : InMux
    port map (
            O => \N__8867\,
            I => \N__8842\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__8864\,
            I => \U712_CHIP_RAM.N_412\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__8861\,
            I => \U712_CHIP_RAM.N_412\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__8856\,
            I => \U712_CHIP_RAM.N_412\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__8851\,
            I => \U712_CHIP_RAM.N_412\
        );

    \I__1937\ : Odrv4
    port map (
            O => \N__8848\,
            I => \U712_CHIP_RAM.N_412\
        );

    \I__1936\ : Odrv4
    port map (
            O => \N__8845\,
            I => \U712_CHIP_RAM.N_412\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__8842\,
            I => \U712_CHIP_RAM.N_412\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__8827\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4_cascade_\
        );

    \I__1933\ : IoInMux
    port map (
            O => \N__8824\,
            I => \N__8821\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__8821\,
            I => \N__8818\
        );

    \I__1931\ : IoSpan4Mux
    port map (
            O => \N__8818\,
            I => \N__8815\
        );

    \I__1930\ : Span4Mux_s3_h
    port map (
            O => \N__8815\,
            I => \N__8812\
        );

    \I__1929\ : Sp12to4
    port map (
            O => \N__8812\,
            I => \N__8809\
        );

    \I__1928\ : Span12Mux_h
    port map (
            O => \N__8809\,
            I => \N__8806\
        );

    \I__1927\ : Odrv12
    port map (
            O => \N__8806\,
            I => \CMA_c_4\
        );

    \I__1926\ : InMux
    port map (
            O => \N__8803\,
            I => \N__8800\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__8800\,
            I => \N__8770\
        );

    \I__1924\ : ClkMux
    port map (
            O => \N__8799\,
            I => \N__8680\
        );

    \I__1923\ : ClkMux
    port map (
            O => \N__8798\,
            I => \N__8680\
        );

    \I__1922\ : ClkMux
    port map (
            O => \N__8797\,
            I => \N__8680\
        );

    \I__1921\ : ClkMux
    port map (
            O => \N__8796\,
            I => \N__8680\
        );

    \I__1920\ : ClkMux
    port map (
            O => \N__8795\,
            I => \N__8680\
        );

    \I__1919\ : ClkMux
    port map (
            O => \N__8794\,
            I => \N__8680\
        );

    \I__1918\ : ClkMux
    port map (
            O => \N__8793\,
            I => \N__8680\
        );

    \I__1917\ : ClkMux
    port map (
            O => \N__8792\,
            I => \N__8680\
        );

    \I__1916\ : ClkMux
    port map (
            O => \N__8791\,
            I => \N__8680\
        );

    \I__1915\ : ClkMux
    port map (
            O => \N__8790\,
            I => \N__8680\
        );

    \I__1914\ : ClkMux
    port map (
            O => \N__8789\,
            I => \N__8680\
        );

    \I__1913\ : ClkMux
    port map (
            O => \N__8788\,
            I => \N__8680\
        );

    \I__1912\ : ClkMux
    port map (
            O => \N__8787\,
            I => \N__8680\
        );

    \I__1911\ : ClkMux
    port map (
            O => \N__8786\,
            I => \N__8680\
        );

    \I__1910\ : ClkMux
    port map (
            O => \N__8785\,
            I => \N__8680\
        );

    \I__1909\ : ClkMux
    port map (
            O => \N__8784\,
            I => \N__8680\
        );

    \I__1908\ : ClkMux
    port map (
            O => \N__8783\,
            I => \N__8680\
        );

    \I__1907\ : ClkMux
    port map (
            O => \N__8782\,
            I => \N__8680\
        );

    \I__1906\ : ClkMux
    port map (
            O => \N__8781\,
            I => \N__8680\
        );

    \I__1905\ : ClkMux
    port map (
            O => \N__8780\,
            I => \N__8680\
        );

    \I__1904\ : ClkMux
    port map (
            O => \N__8779\,
            I => \N__8680\
        );

    \I__1903\ : ClkMux
    port map (
            O => \N__8778\,
            I => \N__8680\
        );

    \I__1902\ : ClkMux
    port map (
            O => \N__8777\,
            I => \N__8680\
        );

    \I__1901\ : ClkMux
    port map (
            O => \N__8776\,
            I => \N__8680\
        );

    \I__1900\ : ClkMux
    port map (
            O => \N__8775\,
            I => \N__8680\
        );

    \I__1899\ : ClkMux
    port map (
            O => \N__8774\,
            I => \N__8680\
        );

    \I__1898\ : ClkMux
    port map (
            O => \N__8773\,
            I => \N__8680\
        );

    \I__1897\ : Glb2LocalMux
    port map (
            O => \N__8770\,
            I => \N__8680\
        );

    \I__1896\ : ClkMux
    port map (
            O => \N__8769\,
            I => \N__8680\
        );

    \I__1895\ : ClkMux
    port map (
            O => \N__8768\,
            I => \N__8680\
        );

    \I__1894\ : ClkMux
    port map (
            O => \N__8767\,
            I => \N__8680\
        );

    \I__1893\ : ClkMux
    port map (
            O => \N__8766\,
            I => \N__8680\
        );

    \I__1892\ : ClkMux
    port map (
            O => \N__8765\,
            I => \N__8680\
        );

    \I__1891\ : ClkMux
    port map (
            O => \N__8764\,
            I => \N__8680\
        );

    \I__1890\ : ClkMux
    port map (
            O => \N__8763\,
            I => \N__8680\
        );

    \I__1889\ : ClkMux
    port map (
            O => \N__8762\,
            I => \N__8680\
        );

    \I__1888\ : ClkMux
    port map (
            O => \N__8761\,
            I => \N__8680\
        );

    \I__1887\ : ClkMux
    port map (
            O => \N__8760\,
            I => \N__8680\
        );

    \I__1886\ : ClkMux
    port map (
            O => \N__8759\,
            I => \N__8680\
        );

    \I__1885\ : GlobalMux
    port map (
            O => \N__8680\,
            I => \CLK80_PLL\
        );

    \I__1884\ : CEMux
    port map (
            O => \N__8677\,
            I => \N__8671\
        );

    \I__1883\ : CEMux
    port map (
            O => \N__8676\,
            I => \N__8668\
        );

    \I__1882\ : CEMux
    port map (
            O => \N__8675\,
            I => \N__8664\
        );

    \I__1881\ : CEMux
    port map (
            O => \N__8674\,
            I => \N__8660\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__8671\,
            I => \N__8655\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__8668\,
            I => \N__8655\
        );

    \I__1878\ : CEMux
    port map (
            O => \N__8667\,
            I => \N__8652\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__8664\,
            I => \N__8649\
        );

    \I__1876\ : CEMux
    port map (
            O => \N__8663\,
            I => \N__8646\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__8660\,
            I => \N__8643\
        );

    \I__1874\ : Span4Mux_v
    port map (
            O => \N__8655\,
            I => \N__8638\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__8652\,
            I => \N__8638\
        );

    \I__1872\ : Span4Mux_h
    port map (
            O => \N__8649\,
            I => \N__8633\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__8646\,
            I => \N__8633\
        );

    \I__1870\ : Span4Mux_h
    port map (
            O => \N__8643\,
            I => \N__8630\
        );

    \I__1869\ : Span4Mux_v
    port map (
            O => \N__8638\,
            I => \N__8627\
        );

    \I__1868\ : Span4Mux_h
    port map (
            O => \N__8633\,
            I => \N__8624\
        );

    \I__1867\ : Odrv4
    port map (
            O => \N__8630\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__8627\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1865\ : Odrv4
    port map (
            O => \N__8624\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1864\ : InMux
    port map (
            O => \N__8617\,
            I => \N__8614\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__8614\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__1862\ : IoInMux
    port map (
            O => \N__8611\,
            I => \N__8608\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__8608\,
            I => \N__8605\
        );

    \I__1860\ : IoSpan4Mux
    port map (
            O => \N__8605\,
            I => \N__8602\
        );

    \I__1859\ : Span4Mux_s2_h
    port map (
            O => \N__8602\,
            I => \N__8599\
        );

    \I__1858\ : Sp12to4
    port map (
            O => \N__8599\,
            I => \N__8596\
        );

    \I__1857\ : Span12Mux_h
    port map (
            O => \N__8596\,
            I => \N__8593\
        );

    \I__1856\ : Odrv12
    port map (
            O => \N__8593\,
            I => \CMA_c_6\
        );

    \I__1855\ : InMux
    port map (
            O => \N__8590\,
            I => \N__8587\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__8587\,
            I => \N__8584\
        );

    \I__1853\ : Span4Mux_v
    port map (
            O => \N__8584\,
            I => \N__8581\
        );

    \I__1852\ : Span4Mux_v
    port map (
            O => \N__8581\,
            I => \N__8578\
        );

    \I__1851\ : Sp12to4
    port map (
            O => \N__8578\,
            I => \N__8575\
        );

    \I__1850\ : Span12Mux_h
    port map (
            O => \N__8575\,
            I => \N__8572\
        );

    \I__1849\ : Odrv12
    port map (
            O => \N__8572\,
            I => \A_c_17\
        );

    \I__1848\ : IoInMux
    port map (
            O => \N__8569\,
            I => \N__8566\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__8566\,
            I => \N__8563\
        );

    \I__1846\ : Span4Mux_s3_h
    port map (
            O => \N__8563\,
            I => \N__8560\
        );

    \I__1845\ : Sp12to4
    port map (
            O => \N__8560\,
            I => \N__8557\
        );

    \I__1844\ : Span12Mux_s9_v
    port map (
            O => \N__8557\,
            I => \N__8554\
        );

    \I__1843\ : Span12Mux_h
    port map (
            O => \N__8554\,
            I => \N__8551\
        );

    \I__1842\ : Odrv12
    port map (
            O => \N__8551\,
            I => \CMA_c_8\
        );

    \I__1841\ : InMux
    port map (
            O => \N__8548\,
            I => \N__8545\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__8545\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__1839\ : IoInMux
    port map (
            O => \N__8542\,
            I => \N__8539\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__8539\,
            I => \N__8536\
        );

    \I__1837\ : Span12Mux_s3_h
    port map (
            O => \N__8536\,
            I => \N__8533\
        );

    \I__1836\ : Span12Mux_h
    port map (
            O => \N__8533\,
            I => \N__8530\
        );

    \I__1835\ : Odrv12
    port map (
            O => \N__8530\,
            I => \CMA_c_7\
        );

    \I__1834\ : InMux
    port map (
            O => \N__8527\,
            I => \N__8524\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__8524\,
            I => \N__8520\
        );

    \I__1832\ : InMux
    port map (
            O => \N__8523\,
            I => \N__8517\
        );

    \I__1831\ : Odrv4
    port map (
            O => \N__8520\,
            I => \U712_CHIP_RAM.CMA_5_i_0_8\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8517\,
            I => \U712_CHIP_RAM.CMA_5_i_0_8\
        );

    \I__1829\ : InMux
    port map (
            O => \N__8512\,
            I => \N__8509\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__8509\,
            I => \N__8506\
        );

    \I__1827\ : Span4Mux_v
    port map (
            O => \N__8506\,
            I => \N__8503\
        );

    \I__1826\ : Span4Mux_v
    port map (
            O => \N__8503\,
            I => \N__8500\
        );

    \I__1825\ : Sp12to4
    port map (
            O => \N__8500\,
            I => \N__8497\
        );

    \I__1824\ : Span12Mux_h
    port map (
            O => \N__8497\,
            I => \N__8494\
        );

    \I__1823\ : Odrv12
    port map (
            O => \N__8494\,
            I => \A_c_19\
        );

    \I__1822\ : IoInMux
    port map (
            O => \N__8491\,
            I => \N__8488\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__8488\,
            I => \N__8485\
        );

    \I__1820\ : Span4Mux_s3_h
    port map (
            O => \N__8485\,
            I => \N__8482\
        );

    \I__1819\ : Sp12to4
    port map (
            O => \N__8482\,
            I => \N__8479\
        );

    \I__1818\ : Span12Mux_s11_v
    port map (
            O => \N__8479\,
            I => \N__8476\
        );

    \I__1817\ : Odrv12
    port map (
            O => \N__8476\,
            I => \CMA_c_9\
        );

    \I__1816\ : InMux
    port map (
            O => \N__8473\,
            I => \N__8470\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__8470\,
            I => \N__8467\
        );

    \I__1814\ : Odrv4
    port map (
            O => \N__8467\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__1813\ : IoInMux
    port map (
            O => \N__8464\,
            I => \N__8461\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__8461\,
            I => \N__8458\
        );

    \I__1811\ : Span4Mux_s2_h
    port map (
            O => \N__8458\,
            I => \N__8455\
        );

    \I__1810\ : Span4Mux_v
    port map (
            O => \N__8455\,
            I => \N__8452\
        );

    \I__1809\ : Sp12to4
    port map (
            O => \N__8452\,
            I => \N__8449\
        );

    \I__1808\ : Span12Mux_h
    port map (
            O => \N__8449\,
            I => \N__8446\
        );

    \I__1807\ : Odrv12
    port map (
            O => \N__8446\,
            I => \CMA_c_3\
        );

    \I__1806\ : InMux
    port map (
            O => \N__8443\,
            I => \N__8440\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__8440\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__1804\ : InMux
    port map (
            O => \N__8437\,
            I => \N__8434\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__8434\,
            I => \N__8431\
        );

    \I__1802\ : Odrv4
    port map (
            O => \N__8431\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8428\,
            I => \N__8425\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__8425\,
            I => \N__8422\
        );

    \I__1799\ : Odrv4
    port map (
            O => \N__8422\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__1798\ : CascadeMux
    port map (
            O => \N__8419\,
            I => \N__8416\
        );

    \I__1797\ : InMux
    port map (
            O => \N__8416\,
            I => \N__8413\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__8413\,
            I => \N__8410\
        );

    \I__1795\ : Odrv4
    port map (
            O => \N__8410\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__1794\ : CascadeMux
    port map (
            O => \N__8407\,
            I => \U712_BYTE_ENABLE.N_563_cascade_\
        );

    \I__1793\ : IoInMux
    port map (
            O => \N__8404\,
            I => \N__8401\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__8401\,
            I => \N__8398\
        );

    \I__1791\ : Span4Mux_s2_v
    port map (
            O => \N__8398\,
            I => \N__8395\
        );

    \I__1790\ : Span4Mux_h
    port map (
            O => \N__8395\,
            I => \N__8392\
        );

    \I__1789\ : Sp12to4
    port map (
            O => \N__8392\,
            I => \N__8389\
        );

    \I__1788\ : Span12Mux_s10_v
    port map (
            O => \N__8389\,
            I => \N__8386\
        );

    \I__1787\ : Odrv12
    port map (
            O => \N__8386\,
            I => \N_56_i\
        );

    \I__1786\ : IoInMux
    port map (
            O => \N__8383\,
            I => \N__8380\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__8380\,
            I => \N__8377\
        );

    \I__1784\ : IoSpan4Mux
    port map (
            O => \N__8377\,
            I => \N__8374\
        );

    \I__1783\ : Sp12to4
    port map (
            O => \N__8374\,
            I => \N__8371\
        );

    \I__1782\ : Span12Mux_s7_v
    port map (
            O => \N__8371\,
            I => \N__8368\
        );

    \I__1781\ : Odrv12
    port map (
            O => \N__8368\,
            I => \WEn_c\
        );

    \I__1780\ : InMux
    port map (
            O => \N__8365\,
            I => \N__8361\
        );

    \I__1779\ : InMux
    port map (
            O => \N__8364\,
            I => \N__8358\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__8361\,
            I => \N__8355\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__8358\,
            I => \N__8347\
        );

    \I__1776\ : Span4Mux_h
    port map (
            O => \N__8355\,
            I => \N__8347\
        );

    \I__1775\ : InMux
    port map (
            O => \N__8354\,
            I => \N__8344\
        );

    \I__1774\ : InMux
    port map (
            O => \N__8353\,
            I => \N__8341\
        );

    \I__1773\ : CascadeMux
    port map (
            O => \N__8352\,
            I => \N__8338\
        );

    \I__1772\ : Span4Mux_v
    port map (
            O => \N__8347\,
            I => \N__8331\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__8344\,
            I => \N__8331\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__8341\,
            I => \N__8331\
        );

    \I__1769\ : InMux
    port map (
            O => \N__8338\,
            I => \N__8328\
        );

    \I__1768\ : Span4Mux_h
    port map (
            O => \N__8331\,
            I => \N__8325\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__8328\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1766\ : Odrv4
    port map (
            O => \N__8325\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1765\ : IoInMux
    port map (
            O => \N__8320\,
            I => \N__8317\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8317\,
            I => \N__8314\
        );

    \I__1763\ : Span4Mux_s3_v
    port map (
            O => \N__8314\,
            I => \N__8311\
        );

    \I__1762\ : Span4Mux_v
    port map (
            O => \N__8311\,
            I => \N__8308\
        );

    \I__1761\ : Span4Mux_h
    port map (
            O => \N__8308\,
            I => \N__8305\
        );

    \I__1760\ : Odrv4
    port map (
            O => \N__8305\,
            I => \CRCSn_c\
        );

    \I__1759\ : InMux
    port map (
            O => \N__8302\,
            I => \N__8299\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__8299\,
            I => \N__8292\
        );

    \I__1757\ : InMux
    port map (
            O => \N__8298\,
            I => \N__8289\
        );

    \I__1756\ : InMux
    port map (
            O => \N__8297\,
            I => \N__8286\
        );

    \I__1755\ : CascadeMux
    port map (
            O => \N__8296\,
            I => \N__8283\
        );

    \I__1754\ : CascadeMux
    port map (
            O => \N__8295\,
            I => \N__8280\
        );

    \I__1753\ : Span4Mux_h
    port map (
            O => \N__8292\,
            I => \N__8277\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__8289\,
            I => \N__8274\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__8286\,
            I => \N__8271\
        );

    \I__1750\ : InMux
    port map (
            O => \N__8283\,
            I => \N__8268\
        );

    \I__1749\ : InMux
    port map (
            O => \N__8280\,
            I => \N__8265\
        );

    \I__1748\ : Span4Mux_v
    port map (
            O => \N__8277\,
            I => \N__8262\
        );

    \I__1747\ : Span4Mux_v
    port map (
            O => \N__8274\,
            I => \N__8259\
        );

    \I__1746\ : Span4Mux_h
    port map (
            O => \N__8271\,
            I => \N__8254\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__8268\,
            I => \N__8254\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__8265\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1743\ : Odrv4
    port map (
            O => \N__8262\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1742\ : Odrv4
    port map (
            O => \N__8259\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1741\ : Odrv4
    port map (
            O => \N__8254\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1740\ : InMux
    port map (
            O => \N__8245\,
            I => \N__8242\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__8242\,
            I => \N__8239\
        );

    \I__1738\ : Odrv12
    port map (
            O => \N__8239\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__1737\ : InMux
    port map (
            O => \N__8236\,
            I => \N__8233\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__8233\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\
        );

    \I__1735\ : InMux
    port map (
            O => \N__8230\,
            I => \N__8227\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__8227\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\
        );

    \I__1733\ : InMux
    port map (
            O => \N__8224\,
            I => \N__8221\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__8221\,
            I => \N__8218\
        );

    \I__1731\ : Odrv12
    port map (
            O => \N__8218\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\
        );

    \I__1730\ : IoInMux
    port map (
            O => \N__8215\,
            I => \N__8212\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__8212\,
            I => \N__8209\
        );

    \I__1728\ : IoSpan4Mux
    port map (
            O => \N__8209\,
            I => \N__8206\
        );

    \I__1727\ : Span4Mux_s2_h
    port map (
            O => \N__8206\,
            I => \N__8203\
        );

    \I__1726\ : Sp12to4
    port map (
            O => \N__8203\,
            I => \N__8200\
        );

    \I__1725\ : Span12Mux_h
    port map (
            O => \N__8200\,
            I => \N__8197\
        );

    \I__1724\ : Odrv12
    port map (
            O => \N__8197\,
            I => \CMA_c_5\
        );

    \I__1723\ : CascadeMux
    port map (
            O => \N__8194\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\
        );

    \I__1722\ : InMux
    port map (
            O => \N__8191\,
            I => \N__8188\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__8188\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__1720\ : InMux
    port map (
            O => \N__8185\,
            I => \N__8179\
        );

    \I__1719\ : InMux
    port map (
            O => \N__8184\,
            I => \N__8176\
        );

    \I__1718\ : InMux
    port map (
            O => \N__8183\,
            I => \N__8173\
        );

    \I__1717\ : InMux
    port map (
            O => \N__8182\,
            I => \N__8170\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__8179\,
            I => \N__8163\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__8176\,
            I => \N__8163\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__8173\,
            I => \N__8163\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__8170\,
            I => \N__8158\
        );

    \I__1712\ : Span4Mux_h
    port map (
            O => \N__8163\,
            I => \N__8158\
        );

    \I__1711\ : Sp12to4
    port map (
            O => \N__8158\,
            I => \N__8155\
        );

    \I__1710\ : Span12Mux_v
    port map (
            O => \N__8155\,
            I => \N__8152\
        );

    \I__1709\ : Odrv12
    port map (
            O => \N__8152\,
            I => \CLK40_PLL_i\
        );

    \I__1708\ : IoInMux
    port map (
            O => \N__8149\,
            I => \N__8145\
        );

    \I__1707\ : IoInMux
    port map (
            O => \N__8148\,
            I => \N__8142\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__8145\,
            I => \N__8138\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__8142\,
            I => \N__8135\
        );

    \I__1704\ : IoInMux
    port map (
            O => \N__8141\,
            I => \N__8132\
        );

    \I__1703\ : Span4Mux_s2_v
    port map (
            O => \N__8138\,
            I => \N__8129\
        );

    \I__1702\ : Span4Mux_s2_v
    port map (
            O => \N__8135\,
            I => \N__8126\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__8132\,
            I => \N__8123\
        );

    \I__1700\ : Span4Mux_v
    port map (
            O => \N__8129\,
            I => \N__8120\
        );

    \I__1699\ : Span4Mux_v
    port map (
            O => \N__8126\,
            I => \N__8117\
        );

    \I__1698\ : Span4Mux_s3_h
    port map (
            O => \N__8123\,
            I => \N__8114\
        );

    \I__1697\ : Sp12to4
    port map (
            O => \N__8120\,
            I => \N__8109\
        );

    \I__1696\ : Sp12to4
    port map (
            O => \N__8117\,
            I => \N__8109\
        );

    \I__1695\ : Span4Mux_h
    port map (
            O => \N__8114\,
            I => \N__8106\
        );

    \I__1694\ : Span12Mux_s8_h
    port map (
            O => \N__8109\,
            I => \N__8103\
        );

    \I__1693\ : Span4Mux_h
    port map (
            O => \N__8106\,
            I => \N__8100\
        );

    \I__1692\ : Span12Mux_v
    port map (
            O => \N__8103\,
            I => \N__8097\
        );

    \I__1691\ : Span4Mux_h
    port map (
            O => \N__8100\,
            I => \N__8094\
        );

    \I__1690\ : Odrv12
    port map (
            O => \N__8097\,
            I => \CLK40_PLL_i_i\
        );

    \I__1689\ : Odrv4
    port map (
            O => \N__8094\,
            I => \CLK40_PLL_i_i\
        );

    \I__1688\ : InMux
    port map (
            O => \N__8089\,
            I => \N__8085\
        );

    \I__1687\ : InMux
    port map (
            O => \N__8088\,
            I => \N__8082\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__8085\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__8082\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1684\ : InMux
    port map (
            O => \N__8077\,
            I => \N__8074\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__8074\,
            I => \U712_CYCLE_TERM.N_598\
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__8071\,
            I => \N__8066\
        );

    \I__1681\ : InMux
    port map (
            O => \N__8070\,
            I => \N__8063\
        );

    \I__1680\ : InMux
    port map (
            O => \N__8069\,
            I => \N__8060\
        );

    \I__1679\ : InMux
    port map (
            O => \N__8066\,
            I => \N__8057\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__8063\,
            I => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__8060\,
            I => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__8057\,
            I => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\
        );

    \I__1675\ : InMux
    port map (
            O => \N__8050\,
            I => \N__8046\
        );

    \I__1674\ : InMux
    port map (
            O => \N__8049\,
            I => \N__8043\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__8046\,
            I => \U712_CYCLE_TERM.N_440\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__8043\,
            I => \U712_CYCLE_TERM.N_440\
        );

    \I__1671\ : InMux
    port map (
            O => \N__8038\,
            I => \N__8035\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__8035\,
            I => \U712_CYCLE_TERM.un13_0\
        );

    \I__1669\ : InMux
    port map (
            O => \N__8032\,
            I => \N__8015\
        );

    \I__1668\ : InMux
    port map (
            O => \N__8031\,
            I => \N__8015\
        );

    \I__1667\ : InMux
    port map (
            O => \N__8030\,
            I => \N__8015\
        );

    \I__1666\ : InMux
    port map (
            O => \N__8029\,
            I => \N__8008\
        );

    \I__1665\ : InMux
    port map (
            O => \N__8028\,
            I => \N__8008\
        );

    \I__1664\ : InMux
    port map (
            O => \N__8027\,
            I => \N__8008\
        );

    \I__1663\ : InMux
    port map (
            O => \N__8026\,
            I => \N__8004\
        );

    \I__1662\ : InMux
    port map (
            O => \N__8025\,
            I => \N__8001\
        );

    \I__1661\ : InMux
    port map (
            O => \N__8024\,
            I => \N__7996\
        );

    \I__1660\ : InMux
    port map (
            O => \N__8023\,
            I => \N__7991\
        );

    \I__1659\ : InMux
    port map (
            O => \N__8022\,
            I => \N__7991\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__8015\,
            I => \N__7979\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__8008\,
            I => \N__7979\
        );

    \I__1656\ : InMux
    port map (
            O => \N__8007\,
            I => \N__7976\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__8004\,
            I => \N__7972\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__8001\,
            I => \N__7969\
        );

    \I__1653\ : InMux
    port map (
            O => \N__8000\,
            I => \N__7964\
        );

    \I__1652\ : InMux
    port map (
            O => \N__7999\,
            I => \N__7964\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__7996\,
            I => \N__7954\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__7991\,
            I => \N__7954\
        );

    \I__1649\ : InMux
    port map (
            O => \N__7990\,
            I => \N__7951\
        );

    \I__1648\ : InMux
    port map (
            O => \N__7989\,
            I => \N__7944\
        );

    \I__1647\ : InMux
    port map (
            O => \N__7988\,
            I => \N__7944\
        );

    \I__1646\ : InMux
    port map (
            O => \N__7987\,
            I => \N__7941\
        );

    \I__1645\ : InMux
    port map (
            O => \N__7986\,
            I => \N__7938\
        );

    \I__1644\ : InMux
    port map (
            O => \N__7985\,
            I => \N__7933\
        );

    \I__1643\ : InMux
    port map (
            O => \N__7984\,
            I => \N__7933\
        );

    \I__1642\ : Span4Mux_v
    port map (
            O => \N__7979\,
            I => \N__7928\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__7976\,
            I => \N__7928\
        );

    \I__1640\ : InMux
    port map (
            O => \N__7975\,
            I => \N__7925\
        );

    \I__1639\ : Span4Mux_v
    port map (
            O => \N__7972\,
            I => \N__7917\
        );

    \I__1638\ : Span4Mux_v
    port map (
            O => \N__7969\,
            I => \N__7917\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__7964\,
            I => \N__7917\
        );

    \I__1636\ : InMux
    port map (
            O => \N__7963\,
            I => \N__7908\
        );

    \I__1635\ : InMux
    port map (
            O => \N__7962\,
            I => \N__7908\
        );

    \I__1634\ : InMux
    port map (
            O => \N__7961\,
            I => \N__7908\
        );

    \I__1633\ : InMux
    port map (
            O => \N__7960\,
            I => \N__7908\
        );

    \I__1632\ : InMux
    port map (
            O => \N__7959\,
            I => \N__7905\
        );

    \I__1631\ : Span4Mux_v
    port map (
            O => \N__7954\,
            I => \N__7900\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__7951\,
            I => \N__7900\
        );

    \I__1629\ : InMux
    port map (
            O => \N__7950\,
            I => \N__7897\
        );

    \I__1628\ : InMux
    port map (
            O => \N__7949\,
            I => \N__7894\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__7944\,
            I => \N__7885\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__7941\,
            I => \N__7885\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__7938\,
            I => \N__7885\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__7933\,
            I => \N__7885\
        );

    \I__1623\ : Span4Mux_v
    port map (
            O => \N__7928\,
            I => \N__7880\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__7925\,
            I => \N__7880\
        );

    \I__1621\ : InMux
    port map (
            O => \N__7924\,
            I => \N__7877\
        );

    \I__1620\ : Span4Mux_h
    port map (
            O => \N__7917\,
            I => \N__7872\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__7908\,
            I => \N__7872\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__7905\,
            I => \N__7865\
        );

    \I__1617\ : Span4Mux_v
    port map (
            O => \N__7900\,
            I => \N__7865\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__7897\,
            I => \N__7865\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__7894\,
            I => \N__7862\
        );

    \I__1614\ : Span4Mux_v
    port map (
            O => \N__7885\,
            I => \N__7857\
        );

    \I__1613\ : Span4Mux_v
    port map (
            O => \N__7880\,
            I => \N__7857\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__7877\,
            I => \N__7854\
        );

    \I__1611\ : Span4Mux_v
    port map (
            O => \N__7872\,
            I => \N__7847\
        );

    \I__1610\ : Span4Mux_v
    port map (
            O => \N__7865\,
            I => \N__7847\
        );

    \I__1609\ : Span4Mux_v
    port map (
            O => \N__7862\,
            I => \N__7847\
        );

    \I__1608\ : Sp12to4
    port map (
            O => \N__7857\,
            I => \N__7844\
        );

    \I__1607\ : Span12Mux_v
    port map (
            O => \N__7854\,
            I => \N__7839\
        );

    \I__1606\ : Sp12to4
    port map (
            O => \N__7847\,
            I => \N__7839\
        );

    \I__1605\ : Span12Mux_h
    port map (
            O => \N__7844\,
            I => \N__7836\
        );

    \I__1604\ : Span12Mux_h
    port map (
            O => \N__7839\,
            I => \N__7833\
        );

    \I__1603\ : Odrv12
    port map (
            O => \N__7836\,
            I => \RESETn_c\
        );

    \I__1602\ : Odrv12
    port map (
            O => \N__7833\,
            I => \RESETn_c\
        );

    \I__1601\ : InMux
    port map (
            O => \N__7828\,
            I => \N__7825\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__7825\,
            I => \U712_CYCLE_TERM.N_566\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__7822\,
            I => \U712_CYCLE_TERM.un13_0_cascade_\
        );

    \I__1598\ : CascadeMux
    port map (
            O => \N__7819\,
            I => \N__7816\
        );

    \I__1597\ : InMux
    port map (
            O => \N__7816\,
            I => \N__7813\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__7813\,
            I => \N__7810\
        );

    \I__1595\ : Odrv12
    port map (
            O => \N__7810\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\
        );

    \I__1594\ : InMux
    port map (
            O => \N__7807\,
            I => \N__7804\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__7804\,
            I => \N__7797\
        );

    \I__1592\ : CascadeMux
    port map (
            O => \N__7803\,
            I => \N__7787\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__7802\,
            I => \N__7784\
        );

    \I__1590\ : InMux
    port map (
            O => \N__7801\,
            I => \N__7779\
        );

    \I__1589\ : InMux
    port map (
            O => \N__7800\,
            I => \N__7776\
        );

    \I__1588\ : Span4Mux_h
    port map (
            O => \N__7797\,
            I => \N__7773\
        );

    \I__1587\ : InMux
    port map (
            O => \N__7796\,
            I => \N__7768\
        );

    \I__1586\ : InMux
    port map (
            O => \N__7795\,
            I => \N__7768\
        );

    \I__1585\ : InMux
    port map (
            O => \N__7794\,
            I => \N__7765\
        );

    \I__1584\ : InMux
    port map (
            O => \N__7793\,
            I => \N__7760\
        );

    \I__1583\ : InMux
    port map (
            O => \N__7792\,
            I => \N__7760\
        );

    \I__1582\ : InMux
    port map (
            O => \N__7791\,
            I => \N__7753\
        );

    \I__1581\ : InMux
    port map (
            O => \N__7790\,
            I => \N__7753\
        );

    \I__1580\ : InMux
    port map (
            O => \N__7787\,
            I => \N__7753\
        );

    \I__1579\ : InMux
    port map (
            O => \N__7784\,
            I => \N__7746\
        );

    \I__1578\ : InMux
    port map (
            O => \N__7783\,
            I => \N__7746\
        );

    \I__1577\ : InMux
    port map (
            O => \N__7782\,
            I => \N__7746\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__7779\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__7776\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1574\ : Odrv4
    port map (
            O => \N__7773\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__7768\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__7765\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__7760\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__7753\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__7746\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1568\ : InMux
    port map (
            O => \N__7729\,
            I => \N__7726\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__7726\,
            I => \N__7723\
        );

    \I__1566\ : Span4Mux_h
    port map (
            O => \N__7723\,
            I => \N__7720\
        );

    \I__1565\ : Odrv4
    port map (
            O => \N__7720\,
            I => \U712_CHIP_RAM.N_93\
        );

    \I__1564\ : IoInMux
    port map (
            O => \N__7717\,
            I => \N__7714\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__7714\,
            I => \N__7711\
        );

    \I__1562\ : IoSpan4Mux
    port map (
            O => \N__7711\,
            I => \N__7707\
        );

    \I__1561\ : InMux
    port map (
            O => \N__7710\,
            I => \N__7704\
        );

    \I__1560\ : Span4Mux_s2_v
    port map (
            O => \N__7707\,
            I => \N__7701\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__7704\,
            I => \N__7698\
        );

    \I__1558\ : Sp12to4
    port map (
            O => \N__7701\,
            I => \N__7695\
        );

    \I__1557\ : Span4Mux_v
    port map (
            O => \N__7698\,
            I => \N__7692\
        );

    \I__1556\ : Span12Mux_s8_v
    port map (
            O => \N__7695\,
            I => \N__7689\
        );

    \I__1555\ : Sp12to4
    port map (
            O => \N__7692\,
            I => \N__7686\
        );

    \I__1554\ : Span12Mux_v
    port map (
            O => \N__7689\,
            I => \N__7681\
        );

    \I__1553\ : Span12Mux_h
    port map (
            O => \N__7686\,
            I => \N__7681\
        );

    \I__1552\ : Span12Mux_h
    port map (
            O => \N__7681\,
            I => \N__7678\
        );

    \I__1551\ : Odrv12
    port map (
            O => \N__7678\,
            I => \A_c_10\
        );

    \I__1550\ : InMux
    port map (
            O => \N__7675\,
            I => \N__7672\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__7672\,
            I => \N__7669\
        );

    \I__1548\ : Odrv12
    port map (
            O => \N__7669\,
            I => \U712_CHIP_RAM.N_455\
        );

    \I__1547\ : IoInMux
    port map (
            O => \N__7666\,
            I => \N__7662\
        );

    \I__1546\ : InMux
    port map (
            O => \N__7665\,
            I => \N__7659\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__7662\,
            I => \N__7656\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__7659\,
            I => \N__7653\
        );

    \I__1543\ : Span12Mux_s9_h
    port map (
            O => \N__7656\,
            I => \N__7649\
        );

    \I__1542\ : Span4Mux_v
    port map (
            O => \N__7653\,
            I => \N__7646\
        );

    \I__1541\ : InMux
    port map (
            O => \N__7652\,
            I => \N__7643\
        );

    \I__1540\ : Span12Mux_v
    port map (
            O => \N__7649\,
            I => \N__7639\
        );

    \I__1539\ : Span4Mux_h
    port map (
            O => \N__7646\,
            I => \N__7636\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7643\,
            I => \N__7633\
        );

    \I__1537\ : InMux
    port map (
            O => \N__7642\,
            I => \N__7630\
        );

    \I__1536\ : Odrv12
    port map (
            O => \N__7639\,
            I => \TACK_OUTn\
        );

    \I__1535\ : Odrv4
    port map (
            O => \N__7636\,
            I => \TACK_OUTn\
        );

    \I__1534\ : Odrv4
    port map (
            O => \N__7633\,
            I => \TACK_OUTn\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__7630\,
            I => \TACK_OUTn\
        );

    \I__1532\ : InMux
    port map (
            O => \N__7621\,
            I => \N__7617\
        );

    \I__1531\ : InMux
    port map (
            O => \N__7620\,
            I => \N__7614\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__7617\,
            I => \U712_CYCLE_TERM.RAM_CYCLEZ0\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__7614\,
            I => \U712_CYCLE_TERM.RAM_CYCLEZ0\
        );

    \I__1528\ : IoInMux
    port map (
            O => \N__7609\,
            I => \N__7606\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7606\,
            I => \N__7603\
        );

    \I__1526\ : Span4Mux_s3_h
    port map (
            O => \N__7603\,
            I => \N__7600\
        );

    \I__1525\ : Span4Mux_h
    port map (
            O => \N__7600\,
            I => \N__7596\
        );

    \I__1524\ : InMux
    port map (
            O => \N__7599\,
            I => \N__7593\
        );

    \I__1523\ : Sp12to4
    port map (
            O => \N__7596\,
            I => \N__7590\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__7593\,
            I => \N__7587\
        );

    \I__1521\ : Span12Mux_v
    port map (
            O => \N__7590\,
            I => \N__7580\
        );

    \I__1520\ : Span12Mux_s7_h
    port map (
            O => \N__7587\,
            I => \N__7580\
        );

    \I__1519\ : InMux
    port map (
            O => \N__7586\,
            I => \N__7577\
        );

    \I__1518\ : InMux
    port map (
            O => \N__7585\,
            I => \N__7574\
        );

    \I__1517\ : Odrv12
    port map (
            O => \N__7580\,
            I => \TACK_EN\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__7577\,
            I => \TACK_EN\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__7574\,
            I => \TACK_EN\
        );

    \I__1514\ : IoInMux
    port map (
            O => \N__7567\,
            I => \N__7564\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__7564\,
            I => \N__7561\
        );

    \I__1512\ : Span4Mux_s2_v
    port map (
            O => \N__7561\,
            I => \N__7558\
        );

    \I__1511\ : Sp12to4
    port map (
            O => \N__7558\,
            I => \N__7555\
        );

    \I__1510\ : Span12Mux_s11_h
    port map (
            O => \N__7555\,
            I => \N__7552\
        );

    \I__1509\ : Span12Mux_v
    port map (
            O => \N__7552\,
            I => \N__7549\
        );

    \I__1508\ : Odrv12
    port map (
            O => \N__7549\,
            I => \U712_CYCLE_TERM_TCIn_0_i\
        );

    \I__1507\ : IoInMux
    port map (
            O => \N__7546\,
            I => \N__7543\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__7543\,
            I => \N__7540\
        );

    \I__1505\ : Span4Mux_s2_v
    port map (
            O => \N__7540\,
            I => \N__7537\
        );

    \I__1504\ : Span4Mux_h
    port map (
            O => \N__7537\,
            I => \N__7534\
        );

    \I__1503\ : Sp12to4
    port map (
            O => \N__7534\,
            I => \N__7530\
        );

    \I__1502\ : InMux
    port map (
            O => \N__7533\,
            I => \N__7527\
        );

    \I__1501\ : Span12Mux_s9_v
    port map (
            O => \N__7530\,
            I => \N__7524\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__7527\,
            I => \N__7521\
        );

    \I__1499\ : Odrv12
    port map (
            O => \N__7524\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1498\ : Odrv12
    port map (
            O => \N__7521\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1497\ : CascadeMux
    port map (
            O => \N__7516\,
            I => \U712_CHIP_RAM.N_412_cascade_\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7513\,
            I => \N__7510\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__7510\,
            I => \N__7507\
        );

    \I__1494\ : Span4Mux_v
    port map (
            O => \N__7507\,
            I => \N__7504\
        );

    \I__1493\ : Sp12to4
    port map (
            O => \N__7504\,
            I => \N__7501\
        );

    \I__1492\ : Span12Mux_h
    port map (
            O => \N__7501\,
            I => \N__7498\
        );

    \I__1491\ : Span12Mux_v
    port map (
            O => \N__7498\,
            I => \N__7495\
        );

    \I__1490\ : Odrv12
    port map (
            O => \N__7495\,
            I => \A_c_3\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7492\,
            I => \N__7489\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__7489\,
            I => \U712_CHIP_RAM.N_478\
        );

    \I__1487\ : InMux
    port map (
            O => \N__7486\,
            I => \N__7483\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__7483\,
            I => \N__7480\
        );

    \I__1485\ : Span4Mux_h
    port map (
            O => \N__7480\,
            I => \N__7477\
        );

    \I__1484\ : Odrv4
    port map (
            O => \N__7477\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\
        );

    \I__1483\ : InMux
    port map (
            O => \N__7474\,
            I => \N__7471\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__7471\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\
        );

    \I__1481\ : CascadeMux
    port map (
            O => \N__7468\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0_cascade_\
        );

    \I__1480\ : IoInMux
    port map (
            O => \N__7465\,
            I => \N__7462\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__7462\,
            I => \N__7459\
        );

    \I__1478\ : Span12Mux_s11_v
    port map (
            O => \N__7459\,
            I => \N__7456\
        );

    \I__1477\ : Odrv12
    port map (
            O => \N__7456\,
            I => \CMA_c_0\
        );

    \I__1476\ : IoInMux
    port map (
            O => \N__7453\,
            I => \N__7450\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__7450\,
            I => \N__7447\
        );

    \I__1474\ : Span4Mux_s3_v
    port map (
            O => \N__7447\,
            I => \N__7444\
        );

    \I__1473\ : Span4Mux_v
    port map (
            O => \N__7444\,
            I => \N__7441\
        );

    \I__1472\ : Span4Mux_v
    port map (
            O => \N__7441\,
            I => \N__7438\
        );

    \I__1471\ : Odrv4
    port map (
            O => \N__7438\,
            I => \CMA_c_2\
        );

    \I__1470\ : InMux
    port map (
            O => \N__7435\,
            I => \N__7432\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__7432\,
            I => \N__7429\
        );

    \I__1468\ : Span4Mux_v
    port map (
            O => \N__7429\,
            I => \N__7426\
        );

    \I__1467\ : Span4Mux_v
    port map (
            O => \N__7426\,
            I => \N__7423\
        );

    \I__1466\ : Sp12to4
    port map (
            O => \N__7423\,
            I => \N__7420\
        );

    \I__1465\ : Span12Mux_h
    port map (
            O => \N__7420\,
            I => \N__7417\
        );

    \I__1464\ : Odrv12
    port map (
            O => \N__7417\,
            I => \A_c_4\
        );

    \I__1463\ : IoInMux
    port map (
            O => \N__7414\,
            I => \N__7411\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__7411\,
            I => \N__7408\
        );

    \I__1461\ : IoSpan4Mux
    port map (
            O => \N__7408\,
            I => \N__7405\
        );

    \I__1460\ : Span4Mux_s2_v
    port map (
            O => \N__7405\,
            I => \N__7402\
        );

    \I__1459\ : Sp12to4
    port map (
            O => \N__7402\,
            I => \N__7398\
        );

    \I__1458\ : InMux
    port map (
            O => \N__7401\,
            I => \N__7395\
        );

    \I__1457\ : Span12Mux_s8_v
    port map (
            O => \N__7398\,
            I => \N__7392\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__7395\,
            I => \N__7389\
        );

    \I__1455\ : Span12Mux_v
    port map (
            O => \N__7392\,
            I => \N__7386\
        );

    \I__1454\ : Span12Mux_v
    port map (
            O => \N__7389\,
            I => \N__7383\
        );

    \I__1453\ : Span12Mux_h
    port map (
            O => \N__7386\,
            I => \N__7380\
        );

    \I__1452\ : Span12Mux_h
    port map (
            O => \N__7383\,
            I => \N__7377\
        );

    \I__1451\ : Odrv12
    port map (
            O => \N__7380\,
            I => \A_c_11\
        );

    \I__1450\ : Odrv12
    port map (
            O => \N__7377\,
            I => \A_c_11\
        );

    \I__1449\ : InMux
    port map (
            O => \N__7372\,
            I => \N__7367\
        );

    \I__1448\ : InMux
    port map (
            O => \N__7371\,
            I => \N__7362\
        );

    \I__1447\ : InMux
    port map (
            O => \N__7370\,
            I => \N__7362\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__7367\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__7362\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1444\ : CascadeMux
    port map (
            O => \N__7357\,
            I => \N__7354\
        );

    \I__1443\ : InMux
    port map (
            O => \N__7354\,
            I => \N__7351\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__7351\,
            I => \N__7345\
        );

    \I__1441\ : InMux
    port map (
            O => \N__7350\,
            I => \N__7338\
        );

    \I__1440\ : InMux
    port map (
            O => \N__7349\,
            I => \N__7338\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7348\,
            I => \N__7338\
        );

    \I__1438\ : Odrv4
    port map (
            O => \N__7345\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__7338\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1436\ : InMux
    port map (
            O => \N__7333\,
            I => \N__7329\
        );

    \I__1435\ : InMux
    port map (
            O => \N__7332\,
            I => \N__7326\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__7329\,
            I => \U712_REG_SM.N_407\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__7326\,
            I => \U712_REG_SM.N_407\
        );

    \I__1432\ : CascadeMux
    port map (
            O => \N__7321\,
            I => \N__7317\
        );

    \I__1431\ : InMux
    port map (
            O => \N__7320\,
            I => \N__7311\
        );

    \I__1430\ : InMux
    port map (
            O => \N__7317\,
            I => \N__7308\
        );

    \I__1429\ : InMux
    port map (
            O => \N__7316\,
            I => \N__7305\
        );

    \I__1428\ : InMux
    port map (
            O => \N__7315\,
            I => \N__7302\
        );

    \I__1427\ : InMux
    port map (
            O => \N__7314\,
            I => \N__7298\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__7311\,
            I => \N__7295\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__7308\,
            I => \N__7290\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__7305\,
            I => \N__7290\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__7302\,
            I => \N__7287\
        );

    \I__1422\ : InMux
    port map (
            O => \N__7301\,
            I => \N__7284\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__7298\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1420\ : Odrv12
    port map (
            O => \N__7295\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1419\ : Odrv4
    port map (
            O => \N__7290\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1418\ : Odrv4
    port map (
            O => \N__7287\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__7284\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1416\ : CascadeMux
    port map (
            O => \N__7273\,
            I => \N__7269\
        );

    \I__1415\ : InMux
    port map (
            O => \N__7272\,
            I => \N__7261\
        );

    \I__1414\ : InMux
    port map (
            O => \N__7269\,
            I => \N__7256\
        );

    \I__1413\ : InMux
    port map (
            O => \N__7268\,
            I => \N__7256\
        );

    \I__1412\ : InMux
    port map (
            O => \N__7267\,
            I => \N__7247\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7266\,
            I => \N__7247\
        );

    \I__1410\ : InMux
    port map (
            O => \N__7265\,
            I => \N__7247\
        );

    \I__1409\ : InMux
    port map (
            O => \N__7264\,
            I => \N__7247\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__7261\,
            I => \N__7240\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__7256\,
            I => \N__7240\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__7247\,
            I => \N__7240\
        );

    \I__1405\ : Odrv4
    port map (
            O => \N__7240\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1404\ : InMux
    port map (
            O => \N__7237\,
            I => \N__7232\
        );

    \I__1403\ : InMux
    port map (
            O => \N__7236\,
            I => \N__7229\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__7235\,
            I => \N__7225\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__7232\,
            I => \N__7222\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__7229\,
            I => \N__7219\
        );

    \I__1399\ : InMux
    port map (
            O => \N__7228\,
            I => \N__7216\
        );

    \I__1398\ : InMux
    port map (
            O => \N__7225\,
            I => \N__7213\
        );

    \I__1397\ : Sp12to4
    port map (
            O => \N__7222\,
            I => \N__7210\
        );

    \I__1396\ : Sp12to4
    port map (
            O => \N__7219\,
            I => \N__7205\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__7216\,
            I => \N__7205\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__7213\,
            I => \N__7202\
        );

    \I__1393\ : Span12Mux_v
    port map (
            O => \N__7210\,
            I => \N__7199\
        );

    \I__1392\ : Span12Mux_h
    port map (
            O => \N__7205\,
            I => \N__7196\
        );

    \I__1391\ : Span12Mux_v
    port map (
            O => \N__7202\,
            I => \N__7193\
        );

    \I__1390\ : Span12Mux_h
    port map (
            O => \N__7199\,
            I => \N__7188\
        );

    \I__1389\ : Span12Mux_v
    port map (
            O => \N__7196\,
            I => \N__7188\
        );

    \I__1388\ : Span12Mux_h
    port map (
            O => \N__7193\,
            I => \N__7185\
        );

    \I__1387\ : Odrv12
    port map (
            O => \N__7188\,
            I => \RnW_c\
        );

    \I__1386\ : Odrv12
    port map (
            O => \N__7185\,
            I => \RnW_c\
        );

    \I__1385\ : InMux
    port map (
            O => \N__7180\,
            I => \N__7175\
        );

    \I__1384\ : InMux
    port map (
            O => \N__7179\,
            I => \N__7172\
        );

    \I__1383\ : InMux
    port map (
            O => \N__7178\,
            I => \N__7169\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__7175\,
            I => \N__7162\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__7172\,
            I => \N__7162\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__7169\,
            I => \N__7157\
        );

    \I__1379\ : InMux
    port map (
            O => \N__7168\,
            I => \N__7154\
        );

    \I__1378\ : InMux
    port map (
            O => \N__7167\,
            I => \N__7151\
        );

    \I__1377\ : Span4Mux_h
    port map (
            O => \N__7162\,
            I => \N__7148\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7161\,
            I => \N__7145\
        );

    \I__1375\ : InMux
    port map (
            O => \N__7160\,
            I => \N__7140\
        );

    \I__1374\ : Span4Mux_h
    port map (
            O => \N__7157\,
            I => \N__7133\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__7154\,
            I => \N__7133\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__7151\,
            I => \N__7133\
        );

    \I__1371\ : Sp12to4
    port map (
            O => \N__7148\,
            I => \N__7129\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__7145\,
            I => \N__7126\
        );

    \I__1369\ : InMux
    port map (
            O => \N__7144\,
            I => \N__7121\
        );

    \I__1368\ : InMux
    port map (
            O => \N__7143\,
            I => \N__7121\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__7140\,
            I => \N__7118\
        );

    \I__1366\ : Span4Mux_v
    port map (
            O => \N__7133\,
            I => \N__7115\
        );

    \I__1365\ : InMux
    port map (
            O => \N__7132\,
            I => \N__7112\
        );

    \I__1364\ : Odrv12
    port map (
            O => \N__7129\,
            I => \WRITE_CYCLEm\
        );

    \I__1363\ : Odrv4
    port map (
            O => \N__7126\,
            I => \WRITE_CYCLEm\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__7121\,
            I => \WRITE_CYCLEm\
        );

    \I__1361\ : Odrv4
    port map (
            O => \N__7118\,
            I => \WRITE_CYCLEm\
        );

    \I__1360\ : Odrv4
    port map (
            O => \N__7115\,
            I => \WRITE_CYCLEm\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__7112\,
            I => \WRITE_CYCLEm\
        );

    \I__1358\ : IoInMux
    port map (
            O => \N__7099\,
            I => \N__7096\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__7096\,
            I => \N__7093\
        );

    \I__1356\ : Span4Mux_s1_h
    port map (
            O => \N__7093\,
            I => \N__7090\
        );

    \I__1355\ : Span4Mux_h
    port map (
            O => \N__7090\,
            I => \N__7087\
        );

    \I__1354\ : Sp12to4
    port map (
            O => \N__7087\,
            I => \N__7084\
        );

    \I__1353\ : Span12Mux_s10_v
    port map (
            O => \N__7084\,
            I => \N__7081\
        );

    \I__1352\ : Span12Mux_h
    port map (
            O => \N__7081\,
            I => \N__7078\
        );

    \I__1351\ : Odrv12
    port map (
            O => \N__7078\,
            I => \N_483\
        );

    \I__1350\ : IoInMux
    port map (
            O => \N__7075\,
            I => \N__7072\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__7072\,
            I => \N__7069\
        );

    \I__1348\ : Span12Mux_s8_v
    port map (
            O => \N__7069\,
            I => \N__7066\
        );

    \I__1347\ : Odrv12
    port map (
            O => \N__7066\,
            I => \CMA_c_10\
        );

    \I__1346\ : IoInMux
    port map (
            O => \N__7063\,
            I => \N__7060\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__7060\,
            I => \N__7057\
        );

    \I__1344\ : Odrv12
    port map (
            O => \N__7057\,
            I => \CMA_c_1\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7054\,
            I => \N__7051\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__7051\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i\
        );

    \I__1341\ : CascadeMux
    port map (
            O => \N__7048\,
            I => \U712_CYCLE_TERM.TACK_EN_RNOZ0Z_0_cascade_\
        );

    \I__1340\ : CascadeMux
    port map (
            O => \N__7045\,
            I => \U712_CYCLE_TERM.N_598_cascade_\
        );

    \I__1339\ : CascadeMux
    port map (
            O => \N__7042\,
            I => \N__7038\
        );

    \I__1338\ : InMux
    port map (
            O => \N__7041\,
            I => \N__7034\
        );

    \I__1337\ : InMux
    port map (
            O => \N__7038\,
            I => \N__7031\
        );

    \I__1336\ : InMux
    port map (
            O => \N__7037\,
            I => \N__7028\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__7034\,
            I => \N__7025\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__7031\,
            I => \N__7022\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__7028\,
            I => \U712_REG_SM.N_422\
        );

    \I__1332\ : Odrv4
    port map (
            O => \N__7025\,
            I => \U712_REG_SM.N_422\
        );

    \I__1331\ : Odrv12
    port map (
            O => \N__7022\,
            I => \U712_REG_SM.N_422\
        );

    \I__1330\ : InMux
    port map (
            O => \N__7015\,
            I => \N__7012\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__7012\,
            I => \N__7009\
        );

    \I__1328\ : Span4Mux_h
    port map (
            O => \N__7009\,
            I => \N__7006\
        );

    \I__1327\ : Odrv4
    port map (
            O => \N__7006\,
            I => \U712_REG_SM.N_514\
        );

    \I__1326\ : CascadeMux
    port map (
            O => \N__7003\,
            I => \N__6999\
        );

    \I__1325\ : InMux
    port map (
            O => \N__7002\,
            I => \N__6994\
        );

    \I__1324\ : InMux
    port map (
            O => \N__6999\,
            I => \N__6987\
        );

    \I__1323\ : InMux
    port map (
            O => \N__6998\,
            I => \N__6987\
        );

    \I__1322\ : InMux
    port map (
            O => \N__6997\,
            I => \N__6987\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__6994\,
            I => \REG_TACK\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__6987\,
            I => \REG_TACK\
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__6982\,
            I => \N__6979\
        );

    \I__1318\ : InMux
    port map (
            O => \N__6979\,
            I => \N__6973\
        );

    \I__1317\ : InMux
    port map (
            O => \N__6978\,
            I => \N__6966\
        );

    \I__1316\ : InMux
    port map (
            O => \N__6977\,
            I => \N__6966\
        );

    \I__1315\ : InMux
    port map (
            O => \N__6976\,
            I => \N__6966\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__6973\,
            I => \N__6963\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__6966\,
            I => \N__6960\
        );

    \I__1312\ : Span4Mux_h
    port map (
            O => \N__6963\,
            I => \N__6957\
        );

    \I__1311\ : Span4Mux_h
    port map (
            O => \N__6960\,
            I => \N__6954\
        );

    \I__1310\ : Odrv4
    port map (
            O => \N__6957\,
            I => \CPU_TACKm\
        );

    \I__1309\ : Odrv4
    port map (
            O => \N__6954\,
            I => \CPU_TACKm\
        );

    \I__1308\ : InMux
    port map (
            O => \N__6949\,
            I => \N__6941\
        );

    \I__1307\ : InMux
    port map (
            O => \N__6948\,
            I => \N__6941\
        );

    \I__1306\ : InMux
    port map (
            O => \N__6947\,
            I => \N__6936\
        );

    \I__1305\ : InMux
    port map (
            O => \N__6946\,
            I => \N__6936\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__6941\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__6936\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1302\ : CascadeMux
    port map (
            O => \N__6931\,
            I => \U712_CYCLE_TERM.N_571_cascade_\
        );

    \I__1301\ : InMux
    port map (
            O => \N__6928\,
            I => \N__6924\
        );

    \I__1300\ : InMux
    port map (
            O => \N__6927\,
            I => \N__6921\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__6924\,
            I => \U712_REG_SM.N_480\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__6921\,
            I => \U712_REG_SM.N_480\
        );

    \I__1297\ : InMux
    port map (
            O => \N__6916\,
            I => \N__6913\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__6913\,
            I => \U712_REG_SM.REG_TACK_RNOZ0Z_0\
        );

    \I__1295\ : InMux
    port map (
            O => \N__6910\,
            I => \N__6906\
        );

    \I__1294\ : InMux
    port map (
            O => \N__6909\,
            I => \N__6903\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__6906\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__6903\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1291\ : InMux
    port map (
            O => \N__6898\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__1290\ : InMux
    port map (
            O => \N__6895\,
            I => \N__6891\
        );

    \I__1289\ : InMux
    port map (
            O => \N__6894\,
            I => \N__6888\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__6891\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__6888\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1286\ : InMux
    port map (
            O => \N__6883\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__1285\ : InMux
    port map (
            O => \N__6880\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__1284\ : InMux
    port map (
            O => \N__6877\,
            I => \N__6873\
        );

    \I__1283\ : InMux
    port map (
            O => \N__6876\,
            I => \N__6870\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__6873\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__6870\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1280\ : ClkMux
    port map (
            O => \N__6865\,
            I => \N__6841\
        );

    \I__1279\ : ClkMux
    port map (
            O => \N__6864\,
            I => \N__6841\
        );

    \I__1278\ : ClkMux
    port map (
            O => \N__6863\,
            I => \N__6841\
        );

    \I__1277\ : ClkMux
    port map (
            O => \N__6862\,
            I => \N__6841\
        );

    \I__1276\ : ClkMux
    port map (
            O => \N__6861\,
            I => \N__6841\
        );

    \I__1275\ : ClkMux
    port map (
            O => \N__6860\,
            I => \N__6841\
        );

    \I__1274\ : ClkMux
    port map (
            O => \N__6859\,
            I => \N__6841\
        );

    \I__1273\ : ClkMux
    port map (
            O => \N__6858\,
            I => \N__6841\
        );

    \I__1272\ : GlobalMux
    port map (
            O => \N__6841\,
            I => \N__6838\
        );

    \I__1271\ : gio2CtrlBuf
    port map (
            O => \N__6838\,
            I => \C1_c_g\
        );

    \I__1270\ : InMux
    port map (
            O => \N__6835\,
            I => \N__6832\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__6832\,
            I => \N__6829\
        );

    \I__1268\ : Span4Mux_v
    port map (
            O => \N__6829\,
            I => \N__6826\
        );

    \I__1267\ : Sp12to4
    port map (
            O => \N__6826\,
            I => \N__6823\
        );

    \I__1266\ : Span12Mux_h
    port map (
            O => \N__6823\,
            I => \N__6820\
        );

    \I__1265\ : Span12Mux_v
    port map (
            O => \N__6820\,
            I => \N__6817\
        );

    \I__1264\ : Odrv12
    port map (
            O => \N__6817\,
            I => \A_c_2\
        );

    \I__1263\ : IoInMux
    port map (
            O => \N__6814\,
            I => \N__6810\
        );

    \I__1262\ : InMux
    port map (
            O => \N__6813\,
            I => \N__6807\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__6810\,
            I => \N__6804\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__6807\,
            I => \N__6801\
        );

    \I__1259\ : Span12Mux_s4_v
    port map (
            O => \N__6804\,
            I => \N__6798\
        );

    \I__1258\ : Span4Mux_h
    port map (
            O => \N__6801\,
            I => \N__6795\
        );

    \I__1257\ : Span12Mux_v
    port map (
            O => \N__6798\,
            I => \N__6792\
        );

    \I__1256\ : Span4Mux_v
    port map (
            O => \N__6795\,
            I => \N__6789\
        );

    \I__1255\ : Span12Mux_h
    port map (
            O => \N__6792\,
            I => \N__6786\
        );

    \I__1254\ : Sp12to4
    port map (
            O => \N__6789\,
            I => \N__6783\
        );

    \I__1253\ : Odrv12
    port map (
            O => \N__6786\,
            I => \A_c_9\
        );

    \I__1252\ : Odrv12
    port map (
            O => \N__6783\,
            I => \A_c_9\
        );

    \I__1251\ : SRMux
    port map (
            O => \N__6778\,
            I => \N__6775\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__6775\,
            I => \N__6772\
        );

    \I__1249\ : Span4Mux_h
    port map (
            O => \N__6772\,
            I => \N__6769\
        );

    \I__1248\ : Odrv4
    port map (
            O => \N__6769\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__1247\ : CascadeMux
    port map (
            O => \N__6766\,
            I => \U712_CHIP_RAM.REFRESH_RST_cascade_\
        );

    \I__1246\ : InMux
    port map (
            O => \N__6763\,
            I => \N__6756\
        );

    \I__1245\ : InMux
    port map (
            O => \N__6762\,
            I => \N__6753\
        );

    \I__1244\ : CascadeMux
    port map (
            O => \N__6761\,
            I => \N__6748\
        );

    \I__1243\ : InMux
    port map (
            O => \N__6760\,
            I => \N__6744\
        );

    \I__1242\ : InMux
    port map (
            O => \N__6759\,
            I => \N__6741\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__6756\,
            I => \N__6731\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__6753\,
            I => \N__6731\
        );

    \I__1239\ : InMux
    port map (
            O => \N__6752\,
            I => \N__6728\
        );

    \I__1238\ : InMux
    port map (
            O => \N__6751\,
            I => \N__6721\
        );

    \I__1237\ : InMux
    port map (
            O => \N__6748\,
            I => \N__6721\
        );

    \I__1236\ : InMux
    port map (
            O => \N__6747\,
            I => \N__6721\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__6744\,
            I => \N__6718\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__6741\,
            I => \N__6715\
        );

    \I__1233\ : InMux
    port map (
            O => \N__6740\,
            I => \N__6710\
        );

    \I__1232\ : InMux
    port map (
            O => \N__6739\,
            I => \N__6710\
        );

    \I__1231\ : InMux
    port map (
            O => \N__6738\,
            I => \N__6707\
        );

    \I__1230\ : InMux
    port map (
            O => \N__6737\,
            I => \N__6704\
        );

    \I__1229\ : InMux
    port map (
            O => \N__6736\,
            I => \N__6701\
        );

    \I__1228\ : Span4Mux_h
    port map (
            O => \N__6731\,
            I => \N__6694\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__6728\,
            I => \N__6694\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__6721\,
            I => \N__6694\
        );

    \I__1225\ : Span4Mux_v
    port map (
            O => \N__6718\,
            I => \N__6689\
        );

    \I__1224\ : Span4Mux_v
    port map (
            O => \N__6715\,
            I => \N__6689\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__6710\,
            I => \N__6686\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__6707\,
            I => \N__6681\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__6704\,
            I => \N__6681\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__6701\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1219\ : Odrv4
    port map (
            O => \N__6694\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1218\ : Odrv4
    port map (
            O => \N__6689\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1217\ : Odrv4
    port map (
            O => \N__6686\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1216\ : Odrv12
    port map (
            O => \N__6681\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__6670\,
            I => \N__6666\
        );

    \I__1214\ : InMux
    port map (
            O => \N__6669\,
            I => \N__6662\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6666\,
            I => \N__6658\
        );

    \I__1212\ : InMux
    port map (
            O => \N__6665\,
            I => \N__6655\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__6662\,
            I => \N__6648\
        );

    \I__1210\ : InMux
    port map (
            O => \N__6661\,
            I => \N__6645\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__6658\,
            I => \N__6642\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__6655\,
            I => \N__6639\
        );

    \I__1207\ : InMux
    port map (
            O => \N__6654\,
            I => \N__6636\
        );

    \I__1206\ : InMux
    port map (
            O => \N__6653\,
            I => \N__6633\
        );

    \I__1205\ : InMux
    port map (
            O => \N__6652\,
            I => \N__6628\
        );

    \I__1204\ : InMux
    port map (
            O => \N__6651\,
            I => \N__6628\
        );

    \I__1203\ : Odrv4
    port map (
            O => \N__6648\,
            I => \U712_CHIP_RAM.N_595\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__6645\,
            I => \U712_CHIP_RAM.N_595\
        );

    \I__1201\ : Odrv4
    port map (
            O => \N__6642\,
            I => \U712_CHIP_RAM.N_595\
        );

    \I__1200\ : Odrv4
    port map (
            O => \N__6639\,
            I => \U712_CHIP_RAM.N_595\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__6636\,
            I => \U712_CHIP_RAM.N_595\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__6633\,
            I => \U712_CHIP_RAM.N_595\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__6628\,
            I => \U712_CHIP_RAM.N_595\
        );

    \I__1196\ : CEMux
    port map (
            O => \N__6613\,
            I => \N__6610\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__6610\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0\
        );

    \I__1194\ : InMux
    port map (
            O => \N__6607\,
            I => \N__6604\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__6604\,
            I => \U712_REG_SM.N_443\
        );

    \I__1192\ : CascadeMux
    port map (
            O => \N__6601\,
            I => \N__6597\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6600\,
            I => \N__6588\
        );

    \I__1190\ : InMux
    port map (
            O => \N__6597\,
            I => \N__6588\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6596\,
            I => \N__6581\
        );

    \I__1188\ : InMux
    port map (
            O => \N__6595\,
            I => \N__6581\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6594\,
            I => \N__6581\
        );

    \I__1186\ : CascadeMux
    port map (
            O => \N__6593\,
            I => \N__6574\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__6588\,
            I => \N__6568\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__6581\,
            I => \N__6568\
        );

    \I__1183\ : InMux
    port map (
            O => \N__6580\,
            I => \N__6565\
        );

    \I__1182\ : InMux
    port map (
            O => \N__6579\,
            I => \N__6562\
        );

    \I__1181\ : InMux
    port map (
            O => \N__6578\,
            I => \N__6559\
        );

    \I__1180\ : InMux
    port map (
            O => \N__6577\,
            I => \N__6552\
        );

    \I__1179\ : InMux
    port map (
            O => \N__6574\,
            I => \N__6552\
        );

    \I__1178\ : InMux
    port map (
            O => \N__6573\,
            I => \N__6552\
        );

    \I__1177\ : Span4Mux_v
    port map (
            O => \N__6568\,
            I => \N__6549\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__6565\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6562\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__6559\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__6552\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1172\ : Odrv4
    port map (
            O => \N__6549\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1171\ : InMux
    port map (
            O => \N__6538\,
            I => \N__6531\
        );

    \I__1170\ : InMux
    port map (
            O => \N__6537\,
            I => \N__6522\
        );

    \I__1169\ : InMux
    port map (
            O => \N__6536\,
            I => \N__6522\
        );

    \I__1168\ : InMux
    port map (
            O => \N__6535\,
            I => \N__6522\
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__6534\,
            I => \N__6519\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__6531\,
            I => \N__6516\
        );

    \I__1165\ : CascadeMux
    port map (
            O => \N__6530\,
            I => \N__6513\
        );

    \I__1164\ : CascadeMux
    port map (
            O => \N__6529\,
            I => \N__6509\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__6522\,
            I => \N__6502\
        );

    \I__1162\ : InMux
    port map (
            O => \N__6519\,
            I => \N__6499\
        );

    \I__1161\ : Span4Mux_v
    port map (
            O => \N__6516\,
            I => \N__6496\
        );

    \I__1160\ : InMux
    port map (
            O => \N__6513\,
            I => \N__6493\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6512\,
            I => \N__6490\
        );

    \I__1158\ : InMux
    port map (
            O => \N__6509\,
            I => \N__6479\
        );

    \I__1157\ : InMux
    port map (
            O => \N__6508\,
            I => \N__6479\
        );

    \I__1156\ : InMux
    port map (
            O => \N__6507\,
            I => \N__6479\
        );

    \I__1155\ : InMux
    port map (
            O => \N__6506\,
            I => \N__6479\
        );

    \I__1154\ : InMux
    port map (
            O => \N__6505\,
            I => \N__6479\
        );

    \I__1153\ : Span4Mux_v
    port map (
            O => \N__6502\,
            I => \N__6476\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__6499\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1151\ : Odrv4
    port map (
            O => \N__6496\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__6493\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__6490\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__6479\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1147\ : Odrv4
    port map (
            O => \N__6476\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1146\ : IoInMux
    port map (
            O => \N__6463\,
            I => \N__6459\
        );

    \I__1145\ : IoInMux
    port map (
            O => \N__6462\,
            I => \N__6456\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__6459\,
            I => \N__6453\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__6456\,
            I => \N__6450\
        );

    \I__1142\ : Span4Mux_s3_v
    port map (
            O => \N__6453\,
            I => \N__6447\
        );

    \I__1141\ : Span4Mux_s3_v
    port map (
            O => \N__6450\,
            I => \N__6444\
        );

    \I__1140\ : Sp12to4
    port map (
            O => \N__6447\,
            I => \N__6441\
        );

    \I__1139\ : Sp12to4
    port map (
            O => \N__6444\,
            I => \N__6438\
        );

    \I__1138\ : Span12Mux_s9_h
    port map (
            O => \N__6441\,
            I => \N__6435\
        );

    \I__1137\ : Span12Mux_s10_h
    port map (
            O => \N__6438\,
            I => \N__6432\
        );

    \I__1136\ : Span12Mux_v
    port map (
            O => \N__6435\,
            I => \N__6426\
        );

    \I__1135\ : Span12Mux_v
    port map (
            O => \N__6432\,
            I => \N__6426\
        );

    \I__1134\ : InMux
    port map (
            O => \N__6431\,
            I => \N__6423\
        );

    \I__1133\ : Odrv12
    port map (
            O => \N__6426\,
            I => \ASn_c\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__6423\,
            I => \ASn_c\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6418\,
            I => \N__6412\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6417\,
            I => \N__6412\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6412\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1128\ : IoInMux
    port map (
            O => \N__6409\,
            I => \N__6406\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__6406\,
            I => \N__6403\
        );

    \I__1126\ : Span4Mux_s3_v
    port map (
            O => \N__6403\,
            I => \N__6400\
        );

    \I__1125\ : Span4Mux_v
    port map (
            O => \N__6400\,
            I => \N__6397\
        );

    \I__1124\ : Span4Mux_v
    port map (
            O => \N__6397\,
            I => \N__6394\
        );

    \I__1123\ : Odrv4
    port map (
            O => \N__6394\,
            I => \RESETn_c_i\
        );

    \I__1122\ : IoInMux
    port map (
            O => \N__6391\,
            I => \N__6388\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__6388\,
            I => \N__6385\
        );

    \I__1120\ : Span4Mux_s3_v
    port map (
            O => \N__6385\,
            I => \N__6382\
        );

    \I__1119\ : Span4Mux_h
    port map (
            O => \N__6382\,
            I => \N__6379\
        );

    \I__1118\ : Span4Mux_v
    port map (
            O => \N__6379\,
            I => \N__6376\
        );

    \I__1117\ : Odrv4
    port map (
            O => \N__6376\,
            I => \N_549\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6373\,
            I => \N__6369\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6372\,
            I => \N__6366\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__6369\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__6366\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__1112\ : InMux
    port map (
            O => \N__6361\,
            I => \bfn_11_5_0_\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6358\,
            I => \N__6354\
        );

    \I__1110\ : InMux
    port map (
            O => \N__6357\,
            I => \N__6351\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__6354\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__6351\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6346\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__1106\ : InMux
    port map (
            O => \N__6343\,
            I => \N__6339\
        );

    \I__1105\ : InMux
    port map (
            O => \N__6342\,
            I => \N__6336\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__6339\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__6336\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__1102\ : InMux
    port map (
            O => \N__6331\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__1101\ : InMux
    port map (
            O => \N__6328\,
            I => \N__6324\
        );

    \I__1100\ : InMux
    port map (
            O => \N__6327\,
            I => \N__6321\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__6324\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__6321\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1097\ : InMux
    port map (
            O => \N__6316\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__1096\ : CascadeMux
    port map (
            O => \N__6313\,
            I => \N__6309\
        );

    \I__1095\ : InMux
    port map (
            O => \N__6312\,
            I => \N__6306\
        );

    \I__1094\ : InMux
    port map (
            O => \N__6309\,
            I => \N__6303\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__6306\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__6303\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1091\ : InMux
    port map (
            O => \N__6298\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__1090\ : InMux
    port map (
            O => \N__6295\,
            I => \N__6292\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__6292\,
            I => \U712_REG_SM.STATE_COUNT_srsts_i_i_i_a2_0_0_0\
        );

    \I__1088\ : InMux
    port map (
            O => \N__6289\,
            I => \N__6283\
        );

    \I__1087\ : InMux
    port map (
            O => \N__6288\,
            I => \N__6276\
        );

    \I__1086\ : InMux
    port map (
            O => \N__6287\,
            I => \N__6276\
        );

    \I__1085\ : InMux
    port map (
            O => \N__6286\,
            I => \N__6276\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__6283\,
            I => \N__6269\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__6276\,
            I => \N__6269\
        );

    \I__1082\ : InMux
    port map (
            O => \N__6275\,
            I => \N__6264\
        );

    \I__1081\ : InMux
    port map (
            O => \N__6274\,
            I => \N__6264\
        );

    \I__1080\ : Odrv12
    port map (
            O => \N__6269\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__6264\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1078\ : InMux
    port map (
            O => \N__6259\,
            I => \N__6256\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__6256\,
            I => \N__6249\
        );

    \I__1076\ : InMux
    port map (
            O => \N__6255\,
            I => \N__6242\
        );

    \I__1075\ : InMux
    port map (
            O => \N__6254\,
            I => \N__6242\
        );

    \I__1074\ : InMux
    port map (
            O => \N__6253\,
            I => \N__6242\
        );

    \I__1073\ : InMux
    port map (
            O => \N__6252\,
            I => \N__6237\
        );

    \I__1072\ : Sp12to4
    port map (
            O => \N__6249\,
            I => \N__6232\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__6242\,
            I => \N__6232\
        );

    \I__1070\ : InMux
    port map (
            O => \N__6241\,
            I => \N__6227\
        );

    \I__1069\ : InMux
    port map (
            O => \N__6240\,
            I => \N__6227\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__6237\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1067\ : Odrv12
    port map (
            O => \N__6232\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__6227\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1065\ : InMux
    port map (
            O => \N__6220\,
            I => \N__6213\
        );

    \I__1064\ : InMux
    port map (
            O => \N__6219\,
            I => \N__6213\
        );

    \I__1063\ : InMux
    port map (
            O => \N__6218\,
            I => \N__6210\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__6213\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__6210\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1060\ : InMux
    port map (
            O => \N__6205\,
            I => \N__6202\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__6202\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_0\
        );

    \I__1058\ : InMux
    port map (
            O => \N__6199\,
            I => \N__6196\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__6196\,
            I => \N__6192\
        );

    \I__1056\ : InMux
    port map (
            O => \N__6195\,
            I => \N__6189\
        );

    \I__1055\ : Odrv12
    port map (
            O => \N__6192\,
            I => \U712_REG_SM.START_RST_0_sqmuxa\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__6189\,
            I => \U712_REG_SM.START_RST_0_sqmuxa\
        );

    \I__1053\ : InMux
    port map (
            O => \N__6184\,
            I => \N__6181\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__6181\,
            I => \U712_REG_SM.un1_STATE_COUNT_4_i_i_0_0\
        );

    \I__1051\ : InMux
    port map (
            O => \N__6178\,
            I => \N__6175\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__6175\,
            I => \U712_REG_SM.DS_EN_RNOZ0Z_0\
        );

    \I__1049\ : CascadeMux
    port map (
            O => \N__6172\,
            I => \N__6169\
        );

    \I__1048\ : InMux
    port map (
            O => \N__6169\,
            I => \N__6166\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__6166\,
            I => \N__6163\
        );

    \I__1046\ : Odrv4
    port map (
            O => \N__6163\,
            I => \U712_REG_SM.N_515\
        );

    \I__1045\ : InMux
    port map (
            O => \N__6160\,
            I => \N__6157\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__6157\,
            I => \N__6154\
        );

    \I__1043\ : Odrv4
    port map (
            O => \N__6154\,
            I => \U712_CHIP_RAM.N_537\
        );

    \I__1042\ : InMux
    port map (
            O => \N__6151\,
            I => \N__6147\
        );

    \I__1041\ : InMux
    port map (
            O => \N__6150\,
            I => \N__6142\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__6147\,
            I => \N__6139\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6146\,
            I => \N__6136\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6145\,
            I => \N__6133\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__6142\,
            I => \N__6130\
        );

    \I__1036\ : Span4Mux_v
    port map (
            O => \N__6139\,
            I => \N__6125\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__6136\,
            I => \N__6125\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__6133\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__1033\ : Odrv4
    port map (
            O => \N__6130\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__1032\ : Odrv4
    port map (
            O => \N__6125\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__1031\ : InMux
    port map (
            O => \N__6118\,
            I => \N__6115\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__6115\,
            I => \N__6112\
        );

    \I__1029\ : Odrv4
    port map (
            O => \N__6112\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_0_0\
        );

    \I__1028\ : InMux
    port map (
            O => \N__6109\,
            I => \N__6098\
        );

    \I__1027\ : InMux
    port map (
            O => \N__6108\,
            I => \N__6098\
        );

    \I__1026\ : CascadeMux
    port map (
            O => \N__6107\,
            I => \N__6094\
        );

    \I__1025\ : CascadeMux
    port map (
            O => \N__6106\,
            I => \N__6090\
        );

    \I__1024\ : InMux
    port map (
            O => \N__6105\,
            I => \N__6083\
        );

    \I__1023\ : InMux
    port map (
            O => \N__6104\,
            I => \N__6077\
        );

    \I__1022\ : InMux
    port map (
            O => \N__6103\,
            I => \N__6077\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__6098\,
            I => \N__6074\
        );

    \I__1020\ : InMux
    port map (
            O => \N__6097\,
            I => \N__6071\
        );

    \I__1019\ : InMux
    port map (
            O => \N__6094\,
            I => \N__6068\
        );

    \I__1018\ : InMux
    port map (
            O => \N__6093\,
            I => \N__6063\
        );

    \I__1017\ : InMux
    port map (
            O => \N__6090\,
            I => \N__6063\
        );

    \I__1016\ : InMux
    port map (
            O => \N__6089\,
            I => \N__6056\
        );

    \I__1015\ : InMux
    port map (
            O => \N__6088\,
            I => \N__6056\
        );

    \I__1014\ : CascadeMux
    port map (
            O => \N__6087\,
            I => \N__6053\
        );

    \I__1013\ : CascadeMux
    port map (
            O => \N__6086\,
            I => \N__6049\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__6083\,
            I => \N__6045\
        );

    \I__1011\ : InMux
    port map (
            O => \N__6082\,
            I => \N__6042\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__6077\,
            I => \N__6039\
        );

    \I__1009\ : Span4Mux_v
    port map (
            O => \N__6074\,
            I => \N__6032\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__6071\,
            I => \N__6032\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__6068\,
            I => \N__6032\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__6063\,
            I => \N__6029\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6062\,
            I => \N__6026\
        );

    \I__1004\ : InMux
    port map (
            O => \N__6061\,
            I => \N__6023\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__6056\,
            I => \N__6020\
        );

    \I__1002\ : InMux
    port map (
            O => \N__6053\,
            I => \N__6017\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6052\,
            I => \N__6014\
        );

    \I__1000\ : InMux
    port map (
            O => \N__6049\,
            I => \N__6009\
        );

    \I__999\ : InMux
    port map (
            O => \N__6048\,
            I => \N__6009\
        );

    \I__998\ : Span4Mux_v
    port map (
            O => \N__6045\,
            I => \N__5998\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__6042\,
            I => \N__5998\
        );

    \I__996\ : Span4Mux_v
    port map (
            O => \N__6039\,
            I => \N__5998\
        );

    \I__995\ : Span4Mux_h
    port map (
            O => \N__6032\,
            I => \N__5998\
        );

    \I__994\ : Span4Mux_v
    port map (
            O => \N__6029\,
            I => \N__5998\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__6026\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__6023\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__991\ : Odrv4
    port map (
            O => \N__6020\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__6017\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__6014\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__6009\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__987\ : Odrv4
    port map (
            O => \N__5998\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__986\ : CascadeMux
    port map (
            O => \N__5983\,
            I => \N__5979\
        );

    \I__985\ : InMux
    port map (
            O => \N__5982\,
            I => \N__5972\
        );

    \I__984\ : InMux
    port map (
            O => \N__5979\,
            I => \N__5969\
        );

    \I__983\ : InMux
    port map (
            O => \N__5978\,
            I => \N__5965\
        );

    \I__982\ : CascadeMux
    port map (
            O => \N__5977\,
            I => \N__5959\
        );

    \I__981\ : CascadeMux
    port map (
            O => \N__5976\,
            I => \N__5955\
        );

    \I__980\ : CascadeMux
    port map (
            O => \N__5975\,
            I => \N__5949\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__5972\,
            I => \N__5943\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__5969\,
            I => \N__5943\
        );

    \I__977\ : InMux
    port map (
            O => \N__5968\,
            I => \N__5938\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__5965\,
            I => \N__5935\
        );

    \I__975\ : InMux
    port map (
            O => \N__5964\,
            I => \N__5928\
        );

    \I__974\ : InMux
    port map (
            O => \N__5963\,
            I => \N__5928\
        );

    \I__973\ : InMux
    port map (
            O => \N__5962\,
            I => \N__5928\
        );

    \I__972\ : InMux
    port map (
            O => \N__5959\,
            I => \N__5922\
        );

    \I__971\ : InMux
    port map (
            O => \N__5958\,
            I => \N__5915\
        );

    \I__970\ : InMux
    port map (
            O => \N__5955\,
            I => \N__5915\
        );

    \I__969\ : InMux
    port map (
            O => \N__5954\,
            I => \N__5915\
        );

    \I__968\ : InMux
    port map (
            O => \N__5953\,
            I => \N__5912\
        );

    \I__967\ : InMux
    port map (
            O => \N__5952\,
            I => \N__5909\
        );

    \I__966\ : InMux
    port map (
            O => \N__5949\,
            I => \N__5906\
        );

    \I__965\ : InMux
    port map (
            O => \N__5948\,
            I => \N__5903\
        );

    \I__964\ : Span12Mux_h
    port map (
            O => \N__5943\,
            I => \N__5900\
        );

    \I__963\ : InMux
    port map (
            O => \N__5942\,
            I => \N__5895\
        );

    \I__962\ : InMux
    port map (
            O => \N__5941\,
            I => \N__5895\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__5938\,
            I => \N__5890\
        );

    \I__960\ : Span4Mux_h
    port map (
            O => \N__5935\,
            I => \N__5890\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__5928\,
            I => \N__5887\
        );

    \I__958\ : InMux
    port map (
            O => \N__5927\,
            I => \N__5884\
        );

    \I__957\ : InMux
    port map (
            O => \N__5926\,
            I => \N__5879\
        );

    \I__956\ : InMux
    port map (
            O => \N__5925\,
            I => \N__5879\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__5922\,
            I => \N__5874\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__5915\,
            I => \N__5874\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__5912\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__5909\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__5906\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__5903\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__949\ : Odrv12
    port map (
            O => \N__5900\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__5895\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__947\ : Odrv4
    port map (
            O => \N__5890\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__946\ : Odrv4
    port map (
            O => \N__5887\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__5884\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__5879\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__943\ : Odrv12
    port map (
            O => \N__5874\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__942\ : InMux
    port map (
            O => \N__5851\,
            I => \N__5847\
        );

    \I__941\ : InMux
    port map (
            O => \N__5850\,
            I => \N__5844\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__5847\,
            I => \U712_CHIP_RAM.N_703\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__5844\,
            I => \U712_CHIP_RAM.N_703\
        );

    \I__938\ : CascadeMux
    port map (
            O => \N__5839\,
            I => \U712_CHIP_RAM.N_530_cascade_\
        );

    \I__937\ : InMux
    port map (
            O => \N__5836\,
            I => \N__5831\
        );

    \I__936\ : InMux
    port map (
            O => \N__5835\,
            I => \N__5826\
        );

    \I__935\ : InMux
    port map (
            O => \N__5834\,
            I => \N__5823\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__5831\,
            I => \N__5820\
        );

    \I__933\ : InMux
    port map (
            O => \N__5830\,
            I => \N__5817\
        );

    \I__932\ : InMux
    port map (
            O => \N__5829\,
            I => \N__5814\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__5826\,
            I => \N__5809\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__5823\,
            I => \N__5809\
        );

    \I__929\ : Odrv4
    port map (
            O => \N__5820\,
            I => \U712_CHIP_RAM.N_600\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__5817\,
            I => \U712_CHIP_RAM.N_600\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__5814\,
            I => \U712_CHIP_RAM.N_600\
        );

    \I__926\ : Odrv4
    port map (
            O => \N__5809\,
            I => \U712_CHIP_RAM.N_600\
        );

    \I__925\ : CascadeMux
    port map (
            O => \N__5800\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_cascade_\
        );

    \I__924\ : CEMux
    port map (
            O => \N__5797\,
            I => \N__5794\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__5794\,
            I => \N__5791\
        );

    \I__922\ : Span4Mux_h
    port map (
            O => \N__5791\,
            I => \N__5788\
        );

    \I__921\ : Odrv4
    port map (
            O => \N__5788\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0\
        );

    \I__920\ : InMux
    port map (
            O => \N__5785\,
            I => \N__5781\
        );

    \I__919\ : InMux
    port map (
            O => \N__5784\,
            I => \N__5778\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__5781\,
            I => \N__5775\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__5778\,
            I => \N__5772\
        );

    \I__916\ : Span4Mux_v
    port map (
            O => \N__5775\,
            I => \N__5769\
        );

    \I__915\ : Span4Mux_v
    port map (
            O => \N__5772\,
            I => \N__5766\
        );

    \I__914\ : Sp12to4
    port map (
            O => \N__5769\,
            I => \N__5763\
        );

    \I__913\ : Span4Mux_h
    port map (
            O => \N__5766\,
            I => \N__5760\
        );

    \I__912\ : Span12Mux_h
    port map (
            O => \N__5763\,
            I => \N__5755\
        );

    \I__911\ : Sp12to4
    port map (
            O => \N__5760\,
            I => \N__5755\
        );

    \I__910\ : Span12Mux_v
    port map (
            O => \N__5755\,
            I => \N__5752\
        );

    \I__909\ : Odrv12
    port map (
            O => \N__5752\,
            I => \AWEn_c\
        );

    \I__908\ : InMux
    port map (
            O => \N__5749\,
            I => \N__5746\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__5746\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\
        );

    \I__906\ : IoInMux
    port map (
            O => \N__5743\,
            I => \N__5740\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__5740\,
            I => \N__5737\
        );

    \I__904\ : IoSpan4Mux
    port map (
            O => \N__5737\,
            I => \N__5734\
        );

    \I__903\ : Span4Mux_s2_v
    port map (
            O => \N__5734\,
            I => \N__5731\
        );

    \I__902\ : Sp12to4
    port map (
            O => \N__5731\,
            I => \N__5727\
        );

    \I__901\ : InMux
    port map (
            O => \N__5730\,
            I => \N__5724\
        );

    \I__900\ : Odrv12
    port map (
            O => \N__5727\,
            I => \DBDIR_c\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__5724\,
            I => \DBDIR_c\
        );

    \I__898\ : InMux
    port map (
            O => \N__5719\,
            I => \N__5716\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__5716\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0\
        );

    \I__896\ : InMux
    port map (
            O => \N__5713\,
            I => \N__5710\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__5710\,
            I => \U712_CHIP_RAM.DBENn_8_0\
        );

    \I__894\ : InMux
    port map (
            O => \N__5707\,
            I => \N__5703\
        );

    \I__893\ : InMux
    port map (
            O => \N__5706\,
            I => \N__5700\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__5703\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__5700\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__890\ : CascadeMux
    port map (
            O => \N__5695\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_\
        );

    \I__889\ : IoInMux
    port map (
            O => \N__5692\,
            I => \N__5689\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__5689\,
            I => \N__5686\
        );

    \I__887\ : Span4Mux_s3_v
    port map (
            O => \N__5686\,
            I => \N__5683\
        );

    \I__886\ : Sp12to4
    port map (
            O => \N__5683\,
            I => \N__5680\
        );

    \I__885\ : Span12Mux_h
    port map (
            O => \N__5680\,
            I => \N__5677\
        );

    \I__884\ : Span12Mux_v
    port map (
            O => \N__5677\,
            I => \N__5673\
        );

    \I__883\ : InMux
    port map (
            O => \N__5676\,
            I => \N__5670\
        );

    \I__882\ : Odrv12
    port map (
            O => \N__5673\,
            I => \LATCH_CLK_c\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__5670\,
            I => \LATCH_CLK_c\
        );

    \I__880\ : CascadeMux
    port map (
            O => \N__5665\,
            I => \N__5661\
        );

    \I__879\ : InMux
    port map (
            O => \N__5664\,
            I => \N__5658\
        );

    \I__878\ : InMux
    port map (
            O => \N__5661\,
            I => \N__5655\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__5658\,
            I => \U712_CHIP_RAM.N_528\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__5655\,
            I => \U712_CHIP_RAM.N_528\
        );

    \I__875\ : InMux
    port map (
            O => \N__5650\,
            I => \N__5647\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__5647\,
            I => \N__5641\
        );

    \I__873\ : InMux
    port map (
            O => \N__5646\,
            I => \N__5638\
        );

    \I__872\ : InMux
    port map (
            O => \N__5645\,
            I => \N__5633\
        );

    \I__871\ : InMux
    port map (
            O => \N__5644\,
            I => \N__5633\
        );

    \I__870\ : Span4Mux_h
    port map (
            O => \N__5641\,
            I => \N__5630\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__5638\,
            I => \N__5625\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__5633\,
            I => \N__5625\
        );

    \I__867\ : Odrv4
    port map (
            O => \N__5630\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__866\ : Odrv12
    port map (
            O => \N__5625\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__865\ : CascadeMux
    port map (
            O => \N__5620\,
            I => \U712_REG_SM.N_482_cascade_\
        );

    \I__864\ : InMux
    port map (
            O => \N__5617\,
            I => \N__5614\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__5614\,
            I => \N__5611\
        );

    \I__862\ : Span4Mux_v
    port map (
            O => \N__5611\,
            I => \N__5608\
        );

    \I__861\ : Span4Mux_h
    port map (
            O => \N__5608\,
            I => \N__5604\
        );

    \I__860\ : IoInMux
    port map (
            O => \N__5607\,
            I => \N__5601\
        );

    \I__859\ : Sp12to4
    port map (
            O => \N__5604\,
            I => \N__5598\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5601\,
            I => \N__5595\
        );

    \I__857\ : Span12Mux_v
    port map (
            O => \N__5598\,
            I => \N__5592\
        );

    \I__856\ : IoSpan4Mux
    port map (
            O => \N__5595\,
            I => \N__5589\
        );

    \I__855\ : Odrv12
    port map (
            O => \N__5592\,
            I => \RAMENn_c\
        );

    \I__854\ : Odrv4
    port map (
            O => \N__5589\,
            I => \RAMENn_c\
        );

    \I__853\ : CascadeMux
    port map (
            O => \N__5584\,
            I => \N__5581\
        );

    \I__852\ : InMux
    port map (
            O => \N__5581\,
            I => \N__5578\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__5578\,
            I => \N__5575\
        );

    \I__850\ : Odrv4
    port map (
            O => \N__5575\,
            I => \U712_CHIP_RAM.N_527\
        );

    \I__849\ : InMux
    port map (
            O => \N__5572\,
            I => \N__5569\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__5569\,
            I => \N__5566\
        );

    \I__847\ : Span4Mux_v
    port map (
            O => \N__5566\,
            I => \N__5562\
        );

    \I__846\ : InMux
    port map (
            O => \N__5565\,
            I => \N__5559\
        );

    \I__845\ : Sp12to4
    port map (
            O => \N__5562\,
            I => \N__5554\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__5559\,
            I => \N__5554\
        );

    \I__843\ : Span12Mux_h
    port map (
            O => \N__5554\,
            I => \N__5551\
        );

    \I__842\ : Span12Mux_v
    port map (
            O => \N__5551\,
            I => \N__5548\
        );

    \I__841\ : Odrv12
    port map (
            O => \N__5548\,
            I => \TSn_c\
        );

    \I__840\ : InMux
    port map (
            O => \N__5545\,
            I => \N__5542\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__5542\,
            I => \N__5537\
        );

    \I__838\ : InMux
    port map (
            O => \N__5541\,
            I => \N__5534\
        );

    \I__837\ : InMux
    port map (
            O => \N__5540\,
            I => \N__5531\
        );

    \I__836\ : Odrv4
    port map (
            O => \N__5537\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__5534\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__5531\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__833\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5520\
        );

    \I__832\ : InMux
    port map (
            O => \N__5523\,
            I => \N__5517\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__5520\,
            I => \N__5514\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__5517\,
            I => \U712_CHIP_RAM.N_553\
        );

    \I__829\ : Odrv12
    port map (
            O => \N__5514\,
            I => \U712_CHIP_RAM.N_553\
        );

    \I__828\ : CascadeMux
    port map (
            O => \N__5509\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1_cascade_\
        );

    \I__827\ : InMux
    port map (
            O => \N__5506\,
            I => \N__5503\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__5503\,
            I => \U712_CHIP_RAM.N_597\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__5500\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_cascade_\
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__5497\,
            I => \U712_REG_SM.N_429_cascade_\
        );

    \I__823\ : CascadeMux
    port map (
            O => \N__5494\,
            I => \U712_REG_SM.N_511_cascade_\
        );

    \I__822\ : InMux
    port map (
            O => \N__5491\,
            I => \N__5488\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__5488\,
            I => \N__5485\
        );

    \I__820\ : Span4Mux_h
    port map (
            O => \N__5485\,
            I => \N__5482\
        );

    \I__819\ : Odrv4
    port map (
            O => \N__5482\,
            I => \U712_REG_SM.N_694\
        );

    \I__818\ : InMux
    port map (
            O => \N__5479\,
            I => \N__5476\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__5476\,
            I => \N__5473\
        );

    \I__816\ : Span4Mux_h
    port map (
            O => \N__5473\,
            I => \N__5470\
        );

    \I__815\ : Odrv4
    port map (
            O => \N__5470\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_0\
        );

    \I__814\ : InMux
    port map (
            O => \N__5467\,
            I => \N__5463\
        );

    \I__813\ : InMux
    port map (
            O => \N__5466\,
            I => \N__5460\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5463\,
            I => \U712_CHIP_RAM.N_700\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__5460\,
            I => \U712_CHIP_RAM.N_700\
        );

    \I__810\ : InMux
    port map (
            O => \N__5455\,
            I => \N__5452\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__5452\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_0_a2_0_1\
        );

    \I__808\ : InMux
    port map (
            O => \N__5449\,
            I => \N__5442\
        );

    \I__807\ : CascadeMux
    port map (
            O => \N__5448\,
            I => \N__5439\
        );

    \I__806\ : CascadeMux
    port map (
            O => \N__5447\,
            I => \N__5436\
        );

    \I__805\ : InMux
    port map (
            O => \N__5446\,
            I => \N__5433\
        );

    \I__804\ : CascadeMux
    port map (
            O => \N__5445\,
            I => \N__5427\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__5442\,
            I => \N__5423\
        );

    \I__802\ : InMux
    port map (
            O => \N__5439\,
            I => \N__5420\
        );

    \I__801\ : InMux
    port map (
            O => \N__5436\,
            I => \N__5417\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__5433\,
            I => \N__5414\
        );

    \I__799\ : InMux
    port map (
            O => \N__5432\,
            I => \N__5411\
        );

    \I__798\ : InMux
    port map (
            O => \N__5431\,
            I => \N__5408\
        );

    \I__797\ : InMux
    port map (
            O => \N__5430\,
            I => \N__5405\
        );

    \I__796\ : InMux
    port map (
            O => \N__5427\,
            I => \N__5399\
        );

    \I__795\ : InMux
    port map (
            O => \N__5426\,
            I => \N__5396\
        );

    \I__794\ : Span4Mux_v
    port map (
            O => \N__5423\,
            I => \N__5393\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__5420\,
            I => \N__5386\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__5417\,
            I => \N__5386\
        );

    \I__791\ : Span4Mux_v
    port map (
            O => \N__5414\,
            I => \N__5386\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__5411\,
            I => \N__5379\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__5408\,
            I => \N__5379\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__5405\,
            I => \N__5379\
        );

    \I__787\ : InMux
    port map (
            O => \N__5404\,
            I => \N__5376\
        );

    \I__786\ : InMux
    port map (
            O => \N__5403\,
            I => \N__5373\
        );

    \I__785\ : InMux
    port map (
            O => \N__5402\,
            I => \N__5370\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__5399\,
            I => \U712_CHIP_RAM.N_578\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__5396\,
            I => \U712_CHIP_RAM.N_578\
        );

    \I__782\ : Odrv4
    port map (
            O => \N__5393\,
            I => \U712_CHIP_RAM.N_578\
        );

    \I__781\ : Odrv4
    port map (
            O => \N__5386\,
            I => \U712_CHIP_RAM.N_578\
        );

    \I__780\ : Odrv12
    port map (
            O => \N__5379\,
            I => \U712_CHIP_RAM.N_578\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__5376\,
            I => \U712_CHIP_RAM.N_578\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__5373\,
            I => \U712_CHIP_RAM.N_578\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__5370\,
            I => \U712_CHIP_RAM.N_578\
        );

    \I__776\ : InMux
    port map (
            O => \N__5353\,
            I => \N__5350\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__5350\,
            I => \N__5343\
        );

    \I__774\ : InMux
    port map (
            O => \N__5349\,
            I => \N__5337\
        );

    \I__773\ : InMux
    port map (
            O => \N__5348\,
            I => \N__5332\
        );

    \I__772\ : InMux
    port map (
            O => \N__5347\,
            I => \N__5332\
        );

    \I__771\ : InMux
    port map (
            O => \N__5346\,
            I => \N__5329\
        );

    \I__770\ : Span4Mux_h
    port map (
            O => \N__5343\,
            I => \N__5326\
        );

    \I__769\ : InMux
    port map (
            O => \N__5342\,
            I => \N__5323\
        );

    \I__768\ : InMux
    port map (
            O => \N__5341\,
            I => \N__5320\
        );

    \I__767\ : InMux
    port map (
            O => \N__5340\,
            I => \N__5317\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__5337\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__5332\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__5329\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__763\ : Odrv4
    port map (
            O => \N__5326\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__5323\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__5320\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__5317\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__759\ : InMux
    port map (
            O => \N__5302\,
            I => \N__5299\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__5299\,
            I => \U712_CHIP_RAM.N_405\
        );

    \I__757\ : InMux
    port map (
            O => \N__5296\,
            I => \N__5291\
        );

    \I__756\ : InMux
    port map (
            O => \N__5295\,
            I => \N__5288\
        );

    \I__755\ : InMux
    port map (
            O => \N__5294\,
            I => \N__5285\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__5291\,
            I => \U712_CHIP_RAM.N_699\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__5288\,
            I => \U712_CHIP_RAM.N_699\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__5285\,
            I => \U712_CHIP_RAM.N_699\
        );

    \I__751\ : CascadeMux
    port map (
            O => \N__5278\,
            I => \U712_CHIP_RAM.N_597_cascade_\
        );

    \I__750\ : CascadeMux
    port map (
            O => \N__5275\,
            I => \N__5272\
        );

    \I__749\ : InMux
    port map (
            O => \N__5272\,
            I => \N__5269\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__5269\,
            I => \N__5266\
        );

    \I__747\ : Odrv4
    port map (
            O => \N__5266\,
            I => \U712_CHIP_RAM.DMA_CYCLE_START_RNOZ0Z_0\
        );

    \I__746\ : InMux
    port map (
            O => \N__5263\,
            I => \N__5260\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__5260\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__744\ : IoInMux
    port map (
            O => \N__5257\,
            I => \N__5253\
        );

    \I__743\ : InMux
    port map (
            O => \N__5256\,
            I => \N__5250\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__5253\,
            I => \N__5247\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__5250\,
            I => \N__5244\
        );

    \I__740\ : IoSpan4Mux
    port map (
            O => \N__5247\,
            I => \N__5241\
        );

    \I__739\ : Span12Mux_h
    port map (
            O => \N__5244\,
            I => \N__5238\
        );

    \I__738\ : IoSpan4Mux
    port map (
            O => \N__5241\,
            I => \N__5235\
        );

    \I__737\ : Span12Mux_v
    port map (
            O => \N__5238\,
            I => \N__5232\
        );

    \I__736\ : IoSpan4Mux
    port map (
            O => \N__5235\,
            I => \N__5229\
        );

    \I__735\ : Odrv12
    port map (
            O => \N__5232\,
            I => \C1_c\
        );

    \I__734\ : Odrv4
    port map (
            O => \N__5229\,
            I => \C1_c\
        );

    \I__733\ : InMux
    port map (
            O => \N__5224\,
            I => \N__5221\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__5221\,
            I => \N__5218\
        );

    \I__731\ : Odrv4
    port map (
            O => \N__5218\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__730\ : CascadeMux
    port map (
            O => \N__5215\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1_cascade_\
        );

    \I__729\ : InMux
    port map (
            O => \N__5212\,
            I => \N__5209\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__5209\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\
        );

    \I__727\ : InMux
    port map (
            O => \N__5206\,
            I => \N__5202\
        );

    \I__726\ : CascadeMux
    port map (
            O => \N__5205\,
            I => \N__5199\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__5202\,
            I => \N__5195\
        );

    \I__724\ : InMux
    port map (
            O => \N__5199\,
            I => \N__5192\
        );

    \I__723\ : InMux
    port map (
            O => \N__5198\,
            I => \N__5189\
        );

    \I__722\ : Span4Mux_h
    port map (
            O => \N__5195\,
            I => \N__5186\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__5192\,
            I => \N__5181\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__5189\,
            I => \N__5181\
        );

    \I__719\ : Odrv4
    port map (
            O => \N__5186\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__718\ : Odrv4
    port map (
            O => \N__5181\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__717\ : InMux
    port map (
            O => \N__5176\,
            I => \N__5173\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__5173\,
            I => \N__5170\
        );

    \I__715\ : Odrv12
    port map (
            O => \N__5170\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5\
        );

    \I__714\ : CascadeMux
    port map (
            O => \N__5167\,
            I => \N__5164\
        );

    \I__713\ : InMux
    port map (
            O => \N__5164\,
            I => \N__5159\
        );

    \I__712\ : InMux
    port map (
            O => \N__5163\,
            I => \N__5154\
        );

    \I__711\ : InMux
    port map (
            O => \N__5162\,
            I => \N__5151\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__5159\,
            I => \N__5146\
        );

    \I__709\ : InMux
    port map (
            O => \N__5158\,
            I => \N__5141\
        );

    \I__708\ : InMux
    port map (
            O => \N__5157\,
            I => \N__5141\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__5154\,
            I => \N__5134\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__5151\,
            I => \N__5134\
        );

    \I__705\ : InMux
    port map (
            O => \N__5150\,
            I => \N__5129\
        );

    \I__704\ : InMux
    port map (
            O => \N__5149\,
            I => \N__5129\
        );

    \I__703\ : Span4Mux_h
    port map (
            O => \N__5146\,
            I => \N__5126\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__5141\,
            I => \N__5123\
        );

    \I__701\ : InMux
    port map (
            O => \N__5140\,
            I => \N__5120\
        );

    \I__700\ : InMux
    port map (
            O => \N__5139\,
            I => \N__5117\
        );

    \I__699\ : Odrv12
    port map (
            O => \N__5134\,
            I => \U712_CHIP_RAM.N_589\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__5129\,
            I => \U712_CHIP_RAM.N_589\
        );

    \I__697\ : Odrv4
    port map (
            O => \N__5126\,
            I => \U712_CHIP_RAM.N_589\
        );

    \I__696\ : Odrv4
    port map (
            O => \N__5123\,
            I => \U712_CHIP_RAM.N_589\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__5120\,
            I => \U712_CHIP_RAM.N_589\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__5117\,
            I => \U712_CHIP_RAM.N_589\
        );

    \I__693\ : CascadeMux
    port map (
            O => \N__5104\,
            I => \N__5100\
        );

    \I__692\ : InMux
    port map (
            O => \N__5103\,
            I => \N__5097\
        );

    \I__691\ : InMux
    port map (
            O => \N__5100\,
            I => \N__5094\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__5097\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__5094\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__688\ : CascadeMux
    port map (
            O => \N__5089\,
            I => \U712_REG_SM.N_694_cascade_\
        );

    \I__687\ : CascadeMux
    port map (
            O => \N__5086\,
            I => \U712_REG_SM.N_522_cascade_\
        );

    \I__686\ : IoInMux
    port map (
            O => \N__5083\,
            I => \N__5080\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__5080\,
            I => \N__5077\
        );

    \I__684\ : IoSpan4Mux
    port map (
            O => \N__5077\,
            I => \N__5074\
        );

    \I__683\ : Span4Mux_s3_h
    port map (
            O => \N__5074\,
            I => \N__5071\
        );

    \I__682\ : Span4Mux_h
    port map (
            O => \N__5071\,
            I => \N__5068\
        );

    \I__681\ : Span4Mux_h
    port map (
            O => \N__5068\,
            I => \N__5065\
        );

    \I__680\ : Span4Mux_h
    port map (
            O => \N__5065\,
            I => \N__5061\
        );

    \I__679\ : InMux
    port map (
            O => \N__5064\,
            I => \N__5058\
        );

    \I__678\ : Sp12to4
    port map (
            O => \N__5061\,
            I => \N__5053\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__5058\,
            I => \N__5053\
        );

    \I__676\ : Span12Mux_h
    port map (
            O => \N__5053\,
            I => \N__5050\
        );

    \I__675\ : Span12Mux_v
    port map (
            O => \N__5050\,
            I => \N__5047\
        );

    \I__674\ : Odrv12
    port map (
            O => \N__5047\,
            I => \C3_c\
        );

    \I__673\ : InMux
    port map (
            O => \N__5044\,
            I => \N__5041\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__5041\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__671\ : InMux
    port map (
            O => \N__5038\,
            I => \N__5034\
        );

    \I__670\ : InMux
    port map (
            O => \N__5037\,
            I => \N__5031\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__5034\,
            I => \U712_CHIP_RAM.N_697\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__5031\,
            I => \U712_CHIP_RAM.N_697\
        );

    \I__667\ : InMux
    port map (
            O => \N__5026\,
            I => \N__5023\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__5023\,
            I => \N__5019\
        );

    \I__665\ : InMux
    port map (
            O => \N__5022\,
            I => \N__5016\
        );

    \I__664\ : Span4Mux_h
    port map (
            O => \N__5019\,
            I => \N__5013\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__5016\,
            I => \N__5010\
        );

    \I__662\ : Odrv4
    port map (
            O => \N__5013\,
            I => \U712_CHIP_RAM.N_551\
        );

    \I__661\ : Odrv4
    port map (
            O => \N__5010\,
            I => \U712_CHIP_RAM.N_551\
        );

    \I__660\ : CascadeMux
    port map (
            O => \N__5005\,
            I => \N__4998\
        );

    \I__659\ : CascadeMux
    port map (
            O => \N__5004\,
            I => \N__4995\
        );

    \I__658\ : CascadeMux
    port map (
            O => \N__5003\,
            I => \N__4992\
        );

    \I__657\ : CascadeMux
    port map (
            O => \N__5002\,
            I => \N__4989\
        );

    \I__656\ : InMux
    port map (
            O => \N__5001\,
            I => \N__4986\
        );

    \I__655\ : InMux
    port map (
            O => \N__4998\,
            I => \N__4981\
        );

    \I__654\ : InMux
    port map (
            O => \N__4995\,
            I => \N__4981\
        );

    \I__653\ : InMux
    port map (
            O => \N__4992\,
            I => \N__4975\
        );

    \I__652\ : InMux
    port map (
            O => \N__4989\,
            I => \N__4975\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__4986\,
            I => \N__4967\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__4981\,
            I => \N__4967\
        );

    \I__649\ : InMux
    port map (
            O => \N__4980\,
            I => \N__4964\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__4975\,
            I => \N__4961\
        );

    \I__647\ : InMux
    port map (
            O => \N__4974\,
            I => \N__4956\
        );

    \I__646\ : InMux
    port map (
            O => \N__4973\,
            I => \N__4956\
        );

    \I__645\ : InMux
    port map (
            O => \N__4972\,
            I => \N__4953\
        );

    \I__644\ : Odrv4
    port map (
            O => \N__4967\,
            I => \U712_CHIP_RAM.N_580\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__4964\,
            I => \U712_CHIP_RAM.N_580\
        );

    \I__642\ : Odrv12
    port map (
            O => \N__4961\,
            I => \U712_CHIP_RAM.N_580\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__4956\,
            I => \U712_CHIP_RAM.N_580\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__4953\,
            I => \U712_CHIP_RAM.N_580\
        );

    \I__639\ : InMux
    port map (
            O => \N__4942\,
            I => \N__4939\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__4939\,
            I => \N__4936\
        );

    \I__637\ : Span4Mux_h
    port map (
            O => \N__4936\,
            I => \N__4933\
        );

    \I__636\ : Odrv4
    port map (
            O => \N__4933\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__635\ : InMux
    port map (
            O => \N__4930\,
            I => \N__4927\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__4927\,
            I => \N__4924\
        );

    \I__633\ : Odrv4
    port map (
            O => \N__4924\,
            I => \U712_CHIP_RAM.N_505\
        );

    \I__632\ : CascadeMux
    port map (
            O => \N__4921\,
            I => \N__4918\
        );

    \I__631\ : InMux
    port map (
            O => \N__4918\,
            I => \N__4915\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__4915\,
            I => \U712_CHIP_RAM.N_437\
        );

    \I__629\ : InMux
    port map (
            O => \N__4912\,
            I => \N__4909\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__4909\,
            I => \U712_CHIP_RAM.N_587\
        );

    \I__627\ : InMux
    port map (
            O => \N__4906\,
            I => \N__4903\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__4903\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__625\ : InMux
    port map (
            O => \N__4900\,
            I => \N__4884\
        );

    \I__624\ : InMux
    port map (
            O => \N__4899\,
            I => \N__4884\
        );

    \I__623\ : InMux
    port map (
            O => \N__4898\,
            I => \N__4884\
        );

    \I__622\ : InMux
    port map (
            O => \N__4897\,
            I => \N__4884\
        );

    \I__621\ : InMux
    port map (
            O => \N__4896\,
            I => \N__4879\
        );

    \I__620\ : InMux
    port map (
            O => \N__4895\,
            I => \N__4879\
        );

    \I__619\ : InMux
    port map (
            O => \N__4894\,
            I => \N__4874\
        );

    \I__618\ : InMux
    port map (
            O => \N__4893\,
            I => \N__4874\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__4884\,
            I => \U712_CHIP_RAM.N_70\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__4879\,
            I => \U712_CHIP_RAM.N_70\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__4874\,
            I => \U712_CHIP_RAM.N_70\
        );

    \I__614\ : CEMux
    port map (
            O => \N__4867\,
            I => \N__4863\
        );

    \I__613\ : CEMux
    port map (
            O => \N__4866\,
            I => \N__4860\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__4863\,
            I => \N__4857\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__4860\,
            I => \N__4854\
        );

    \I__610\ : Span4Mux_h
    port map (
            O => \N__4857\,
            I => \N__4851\
        );

    \I__609\ : Odrv4
    port map (
            O => \N__4854\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__608\ : Odrv4
    port map (
            O => \N__4851\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__607\ : InMux
    port map (
            O => \N__4846\,
            I => \N__4843\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__4843\,
            I => \N__4840\
        );

    \I__605\ : Span4Mux_v
    port map (
            O => \N__4840\,
            I => \N__4837\
        );

    \I__604\ : Sp12to4
    port map (
            O => \N__4837\,
            I => \N__4834\
        );

    \I__603\ : Span12Mux_h
    port map (
            O => \N__4834\,
            I => \N__4831\
        );

    \I__602\ : Odrv12
    port map (
            O => \N__4831\,
            I => \REGSPACEn_c\
        );

    \I__601\ : CascadeMux
    port map (
            O => \N__4828\,
            I => \U712_REG_SM.N_513_cascade_\
        );

    \I__600\ : InMux
    port map (
            O => \N__4825\,
            I => \N__4816\
        );

    \I__599\ : InMux
    port map (
            O => \N__4824\,
            I => \N__4805\
        );

    \I__598\ : InMux
    port map (
            O => \N__4823\,
            I => \N__4802\
        );

    \I__597\ : InMux
    port map (
            O => \N__4822\,
            I => \N__4797\
        );

    \I__596\ : InMux
    port map (
            O => \N__4821\,
            I => \N__4797\
        );

    \I__595\ : InMux
    port map (
            O => \N__4820\,
            I => \N__4792\
        );

    \I__594\ : InMux
    port map (
            O => \N__4819\,
            I => \N__4792\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__4816\,
            I => \N__4789\
        );

    \I__592\ : InMux
    port map (
            O => \N__4815\,
            I => \N__4786\
        );

    \I__591\ : InMux
    port map (
            O => \N__4814\,
            I => \N__4783\
        );

    \I__590\ : InMux
    port map (
            O => \N__4813\,
            I => \N__4778\
        );

    \I__589\ : InMux
    port map (
            O => \N__4812\,
            I => \N__4778\
        );

    \I__588\ : InMux
    port map (
            O => \N__4811\,
            I => \N__4775\
        );

    \I__587\ : InMux
    port map (
            O => \N__4810\,
            I => \N__4768\
        );

    \I__586\ : InMux
    port map (
            O => \N__4809\,
            I => \N__4768\
        );

    \I__585\ : InMux
    port map (
            O => \N__4808\,
            I => \N__4768\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__4805\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__4802\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__4797\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__4792\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__580\ : Odrv4
    port map (
            O => \N__4789\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__4786\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__4783\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__4778\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__4775\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__4768\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__574\ : InMux
    port map (
            O => \N__4747\,
            I => \N__4744\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__4744\,
            I => \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1\
        );

    \I__572\ : CascadeMux
    port map (
            O => \N__4741\,
            I => \U712_CHIP_RAM.N_697_cascade_\
        );

    \I__571\ : InMux
    port map (
            O => \N__4738\,
            I => \N__4735\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__4735\,
            I => \N__4732\
        );

    \I__569\ : Odrv4
    port map (
            O => \N__4732\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_2\
        );

    \I__568\ : CascadeMux
    port map (
            O => \N__4729\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_2_cascade_\
        );

    \I__567\ : InMux
    port map (
            O => \N__4726\,
            I => \N__4723\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__4723\,
            I => \U712_CHIP_RAM.N_539\
        );

    \I__565\ : CascadeMux
    port map (
            O => \N__4720\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_\
        );

    \I__564\ : CEMux
    port map (
            O => \N__4717\,
            I => \N__4714\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__4714\,
            I => \N__4711\
        );

    \I__562\ : Odrv4
    port map (
            O => \N__4711\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0\
        );

    \I__561\ : InMux
    port map (
            O => \N__4708\,
            I => \N__4705\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__4705\,
            I => \N__4698\
        );

    \I__559\ : InMux
    port map (
            O => \N__4704\,
            I => \N__4695\
        );

    \I__558\ : InMux
    port map (
            O => \N__4703\,
            I => \N__4692\
        );

    \I__557\ : InMux
    port map (
            O => \N__4702\,
            I => \N__4687\
        );

    \I__556\ : InMux
    port map (
            O => \N__4701\,
            I => \N__4687\
        );

    \I__555\ : Odrv4
    port map (
            O => \N__4698\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__4695\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__4692\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__4687\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__551\ : CascadeMux
    port map (
            O => \N__4678\,
            I => \U712_CHIP_RAM.N_442_cascade_\
        );

    \I__550\ : InMux
    port map (
            O => \N__4675\,
            I => \N__4672\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__4672\,
            I => \U712_CHIP_RAM.BANK0_RNOZ0Z_3\
        );

    \I__548\ : CascadeMux
    port map (
            O => \N__4669\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_\
        );

    \I__547\ : InMux
    port map (
            O => \N__4666\,
            I => \N__4663\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__4663\,
            I => \U712_CHIP_RAM.BANK0_RNOZ0Z_1\
        );

    \I__545\ : InMux
    port map (
            O => \N__4660\,
            I => \N__4657\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__4657\,
            I => \N__4654\
        );

    \I__543\ : Span4Mux_h
    port map (
            O => \N__4654\,
            I => \N__4651\
        );

    \I__542\ : Span4Mux_v
    port map (
            O => \N__4651\,
            I => \N__4648\
        );

    \I__541\ : Sp12to4
    port map (
            O => \N__4648\,
            I => \N__4645\
        );

    \I__540\ : Odrv12
    port map (
            O => \N__4645\,
            I => \A_c_20\
        );

    \I__539\ : InMux
    port map (
            O => \N__4642\,
            I => \N__4639\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__4639\,
            I => \N__4636\
        );

    \I__537\ : Odrv12
    port map (
            O => \N__4636\,
            I => \U712_CHIP_RAM.BANK0_RNOZ0Z_2\
        );

    \I__536\ : CascadeMux
    port map (
            O => \N__4633\,
            I => \U712_CHIP_RAM.N_605_cascade_\
        );

    \I__535\ : InMux
    port map (
            O => \N__4630\,
            I => \N__4626\
        );

    \I__534\ : InMux
    port map (
            O => \N__4629\,
            I => \N__4623\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__4626\,
            I => \N__4620\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__4623\,
            I => \U712_CHIP_RAM.N_605\
        );

    \I__531\ : Odrv4
    port map (
            O => \N__4620\,
            I => \U712_CHIP_RAM.N_605\
        );

    \I__530\ : CascadeMux
    port map (
            O => \N__4615\,
            I => \U712_CHIP_RAM.N_554_cascade_\
        );

    \I__529\ : IoInMux
    port map (
            O => \N__4612\,
            I => \N__4609\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__4609\,
            I => \N__4606\
        );

    \I__527\ : Span4Mux_s1_v
    port map (
            O => \N__4606\,
            I => \N__4603\
        );

    \I__526\ : Sp12to4
    port map (
            O => \N__4603\,
            I => \N__4600\
        );

    \I__525\ : Span12Mux_h
    port map (
            O => \N__4600\,
            I => \N__4597\
        );

    \I__524\ : Span12Mux_v
    port map (
            O => \N__4597\,
            I => \N__4593\
        );

    \I__523\ : InMux
    port map (
            O => \N__4596\,
            I => \N__4590\
        );

    \I__522\ : Odrv12
    port map (
            O => \N__4593\,
            I => \BANK0_c\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__4590\,
            I => \BANK0_c\
        );

    \I__520\ : InMux
    port map (
            O => \N__4585\,
            I => \N__4582\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__4582\,
            I => \U712_CHIP_RAM.N_588\
        );

    \I__518\ : CascadeMux
    port map (
            O => \N__4579\,
            I => \U712_CHIP_RAM.N_553_cascade_\
        );

    \I__517\ : CascadeMux
    port map (
            O => \N__4576\,
            I => \U712_CHIP_RAM.N_437_cascade_\
        );

    \I__516\ : InMux
    port map (
            O => \N__4573\,
            I => \N__4569\
        );

    \I__515\ : InMux
    port map (
            O => \N__4572\,
            I => \N__4566\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__4569\,
            I => \U712_CHIP_RAM.N_414\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__4566\,
            I => \U712_CHIP_RAM.N_414\
        );

    \I__512\ : InMux
    port map (
            O => \N__4561\,
            I => \N__4558\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__4558\,
            I => \U712_CHIP_RAM.N_507\
        );

    \I__510\ : CascadeMux
    port map (
            O => \N__4555\,
            I => \U712_CHIP_RAM.N_507_cascade_\
        );

    \I__509\ : InMux
    port map (
            O => \N__4552\,
            I => \N__4549\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__4549\,
            I => \N__4546\
        );

    \I__507\ : Odrv4
    port map (
            O => \N__4546\,
            I => \U712_CHIP_RAM.N_506\
        );

    \I__506\ : CascadeMux
    port map (
            O => \N__4543\,
            I => \N__4539\
        );

    \I__505\ : InMux
    port map (
            O => \N__4542\,
            I => \N__4536\
        );

    \I__504\ : InMux
    port map (
            O => \N__4539\,
            I => \N__4532\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4536\,
            I => \N__4529\
        );

    \I__502\ : InMux
    port map (
            O => \N__4535\,
            I => \N__4526\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__4532\,
            I => \U712_CHIP_RAM.N_696\
        );

    \I__500\ : Odrv4
    port map (
            O => \N__4529\,
            I => \U712_CHIP_RAM.N_696\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__4526\,
            I => \U712_CHIP_RAM.N_696\
        );

    \I__498\ : InMux
    port map (
            O => \N__4519\,
            I => \N__4516\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__4516\,
            I => \N__4513\
        );

    \I__496\ : Odrv4
    port map (
            O => \N__4513\,
            I => \U712_CHIP_RAM.N_534\
        );

    \I__495\ : InMux
    port map (
            O => \N__4510\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__494\ : InMux
    port map (
            O => \N__4507\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__493\ : InMux
    port map (
            O => \N__4504\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__492\ : InMux
    port map (
            O => \N__4501\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__491\ : InMux
    port map (
            O => \N__4498\,
            I => \N__4494\
        );

    \I__490\ : InMux
    port map (
            O => \N__4497\,
            I => \N__4491\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__4494\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__4491\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__487\ : InMux
    port map (
            O => \N__4486\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__486\ : InMux
    port map (
            O => \N__4483\,
            I => \N__4479\
        );

    \I__485\ : InMux
    port map (
            O => \N__4482\,
            I => \N__4476\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__4479\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__4476\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__482\ : InMux
    port map (
            O => \N__4471\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__481\ : InMux
    port map (
            O => \N__4468\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__480\ : InMux
    port map (
            O => \N__4465\,
            I => \N__4461\
        );

    \I__479\ : InMux
    port map (
            O => \N__4464\,
            I => \N__4458\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__4461\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__4458\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__476\ : InMux
    port map (
            O => \N__4453\,
            I => \N__4450\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__4450\,
            I => \N__4447\
        );

    \I__474\ : Span4Mux_h
    port map (
            O => \N__4447\,
            I => \N__4444\
        );

    \I__473\ : Sp12to4
    port map (
            O => \N__4444\,
            I => \N__4441\
        );

    \I__472\ : Span12Mux_v
    port map (
            O => \N__4441\,
            I => \N__4438\
        );

    \I__471\ : Odrv12
    port map (
            O => \N__4438\,
            I => \A_c_8\
        );

    \I__470\ : InMux
    port map (
            O => \N__4435\,
            I => \N__4432\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__4432\,
            I => \N__4429\
        );

    \I__468\ : Span12Mux_v
    port map (
            O => \N__4429\,
            I => \N__4426\
        );

    \I__467\ : Odrv12
    port map (
            O => \N__4426\,
            I => \A_c_15\
        );

    \I__466\ : CascadeMux
    port map (
            O => \N__4423\,
            I => \U712_CHIP_RAM.N_578_cascade_\
        );

    \I__465\ : InMux
    port map (
            O => \N__4420\,
            I => \N__4417\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__4417\,
            I => \U712_CHIP_RAM.N_545\
        );

    \I__463\ : CascadeMux
    port map (
            O => \N__4414\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER18_cascade_\
        );

    \I__462\ : CascadeMux
    port map (
            O => \N__4411\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0_cascade_\
        );

    \I__461\ : InMux
    port map (
            O => \N__4408\,
            I => \N__4405\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__4405\,
            I => \U712_CHIP_RAM.N_552\
        );

    \I__459\ : CascadeMux
    port map (
            O => \N__4402\,
            I => \U712_CHIP_RAM.N_504_cascade_\
        );

    \I__458\ : InMux
    port map (
            O => \N__4399\,
            I => \N__4396\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__4396\,
            I => \N__4393\
        );

    \I__456\ : Odrv4
    port map (
            O => \N__4393\,
            I => \U712_CHIP_RAM.N_404\
        );

    \I__455\ : CascadeMux
    port map (
            O => \N__4390\,
            I => \U712_CHIP_RAM.N_404_cascade_\
        );

    \I__454\ : InMux
    port map (
            O => \N__4387\,
            I => \N__4384\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__4384\,
            I => \N__4381\
        );

    \I__452\ : Span4Mux_v
    port map (
            O => \N__4381\,
            I => \N__4378\
        );

    \I__451\ : Span4Mux_v
    port map (
            O => \N__4378\,
            I => \N__4375\
        );

    \I__450\ : Sp12to4
    port map (
            O => \N__4375\,
            I => \N__4372\
        );

    \I__449\ : Odrv12
    port map (
            O => \N__4372\,
            I => \A_c_5\
        );

    \I__448\ : InMux
    port map (
            O => \N__4369\,
            I => \N__4366\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__4366\,
            I => \N__4363\
        );

    \I__446\ : Span4Mux_v
    port map (
            O => \N__4363\,
            I => \N__4360\
        );

    \I__445\ : Sp12to4
    port map (
            O => \N__4360\,
            I => \N__4357\
        );

    \I__444\ : Odrv12
    port map (
            O => \N__4357\,
            I => \A_c_12\
        );

    \I__443\ : InMux
    port map (
            O => \N__4354\,
            I => \N__4351\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__4351\,
            I => \U712_CHIP_RAM.N_591\
        );

    \I__441\ : IoInMux
    port map (
            O => \N__4348\,
            I => \N__4345\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__4345\,
            I => \N__4342\
        );

    \I__439\ : Span12Mux_s9_v
    port map (
            O => \N__4342\,
            I => \N__4339\
        );

    \I__438\ : Odrv12
    port map (
            O => \N__4339\,
            I => \VBENn_c\
        );

    \I__437\ : InMux
    port map (
            O => \N__4336\,
            I => \N__4333\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__4333\,
            I => \N__4330\
        );

    \I__435\ : Span4Mux_v
    port map (
            O => \N__4330\,
            I => \N__4327\
        );

    \I__434\ : Span4Mux_v
    port map (
            O => \N__4327\,
            I => \N__4324\
        );

    \I__433\ : Sp12to4
    port map (
            O => \N__4324\,
            I => \N__4321\
        );

    \I__432\ : Odrv12
    port map (
            O => \N__4321\,
            I => \A_c_14\
        );

    \I__431\ : InMux
    port map (
            O => \N__4318\,
            I => \N__4315\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__4315\,
            I => \N__4312\
        );

    \I__429\ : Span4Mux_v
    port map (
            O => \N__4312\,
            I => \N__4309\
        );

    \I__428\ : Span4Mux_v
    port map (
            O => \N__4309\,
            I => \N__4306\
        );

    \I__427\ : Sp12to4
    port map (
            O => \N__4306\,
            I => \N__4303\
        );

    \I__426\ : Odrv12
    port map (
            O => \N__4303\,
            I => \A_c_7\
        );

    \I__425\ : CascadeMux
    port map (
            O => \N__4300\,
            I => \U712_CHIP_RAM.N_543_cascade_\
        );

    \I__424\ : CascadeMux
    port map (
            O => \N__4297\,
            I => \U712_CHIP_RAM.N_322_cascade_\
        );

    \I__423\ : InMux
    port map (
            O => \N__4294\,
            I => \N__4291\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__4291\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_a2_0_0\
        );

    \I__421\ : InMux
    port map (
            O => \N__4288\,
            I => \N__4285\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__4285\,
            I => \U712_CHIP_RAM.CLK_EN_6_0_a3_0_a2_1\
        );

    \I__419\ : CascadeMux
    port map (
            O => \N__4282\,
            I => \U712_CHIP_RAM.N_599_cascade_\
        );

    \I__418\ : InMux
    port map (
            O => \N__4279\,
            I => \N__4276\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__4276\,
            I => \U712_CHIP_RAM.CLK_EN_6_0\
        );

    \I__416\ : IoInMux
    port map (
            O => \N__4273\,
            I => \N__4270\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__4270\,
            I => \N__4267\
        );

    \I__414\ : Span4Mux_s1_v
    port map (
            O => \N__4267\,
            I => \N__4264\
        );

    \I__413\ : Span4Mux_v
    port map (
            O => \N__4264\,
            I => \N__4261\
        );

    \I__412\ : Span4Mux_v
    port map (
            O => \N__4261\,
            I => \N__4258\
        );

    \I__411\ : Span4Mux_v
    port map (
            O => \N__4258\,
            I => \N__4255\
        );

    \I__410\ : Odrv4
    port map (
            O => \N__4255\,
            I => \U712_CYCLE_TERM_TBIn_0_i\
        );

    \I__409\ : IoInMux
    port map (
            O => \N__4252\,
            I => \N__4249\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__4249\,
            I => \N__4246\
        );

    \I__407\ : Span4Mux_s2_v
    port map (
            O => \N__4246\,
            I => \N__4243\
        );

    \I__406\ : Span4Mux_v
    port map (
            O => \N__4243\,
            I => \N__4240\
        );

    \I__405\ : Span4Mux_h
    port map (
            O => \N__4240\,
            I => \N__4237\
        );

    \I__404\ : Odrv4
    port map (
            O => \N__4237\,
            I => \CLK80_PLL_i_i\
        );

    \I__403\ : IoInMux
    port map (
            O => \N__4234\,
            I => \N__4231\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__4231\,
            I => \N__4228\
        );

    \I__401\ : IoSpan4Mux
    port map (
            O => \N__4228\,
            I => \N__4225\
        );

    \I__400\ : Span4Mux_s3_h
    port map (
            O => \N__4225\,
            I => \N__4222\
        );

    \I__399\ : Span4Mux_h
    port map (
            O => \N__4222\,
            I => \N__4219\
        );

    \I__398\ : Odrv4
    port map (
            O => \N__4219\,
            I => \DBRn_c_i_0\
        );

    \I__397\ : IoInMux
    port map (
            O => \N__4216\,
            I => \N__4213\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__4213\,
            I => \N__4210\
        );

    \I__395\ : Span12Mux_s10_h
    port map (
            O => \N__4210\,
            I => \N__4207\
        );

    \I__394\ : Span12Mux_h
    port map (
            O => \N__4207\,
            I => \N__4203\
        );

    \I__393\ : InMux
    port map (
            O => \N__4206\,
            I => \N__4200\
        );

    \I__392\ : Odrv12
    port map (
            O => \N__4203\,
            I => \CLK_EN_c\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__4200\,
            I => \CLK_EN_c\
        );

    \I__390\ : InMux
    port map (
            O => \N__4195\,
            I => \N__4191\
        );

    \I__389\ : InMux
    port map (
            O => \N__4194\,
            I => \N__4188\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__4191\,
            I => \N__4183\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__4188\,
            I => \N__4183\
        );

    \I__386\ : Span12Mux_h
    port map (
            O => \N__4183\,
            I => \N__4180\
        );

    \I__385\ : Span12Mux_v
    port map (
            O => \N__4180\,
            I => \N__4177\
        );

    \I__384\ : Odrv12
    port map (
            O => \N__4177\,
            I => \DBRn_c\
        );

    \I__383\ : InMux
    port map (
            O => \N__4174\,
            I => \N__4171\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__4171\,
            I => \N__4168\
        );

    \I__381\ : Odrv4
    port map (
            O => \N__4168\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__380\ : InMux
    port map (
            O => \N__4165\,
            I => \N__4162\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__4162\,
            I => \N__4159\
        );

    \I__378\ : Span4Mux_v
    port map (
            O => \N__4159\,
            I => \N__4156\
        );

    \I__377\ : Span4Mux_v
    port map (
            O => \N__4156\,
            I => \N__4153\
        );

    \I__376\ : Sp12to4
    port map (
            O => \N__4153\,
            I => \N__4150\
        );

    \I__375\ : Odrv12
    port map (
            O => \N__4150\,
            I => \A_c_18\
        );

    \I__374\ : InMux
    port map (
            O => \N__4147\,
            I => \N__4144\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__4144\,
            I => \N__4141\
        );

    \I__372\ : Span4Mux_v
    port map (
            O => \N__4141\,
            I => \N__4138\
        );

    \I__371\ : Span4Mux_v
    port map (
            O => \N__4138\,
            I => \N__4135\
        );

    \I__370\ : Sp12to4
    port map (
            O => \N__4135\,
            I => \N__4132\
        );

    \I__369\ : Odrv12
    port map (
            O => \N__4132\,
            I => \A_c_16\
        );

    \I__368\ : InMux
    port map (
            O => \N__4129\,
            I => \N__4126\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__4126\,
            I => \N__4123\
        );

    \I__366\ : Span4Mux_v
    port map (
            O => \N__4123\,
            I => \N__4120\
        );

    \I__365\ : Span4Mux_v
    port map (
            O => \N__4120\,
            I => \N__4117\
        );

    \I__364\ : Sp12to4
    port map (
            O => \N__4117\,
            I => \N__4114\
        );

    \I__363\ : Odrv12
    port map (
            O => \N__4114\,
            I => \A_c_6\
        );

    \I__362\ : InMux
    port map (
            O => \N__4111\,
            I => \N__4108\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__4108\,
            I => \N__4105\
        );

    \I__360\ : Odrv12
    port map (
            O => \N__4105\,
            I => \A_c_13\
        );

    \I__359\ : IoInMux
    port map (
            O => \N__4102\,
            I => \N__4099\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__4099\,
            I => \N__4096\
        );

    \I__357\ : IoSpan4Mux
    port map (
            O => \N__4096\,
            I => \N__4093\
        );

    \I__356\ : Span4Mux_s2_v
    port map (
            O => \N__4093\,
            I => \N__4090\
        );

    \I__355\ : Sp12to4
    port map (
            O => \N__4090\,
            I => \N__4087\
        );

    \I__354\ : Span12Mux_v
    port map (
            O => \N__4087\,
            I => \N__4084\
        );

    \I__353\ : Odrv12
    port map (
            O => \N__4084\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__6861\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            I => \N__6863\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            I => \N__6865\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            I => \N__6860\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__6862\
        );

    \INVU712_CHIP_RAM.DMA_A20C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A20C_net\,
            I => \N__6858\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            I => \N__6859\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_11_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_5_0_\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5257\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6409\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4234\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5083\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_OUTn_RNI3QLB_LC_3_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__7665\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7599\,
            lcout => \U712_CYCLE_TERM_TBIn_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8803\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBRn_ibuf_RNIBAB_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4194\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBRn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9285\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10279\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__4206\,
            in1 => \N__4279\,
            in2 => \_gnd_net_\,
            in3 => \N__5479\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8787\,
            ce => 'H',
            sr => \N__10259\
        );

    \DBR_SYNC_1_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4174\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8791\,
            ce => 'H',
            sr => \N__10256\
        );

    \DBR_SYNC_0_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4195\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8797\,
            ce => 'H',
            sr => \N__10244\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4165\,
            in1 => \N__4147\,
            in2 => \_gnd_net_\,
            in3 => \N__9035\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4129\,
            in1 => \N__4111\,
            in2 => \_gnd_net_\,
            in3 => \N__8997\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_3_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__9585\,
            in1 => \N__7178\,
            in2 => \_gnd_net_\,
            in3 => \N__5978\,
            lcout => \U712_CHIP_RAM.CLK_EN_6_0_a3_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4336\,
            in1 => \N__4318\,
            in2 => \_gnd_net_\,
            in3 => \N__8996\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4399\,
            in1 => \N__4630\,
            in2 => \N__5448\,
            in3 => \N__5348\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_543_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__4294\,
            in1 => \N__4420\,
            in2 => \N__4300\,
            in3 => \N__5001\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_322_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6151\,
            in2 => \N__4297\,
            in3 => \N__9002\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8782\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__4821\,
            in1 => \N__8026\,
            in2 => \N__5983\,
            in3 => \N__6109\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_2_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__4822\,
            in1 => \N__7801\,
            in2 => \_gnd_net_\,
            in3 => \N__6108\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_599_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__4288\,
            in1 => \N__5347\,
            in2 => \N__4282\,
            in3 => \N__5426\,
            lcout => \U712_CHIP_RAM.CLK_EN_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101110"
        )
    port map (
            in0 => \N__4519\,
            in1 => \N__9633\,
            in2 => \N__7802\,
            in3 => \N__7161\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8788\,
            ce => \N__4717\,
            sr => \N__10250\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_1_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__7783\,
            in1 => \N__4972\,
            in2 => \N__6106\,
            in3 => \N__4812\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_504_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5PDS6_3_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__4813\,
            in1 => \N__6093\,
            in2 => \N__4402\,
            in3 => \N__4535\,
            lcout => \U712_CHIP_RAM.N_414\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI85LA2_4_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7782\,
            in1 => \N__5341\,
            in2 => \_gnd_net_\,
            in3 => \N__5402\,
            lcout => \U712_CHIP_RAM.N_696\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001101000000"
        )
    port map (
            in0 => \N__4814\,
            in1 => \N__6097\,
            in2 => \N__5976\,
            in3 => \N__7793\,
            lcout => \U712_CHIP_RAM.N_404\,
            ltout => \U712_CHIP_RAM.N_404_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIM81M2_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__5342\,
            in1 => \_gnd_net_\,
            in2 => \N__4390\,
            in3 => \N__4708\,
            lcout => \U712_CHIP_RAM.N_591\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5958\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4573\,
            lcout => \U712_CHIP_RAM.N_505\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4387\,
            in1 => \N__4369\,
            in2 => \_gnd_net_\,
            in3 => \N__9022\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010001000"
        )
    port map (
            in0 => \N__5954\,
            in1 => \N__7792\,
            in2 => \N__6107\,
            in3 => \N__7132\,
            lcout => \U712_CHIP_RAM.N_588\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIF4EE6_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__4354\,
            in1 => \N__8025\,
            in2 => \N__5167\,
            in3 => \N__5446\,
            lcout => \U712_CHIP_RAM.N_551\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_0_a3_0_a2_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9616\,
            in2 => \_gnd_net_\,
            in3 => \N__10119\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4453\,
            in1 => \N__4435\,
            in2 => \_gnd_net_\,
            in3 => \N__9001\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4464\,
            in1 => \N__4482\,
            in2 => \_gnd_net_\,
            in3 => \N__4497\,
            lcout => \U712_CHIP_RAM.N_578\,
            ltout => \U712_CHIP_RAM.N_578_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__5340\,
            in1 => \_gnd_net_\,
            in2 => \N__4423\,
            in3 => \N__4701\,
            lcout => \U712_CHIP_RAM.N_580\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5206\,
            in1 => \N__8030\,
            in2 => \N__6670\,
            in3 => \N__6759\,
            lcout => \U712_CHIP_RAM.N_545\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5982\,
            in1 => \N__6104\,
            in2 => \N__4543\,
            in3 => \N__4824\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__4702\,
            in1 => \_gnd_net_\,
            in2 => \N__4414\,
            in3 => \N__8031\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8778\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011010001"
        )
    port map (
            in0 => \N__4408\,
            in1 => \N__6150\,
            in2 => \N__9161\,
            in3 => \N__5022\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8778\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIM2QU_3_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8032\,
            in2 => \_gnd_net_\,
            in3 => \N__4811\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIMEP34_1_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000000000000"
        )
    port map (
            in0 => \N__7794\,
            in1 => \N__6103\,
            in2 => \N__4411\,
            in3 => \N__4980\,
            lcout => \U712_CHIP_RAM.N_506\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6062\,
            in2 => \_gnd_net_\,
            in3 => \N__5037\,
            lcout => \U712_CHIP_RAM.N_552\,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4897\,
            in1 => \N__7800\,
            in2 => \_gnd_net_\,
            in3 => \N__4510\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__8783\,
            ce => \N__4866\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5953\,
            in2 => \_gnd_net_\,
            in3 => \N__4507\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4898\,
            in1 => \N__4823\,
            in2 => \_gnd_net_\,
            in3 => \N__4504\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__8783\,
            ce => \N__4866\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4893\,
            in1 => \N__5349\,
            in2 => \_gnd_net_\,
            in3 => \N__4501\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__8783\,
            ce => \N__4866\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4899\,
            in1 => \N__4498\,
            in2 => \_gnd_net_\,
            in3 => \N__4486\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__8783\,
            ce => \N__4866\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4894\,
            in1 => \N__4483\,
            in2 => \_gnd_net_\,
            in3 => \N__4471\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__8783\,
            ce => \N__4866\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4900\,
            in1 => \N__4465\,
            in2 => \_gnd_net_\,
            in3 => \N__4468\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8783\,
            ce => \N__4866\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__5830\,
            in1 => \N__6760\,
            in2 => \N__5003\,
            in3 => \N__5150\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_554_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__4596\,
            in1 => \N__5523\,
            in2 => \N__4615\,
            in3 => \N__4666\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8789\,
            ce => 'H',
            sr => \N__10236\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITIV55_3_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__4912\,
            in1 => \N__4815\,
            in2 => \N__5002\,
            in3 => \N__4585\,
            lcout => \U712_CHIP_RAM.N_553\,
            ltout => \U712_CHIP_RAM.N_553_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIJSRL5_3_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4579\,
            in3 => \N__7988\,
            lcout => \U712_CHIP_RAM.N_437\,
            ltout => \U712_CHIP_RAM.N_437_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIG9KPG_2_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__4561\,
            in1 => \N__5432\,
            in2 => \N__4576\,
            in3 => \N__5149\,
            lcout => \U712_CHIP_RAM.N_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQQ7R7_2_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5948\,
            in1 => \N__7989\,
            in2 => \_gnd_net_\,
            in3 => \N__4572\,
            lcout => \U712_CHIP_RAM.N_507\,
            ltout => \U712_CHIP_RAM.N_507_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVVPHH_1_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__6653\,
            in1 => \N__4738\,
            in2 => \N__4555\,
            in3 => \N__4552\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7143\,
            in1 => \N__4542\,
            in2 => \N__5975\,
            in3 => \N__4747\,
            lcout => \U712_CHIP_RAM.N_534\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_3_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__5157\,
            in1 => \N__6747\,
            in2 => \_gnd_net_\,
            in3 => \N__5430\,
            lcout => \U712_CHIP_RAM.BANK0_RNOZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__6751\,
            in1 => \N__7228\,
            in2 => \_gnd_net_\,
            in3 => \N__5784\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_442_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__8007\,
            in1 => \N__5103\,
            in2 => \N__4678\,
            in3 => \N__7144\,
            lcout => \WRITE_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8792\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIURFN4_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5834\,
            in1 => \N__5431\,
            in2 => \N__6761\,
            in3 => \N__5158\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_1_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101010000"
        )
    port map (
            in0 => \N__4642\,
            in1 => \N__4675\,
            in2 => \N__4669\,
            in3 => \N__9274\,
            lcout => \U712_CHIP_RAM.BANK0_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7533\,
            in2 => \_gnd_net_\,
            in3 => \N__6105\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_2_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__4660\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10613\,
            lcout => \U712_CHIP_RAM.BANK0_RNOZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5836\,
            in1 => \N__5163\,
            in2 => \N__5445\,
            in3 => \N__6738\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8773\,
            ce => \N__5797\,
            sr => \N__10251\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__8028\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4704\,
            lcout => \U712_CHIP_RAM.N_605\,
            ltout => \U712_CHIP_RAM.N_605_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__5963\,
            in1 => \N__4820\,
            in2 => \N__4633\,
            in3 => \N__6088\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_0_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKCP34_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4629\,
            in1 => \N__5140\,
            in2 => \_gnd_net_\,
            in3 => \N__5404\,
            lcout => \U712_CHIP_RAM.N_700\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIONRK3_1_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5964\,
            in1 => \N__8029\,
            in2 => \N__5005\,
            in3 => \N__7796\,
            lcout => \U712_CHIP_RAM.N_697\,
            ltout => \U712_CHIP_RAM.N_697_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__6089\,
            in1 => \_gnd_net_\,
            in2 => \N__4741\,
            in3 => \N__7160\,
            lcout => \U712_CHIP_RAM.N_537\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIHJRU1_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__5302\,
            in1 => \N__8027\,
            in2 => \N__5205\,
            in3 => \N__6737\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_2\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4TF5A_4_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__5467\,
            in1 => \N__6654\,
            in2 => \N__4729\,
            in3 => \N__5346\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5962\,
            in1 => \N__4819\,
            in2 => \N__5004\,
            in3 => \N__7795\,
            lcout => \U712_CHIP_RAM.N_539\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__4726\,
            in1 => \N__5926\,
            in2 => \N__5665\,
            in3 => \N__5295\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4720\,
            in3 => \N__10278\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU2TJ3_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5139\,
            in1 => \N__4703\,
            in2 => \_gnd_net_\,
            in3 => \N__5403\,
            lcout => \U712_CHIP_RAM.N_595\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIEH9V_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__5646\,
            in1 => \N__5198\,
            in2 => \_gnd_net_\,
            in3 => \N__5541\,
            lcout => \U712_CHIP_RAM.N_600\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_1_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4809\,
            in1 => \N__7790\,
            in2 => \_gnd_net_\,
            in3 => \N__4973\,
            lcout => \U712_CHIP_RAM.N_703\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011010001"
        )
    port map (
            in0 => \N__5038\,
            in1 => \N__6145\,
            in2 => \N__8352\,
            in3 => \N__5026\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8779\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_1_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__4810\,
            in1 => \N__7791\,
            in2 => \N__6086\,
            in3 => \N__4974\,
            lcout => \U712_CHIP_RAM.N_699\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_1_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5925\,
            in1 => \N__6048\,
            in2 => \N__7803\,
            in3 => \N__4808\,
            lcout => \U712_CHIP_RAM.N_589\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001110101010"
        )
    port map (
            in0 => \N__4942\,
            in1 => \N__4930\,
            in2 => \N__4921\,
            in3 => \N__4895\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8784\,
            ce => \N__4867\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI57LV_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9770\,
            in1 => \N__5927\,
            in2 => \_gnd_net_\,
            in3 => \N__6052\,
            lcout => \U712_CHIP_RAM.N_587\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__7987\,
            in1 => \N__4906\,
            in2 => \N__5104\,
            in3 => \N__4896\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8784\,
            ce => \N__4867\,
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5706\,
            in2 => \_gnd_net_\,
            in3 => \N__6218\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_513_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011000100"
        )
    port map (
            in0 => \N__4846\,
            in1 => \N__7986\,
            in2 => \N__4828\,
            in3 => \N__5565\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8790\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__9579\,
            in1 => \N__4825\,
            in2 => \_gnd_net_\,
            in3 => \N__6061\,
            lcout => \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5162\,
            in1 => \N__5449\,
            in2 => \_gnd_net_\,
            in3 => \N__9967\,
            lcout => \U712_CHIP_RAM.DBENn_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIPCS25_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__6752\,
            in1 => \N__5835\,
            in2 => \_gnd_net_\,
            in3 => \N__6665\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI347S_1_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6578\,
            in1 => \N__6512\,
            in2 => \_gnd_net_\,
            in3 => \N__5650\,
            lcout => \U712_REG_SM.N_694\,
            ltout => \U712_REG_SM.N_694_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_0_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5089\,
            in3 => \N__6259\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_522_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011100100"
        )
    port map (
            in0 => \N__7985\,
            in1 => \N__10106\,
            in2 => \N__5086\,
            in3 => \N__6928\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8793\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011101100"
        )
    port map (
            in0 => \N__7984\,
            in1 => \N__6736\,
            in2 => \N__5275\,
            in3 => \N__9774\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8793\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_0_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5064\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8795\,
            ce => 'H',
            sr => \N__10215\
        );

    \U712_REG_SM.C3_SYNC_1_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5044\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8795\,
            ce => 'H',
            sr => \N__10215\
        );

    \U712_REG_SM.C1_SYNC_1_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5224\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8795\,
            ce => 'H',
            sr => \N__10215\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5263\,
            in2 => \_gnd_net_\,
            in3 => \N__6417\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_START_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6418\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7975\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8798\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_0_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5256\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8799\,
            ce => 'H',
            sr => \N__10213\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__6342\,
            in1 => \N__6357\,
            in2 => \N__6313\,
            in3 => \N__6372\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6876\,
            in1 => \N__6894\,
            in2 => \_gnd_net_\,
            in3 => \N__6909\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010001100"
        )
    port map (
            in0 => \N__6327\,
            in1 => \N__8024\,
            in2 => \N__5215\,
            in3 => \N__5212\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8766\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__5545\,
            in1 => \N__9578\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_527\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__9577\,
            in1 => \N__5176\,
            in2 => \N__9301\,
            in3 => \N__9068\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__7301\,
            in1 => \N__6594\,
            in2 => \_gnd_net_\,
            in3 => \N__6535\,
            lcout => \U712_REG_SM.N_514\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6240\,
            in2 => \_gnd_net_\,
            in3 => \N__6274\,
            lcout => \U712_REG_SM.N_422\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6595\,
            in2 => \_gnd_net_\,
            in3 => \N__6536\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_429_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__8022\,
            in1 => \N__6199\,
            in2 => \N__5497\,
            in3 => \N__6275\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8774\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__6241\,
            in1 => \N__6596\,
            in2 => \_gnd_net_\,
            in3 => \N__6537\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_511_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__8023\,
            in1 => \N__7037\,
            in2 => \N__5494\,
            in3 => \N__5491\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8774\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__9739\,
            in1 => \N__5968\,
            in2 => \_gnd_net_\,
            in3 => \N__5296\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101010"
        )
    port map (
            in0 => \N__5466\,
            in1 => \N__5455\,
            in2 => \N__5447\,
            in3 => \N__5353\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__5540\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5644\,
            lcout => \U712_CHIP_RAM.N_405\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8MK44_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9757\,
            in1 => \N__5942\,
            in2 => \_gnd_net_\,
            in3 => \N__5294\,
            lcout => \U712_CHIP_RAM.N_597\,
            ltout => \U712_CHIP_RAM.N_597_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__6762\,
            in1 => \N__6661\,
            in2 => \N__5278\,
            in3 => \N__5664\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100010101000"
        )
    port map (
            in0 => \N__7999\,
            in1 => \N__5676\,
            in2 => \N__5695\,
            in3 => \N__7729\,
            lcout => \LATCH_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIOBA64_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__5941\,
            in1 => \N__7167\,
            in2 => \N__6087\,
            in3 => \N__5850\,
            lcout => \U712_CHIP_RAM.N_528\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001111111"
        )
    port map (
            in0 => \N__5645\,
            in1 => \N__6252\,
            in2 => \N__6601\,
            in3 => \N__7314\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_482_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100000000"
        )
    port map (
            in0 => \N__6538\,
            in1 => \N__6600\,
            in2 => \N__5620\,
            in3 => \N__8000\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011000100"
        )
    port map (
            in0 => \N__5617\,
            in1 => \N__7990\,
            in2 => \N__5584\,
            in3 => \N__5572\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8780\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6740\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6652\,
            lcout => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.BANK0_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIFS4TD_2_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__5952\,
            in1 => \N__5524\,
            in2 => \N__5509\,
            in3 => \N__5506\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10276\,
            in1 => \_gnd_net_\,
            in2 => \N__5500\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011010001"
        )
    port map (
            in0 => \N__6160\,
            in1 => \N__6146\,
            in2 => \N__8295\,
            in3 => \N__6118\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8780\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000000000"
        )
    port map (
            in0 => \N__7168\,
            in1 => \N__6082\,
            in2 => \N__5977\,
            in3 => \N__5851\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_530_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__6651\,
            in1 => \N__6739\,
            in2 => \N__5839\,
            in3 => \N__5829\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10275\,
            in1 => \_gnd_net_\,
            in2 => \N__5800\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110001010"
        )
    port map (
            in0 => \N__7642\,
            in1 => \N__8184\,
            in2 => \N__7357\,
            in3 => \N__7372\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8785\,
            ce => 'H',
            sr => \N__10217\
        );

    \U712_CHIP_RAM.DBDIR_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__5730\,
            in1 => \N__5785\,
            in2 => \_gnd_net_\,
            in3 => \N__5749\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8785\,
            ce => 'H',
            sr => \N__10217\
        );

    \U712_CHIP_RAM.DBENn_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__9808\,
            in1 => \N__5719\,
            in2 => \_gnd_net_\,
            in3 => \N__5713\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8785\,
            ce => 'H',
            sr => \N__10217\
        );

    \U712_REG_SM.START_RST_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__5707\,
            in1 => \N__6195\,
            in2 => \_gnd_net_\,
            in3 => \N__6289\,
            lcout => \U712_REG_SM.START_RSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8785\,
            ce => 'H',
            sr => \N__10217\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000101000001011"
        )
    port map (
            in0 => \N__6295\,
            in1 => \N__7320\,
            in2 => \N__7042\,
            in3 => \N__7332\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8785\,
            ce => 'H',
            sr => \N__10217\
        );

    \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__6508\,
            in1 => \N__7266\,
            in2 => \_gnd_net_\,
            in3 => \N__6579\,
            lcout => \U712_REG_SM.N_407\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_0_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__7265\,
            in1 => \N__7237\,
            in2 => \_gnd_net_\,
            in3 => \N__6253\,
            lcout => \U712_REG_SM.DS_EN_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_RNO_0_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__6507\,
            in1 => \_gnd_net_\,
            in2 => \N__7273\,
            in3 => \N__6287\,
            lcout => \U712_REG_SM.N_443\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6220\,
            in1 => \N__7268\,
            in2 => \_gnd_net_\,
            in3 => \N__7315\,
            lcout => \U712_REG_SM.STATE_COUNT_srsts_i_i_i_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_1_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__6254\,
            in1 => \N__7267\,
            in2 => \N__6529\,
            in3 => \N__6288\,
            lcout => \U712_REG_SM.N_515\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_2_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__6286\,
            in1 => \N__6577\,
            in2 => \N__6530\,
            in3 => \N__6255\,
            lcout => \U712_REG_SM.un1_STATE_COUNT_4_i_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6506\,
            in1 => \N__6219\,
            in2 => \N__6593\,
            in3 => \N__6205\,
            lcout => \U712_REG_SM.START_RST_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__7264\,
            in1 => \N__6573\,
            in2 => \_gnd_net_\,
            in3 => \N__6505\,
            lcout => \U712_REG_SM.N_480\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101100000001"
        )
    port map (
            in0 => \N__6184\,
            in1 => \N__6178\,
            in2 => \N__6172\,
            in3 => \N__9324\,
            lcout => \DS_ENm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8794\,
            ce => 'H',
            sr => \N__10214\
        );

    \U712_REG_SM.ASn_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__6607\,
            in1 => \N__6580\,
            in2 => \N__6534\,
            in3 => \N__6431\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8794\,
            ce => 'H',
            sr => \N__10214\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__11245\,
            in1 => \N__11324\,
            in2 => \_gnd_net_\,
            in3 => \N__7950\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__7959\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DMA_LATCH_EN_i_i_a2_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__7179\,
            in1 => \N__11329\,
            in2 => \_gnd_net_\,
            in3 => \N__11256\,
            lcout => \N_549\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6373\,
            in2 => \_gnd_net_\,
            in3 => \N__6361\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_11_5_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__6864\,
            ce => 'H',
            sr => \N__6778\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6358\,
            in2 => \_gnd_net_\,
            in3 => \N__6346\,
            lcout => \U712_CHIP_RAM.REFRESH5lto1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__6864\,
            ce => 'H',
            sr => \N__6778\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6343\,
            in2 => \_gnd_net_\,
            in3 => \N__6331\,
            lcout => \U712_CHIP_RAM.REFRESH5lto2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__6864\,
            ce => 'H',
            sr => \N__6778\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6328\,
            in2 => \_gnd_net_\,
            in3 => \N__6316\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__6864\,
            ce => 'H',
            sr => \N__6778\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6312\,
            in2 => \_gnd_net_\,
            in3 => \N__6298\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__6864\,
            ce => 'H',
            sr => \N__6778\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6910\,
            in2 => \_gnd_net_\,
            in3 => \N__6898\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__6864\,
            ce => 'H',
            sr => \N__6778\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6895\,
            in2 => \_gnd_net_\,
            in3 => \N__6883\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__6864\,
            ce => 'H',
            sr => \N__6778\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6877\,
            in2 => \_gnd_net_\,
            in3 => \N__6880\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6864\,
            ce => 'H',
            sr => \N__6778\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9005\,
            in1 => \N__6835\,
            in2 => \_gnd_net_\,
            in3 => \N__6813\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__9147\,
            in1 => \N__9003\,
            in2 => \N__8296\,
            in3 => \N__8353\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => \U712_CHIP_RAM.REFRESH_RST_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__9004\,
            in1 => \N__8354\,
            in2 => \N__6766\,
            in3 => \N__9148\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6763\,
            in2 => \_gnd_net_\,
            in3 => \N__6669\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8775\,
            ce => \N__6613\,
            sr => \N__10222\
        );

    \U712_CYCLE_TERM.RAM_CYCLE_RNO_0_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6977\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6946\,
            lcout => \U712_CYCLE_TERM.N_566\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__6947\,
            in1 => \N__6998\,
            in2 => \_gnd_net_\,
            in3 => \N__6978\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.TACK_EN_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7585\,
            in2 => \N__7048\,
            in3 => \N__8038\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8777\,
            ce => 'H',
            sr => \N__10218\
        );

    \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_0_a2_1_0_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6997\,
            in2 => \_gnd_net_\,
            in3 => \N__6976\,
            lcout => \U712_CYCLE_TERM.N_598\,
            ltout => \U712_CYCLE_TERM.N_598_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010001000110010"
        )
    port map (
            in0 => \N__8089\,
            in1 => \N__8069\,
            in2 => \N__7045\,
            in3 => \N__8050\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8777\,
            ce => 'H',
            sr => \N__10218\
        );

    \U712_REG_SM.REG_TACK_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__7041\,
            in1 => \N__7015\,
            in2 => \N__7003\,
            in3 => \N__6916\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8777\,
            ce => 'H',
            sr => \N__10218\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100110011"
        )
    port map (
            in0 => \N__7002\,
            in1 => \N__7349\,
            in2 => \N__6982\,
            in3 => \N__6948\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_571_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__6949\,
            in1 => \N__7960\,
            in2 => \N__6931\,
            in3 => \N__8185\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8781\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7963\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7371\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8781\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__7316\,
            in1 => \N__7236\,
            in2 => \_gnd_net_\,
            in3 => \N__6927\,
            lcout => \U712_REG_SM.REG_TACK_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7961\,
            in1 => \N__8183\,
            in2 => \_gnd_net_\,
            in3 => \N__7350\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8781\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7962\,
            in2 => \_gnd_net_\,
            in3 => \N__8070\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8781\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNI05SV_3_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7370\,
            in2 => \_gnd_net_\,
            in3 => \N__7348\,
            lcout => \U712_CYCLE_TERM.N_440\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__7949\,
            in1 => \N__7333\,
            in2 => \N__7321\,
            in3 => \N__7272\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8786\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100001111111"
        )
    port map (
            in0 => \N__11325\,
            in1 => \N__11255\,
            in2 => \N__7235\,
            in3 => \N__7180\,
            lcout => \N_483\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__8888\,
            in1 => \N__8364\,
            in2 => \_gnd_net_\,
            in3 => \N__9073\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8759\,
            ce => \N__8667\,
            sr => \N__10243\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000011"
        )
    port map (
            in0 => \N__7675\,
            in1 => \N__9072\,
            in2 => \N__8893\,
            in3 => \N__7492\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8761\,
            ce => \N__8677\,
            sr => \N__10235\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10277\,
            in2 => \_gnd_net_\,
            in3 => \N__7054\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110001111"
        )
    port map (
            in0 => \N__10039\,
            in1 => \N__8867\,
            in2 => \N__9086\,
            in3 => \N__9644\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9160\,
            in2 => \_gnd_net_\,
            in3 => \N__8298\,
            lcout => \U712_CHIP_RAM.N_412\,
            ltout => \U712_CHIP_RAM.N_412_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100000101"
        )
    port map (
            in0 => \N__9075\,
            in1 => \N__9620\,
            in2 => \N__7516\,
            in3 => \N__10038\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9621\,
            in1 => \N__7513\,
            in2 => \_gnd_net_\,
            in3 => \N__9421\,
            lcout => \U712_CHIP_RAM.N_478\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9076\,
            in1 => \N__7486\,
            in2 => \N__9663\,
            in3 => \N__8428\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9643\,
            in2 => \_gnd_net_\,
            in3 => \N__9074\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__7474\,
            in1 => \N__9021\,
            in2 => \N__9659\,
            in3 => \N__9472\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__8874\,
            in1 => \N__8927\,
            in2 => \N__7468\,
            in3 => \N__9880\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8763\,
            ce => \N__8676\,
            sr => \N__10221\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__8875\,
            in1 => \N__8928\,
            in2 => \N__8419\,
            in3 => \N__8191\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8763\,
            ce => \N__8676\,
            sr => \N__10221\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7435\,
            in1 => \N__7401\,
            in2 => \_gnd_net_\,
            in3 => \N__9070\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9071\,
            in1 => \N__9636\,
            in2 => \N__8194\,
            in3 => \N__8443\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_RNI8MQ3_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8182\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNIDG0M2_4_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110100"
        )
    port map (
            in0 => \N__8088\,
            in1 => \N__8077\,
            in2 => \N__8071\,
            in3 => \N__8049\,
            lcout => \U712_CYCLE_TERM.un13_0\,
            ltout => \U712_CYCLE_TERM.un13_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.RAM_CYCLE_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__7924\,
            in1 => \N__7828\,
            in2 => \N__7822\,
            in3 => \N__7620\,
            lcout => \U712_CYCLE_TERM.RAM_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9635\,
            in1 => \N__9069\,
            in2 => \N__7819\,
            in3 => \N__9367\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9738\,
            in2 => \_gnd_net_\,
            in3 => \N__7807\,
            lcout => \U712_CHIP_RAM.N_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7710\,
            in1 => \N__9634\,
            in2 => \_gnd_net_\,
            in3 => \N__9976\,
            lcout => \U712_CHIP_RAM.N_455\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.RAM_CYCLE_RNILITE_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__7652\,
            in1 => \N__7621\,
            in2 => \_gnd_net_\,
            in3 => \N__7586\,
            lcout => \U712_CYCLE_TERM_TCIn_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000110000"
        )
    port map (
            in0 => \N__11005\,
            in1 => \N__11158\,
            in2 => \N__9667\,
            in3 => \N__9228\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_563_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_56_i_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001101"
        )
    port map (
            in0 => \N__9781\,
            in1 => \N__9834\,
            in2 => \N__8407\,
            in3 => \N__11320\,
            lcout => \N_56_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_LDSn_i_0_0_o2_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11053\,
            in2 => \_gnd_net_\,
            in3 => \N__10869\,
            lcout => \U712_BYTE_ENABLE.N_410\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WEn_LC_13_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8302\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8760\,
            ce => 'H',
            sr => \N__10257\
        );

    \U712_CHIP_RAM.CRCSn_LC_13_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8365\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8760\,
            ce => 'H',
            sr => \N__10257\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__9168\,
            in1 => \N__9050\,
            in2 => \_gnd_net_\,
            in3 => \N__8297\,
            lcout => \U712_CHIP_RAM.CMA_5_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9051\,
            in1 => \N__8245\,
            in2 => \N__9664\,
            in3 => \N__8437\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8236\,
            in1 => \N__8230\,
            in2 => \_gnd_net_\,
            in3 => \N__8224\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8764\,
            ce => \N__8675\,
            sr => \N__10237\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__8921\,
            in1 => \N__10684\,
            in2 => \N__8890\,
            in3 => \N__8617\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8764\,
            ce => \N__8675\,
            sr => \N__10237\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__8523\,
            in1 => \N__8590\,
            in2 => \N__9658\,
            in3 => \N__10630\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8764\,
            ce => \N__8675\,
            sr => \N__10237\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__8922\,
            in1 => \N__9478\,
            in2 => \N__8891\,
            in3 => \N__8548\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8764\,
            ce => \N__8675\,
            sr => \N__10237\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__8527\,
            in1 => \N__8512\,
            in2 => \N__9665\,
            in3 => \N__10372\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8767\,
            ce => \N__8674\,
            sr => \N__10232\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__8926\,
            in1 => \N__9484\,
            in2 => \N__8892\,
            in3 => \N__8473\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8767\,
            ce => \N__8674\,
            sr => \N__10232\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9460\,
            in1 => \N__9407\,
            in2 => \_gnd_net_\,
            in3 => \N__10594\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__10316\,
            sr => \N__10223\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10596\,
            in1 => \N__10428\,
            in2 => \_gnd_net_\,
            in3 => \N__10675\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__10316\,
            sr => \N__10223\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10595\,
            in1 => \N__10731\,
            in2 => \_gnd_net_\,
            in3 => \N__10674\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__10316\,
            sr => \N__10223\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10587\,
            in1 => \N__9456\,
            in2 => \_gnd_net_\,
            in3 => \N__10018\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10355\,
            ce => \N__10314\,
            sr => \N__10219\
        );

    \U712_CHIP_RAM.DMA_A20_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__9289\,
            in1 => \N__10421\,
            in2 => \N__10591\,
            in3 => \N__9270\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A20C_net\,
            ce => 'H',
            sr => \N__10216\
        );

    \U712_BYTE_ENABLE.N_58_i_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__9835\,
            in1 => \N__11316\,
            in2 => \N__9211\,
            in3 => \N__9783\,
            lcout => \N_58_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100000000"
        )
    port map (
            in0 => \N__11018\,
            in1 => \N__11157\,
            in2 => \N__9232\,
            in3 => \N__9666\,
            lcout => \U712_BYTE_ENABLE.N_559\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_129_i_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011100000"
        )
    port map (
            in0 => \N__11006\,
            in1 => \N__11065\,
            in2 => \N__10927\,
            in3 => \N__10841\,
            lcout => \N_129_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CASn_LC_14_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9088\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8762\,
            ce => 'H',
            sr => \N__10260\
        );

    \U712_CHIP_RAM.RASn_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9169\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8765\,
            ce => 'H',
            sr => \N__10252\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9648\,
            in1 => \N__9100\,
            in2 => \N__9087\,
            in3 => \N__10090\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__8929\,
            in1 => \N__8889\,
            in2 => \N__8827\,
            in3 => \N__9490\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8768\,
            ce => \N__8663\,
            sr => \N__10245\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10617\,
            in1 => \N__9409\,
            in2 => \_gnd_net_\,
            in3 => \N__10068\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10357\,
            ce => \N__10321\,
            sr => \N__10238\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__9408\,
            in1 => \N__9455\,
            in2 => \_gnd_net_\,
            in3 => \N__10616\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10357\,
            ce => \N__10321\,
            sr => \N__10238\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10673\,
            in1 => \N__10735\,
            in2 => \_gnd_net_\,
            in3 => \N__10618\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10357\,
            ce => \N__10321\,
            sr => \N__10238\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9955\,
            in1 => \N__10020\,
            in2 => \_gnd_net_\,
            in3 => \N__10530\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__10319\,
            sr => \N__10233\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__10531\,
            in1 => \_gnd_net_\,
            in2 => \N__10024\,
            in3 => \N__9448\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__10319\,
            sr => \N__10233\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10067\,
            in1 => \N__9398\,
            in2 => \_gnd_net_\,
            in3 => \N__10555\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            ce => \N__10317\,
            sr => \N__10224\
        );

    \U712_BYTE_ENABLE.un1_UDSn_i_0_0_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100011111111"
        )
    port map (
            in0 => \N__10843\,
            in1 => \N__11086\,
            in2 => \N__10929\,
            in3 => \N__9340\,
            lcout => \un1_UDSn_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_LDSn_i_0_0_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011111111"
        )
    port map (
            in0 => \N__10842\,
            in1 => \N__11085\,
            in2 => \N__10928\,
            in3 => \N__9339\,
            lcout => \un1_LDSn_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10615\,
            in1 => \N__10786\,
            in2 => \_gnd_net_\,
            in3 => \N__10730\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__10324\,
            sr => \N__10253\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10614\,
            in1 => \N__10084\,
            in2 => \_gnd_net_\,
            in3 => \N__10778\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__10323\,
            sr => \N__10246\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10521\,
            in1 => \N__10080\,
            in2 => \_gnd_net_\,
            in3 => \N__10769\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10353\,
            ce => \N__10322\,
            sr => \N__10239\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10019\,
            in1 => \N__9954\,
            in2 => \_gnd_net_\,
            in3 => \N__10599\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10352\,
            ce => \N__10320\,
            sr => \N__10234\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10598\,
            in1 => \N__9913\,
            in2 => \_gnd_net_\,
            in3 => \N__9946\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10318\,
            sr => \N__10225\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__9953\,
            in1 => \N__9909\,
            in2 => \_gnd_net_\,
            in3 => \N__10597\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10351\,
            ce => \N__10315\,
            sr => \N__10220\
        );

    \U712_BYTE_ENABLE.N_57_i_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100011"
        )
    port map (
            in0 => \N__11224\,
            in1 => \N__11167\,
            in2 => \N__9787\,
            in3 => \N__9845\,
            lcout => \N_57_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_59_i_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__11257\,
            in1 => \N__9673\,
            in2 => \N__9850\,
            in3 => \N__9782\,
            lcout => \N_59_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100000000"
        )
    port map (
            in0 => \N__11084\,
            in1 => \N__11020\,
            in2 => \N__11156\,
            in3 => \N__9629\,
            lcout => \U712_BYTE_ENABLE.N_557\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100000000"
        )
    port map (
            in0 => \N__11083\,
            in1 => \N__11019\,
            in2 => \N__11155\,
            in3 => \N__9628\,
            lcout => \U712_BYTE_ENABLE.N_561\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LLBE_i_o2_0_x2_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10942\,
            in2 => \_gnd_net_\,
            in3 => \N__10870\,
            lcout => \U712_BYTE_ENABLE.N_397_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_130_i_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111010000"
        )
    port map (
            in0 => \N__11012\,
            in1 => \N__11089\,
            in2 => \N__10868\,
            in3 => \N__10936\,
            lcout => \N_130_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_127_i_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011010000"
        )
    port map (
            in0 => \N__11087\,
            in1 => \N__11010\,
            in2 => \N__10940\,
            in3 => \N__10857\,
            lcout => \N_127_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_128_i_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001101110000"
        )
    port map (
            in0 => \N__11088\,
            in1 => \N__11011\,
            in2 => \N__10941\,
            in3 => \N__10858\,
            lcout => \N_128_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10593\,
            in1 => \N__10785\,
            in2 => \_gnd_net_\,
            in3 => \N__10720\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10356\,
            ce => \N__10327\,
            sr => \N__10258\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10592\,
            in1 => \N__10429\,
            in2 => \_gnd_net_\,
            in3 => \N__10667\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10354\,
            ce => \N__10325\,
            sr => \N__10254\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10569\,
            in1 => \N__10438\,
            in2 => \_gnd_net_\,
            in3 => \N__10403\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10350\,
            ce => \N__10326\,
            sr => \N__10255\
        );

    \U712_BUFFERS.un1_DRDENn_0_a2_LC_24_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__10126\,
            in1 => \N__11300\,
            in2 => \_gnd_net_\,
            in3 => \N__11218\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jul 2 2025 17:00:31

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    DA : out std_logic_vector(2 downto 0);
    A : in std_logic_vector(20 downto 0);
    TBIn : out std_logic;
    RAMSPACEn : in std_logic;
    DBRn : in std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    PRnW : out std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    BLSn : out std_logic;
    TCIn : out std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__13257\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13248\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13239\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13230\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13219\ : std_logic;
signal \N__13212\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13203\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13192\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13149\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13084\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13048\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__12996\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12976\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12931\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12913\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12904\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12895\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12877\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12868\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12841\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12814\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12778\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12769\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12760\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12733\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12589\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12037\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10629\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9753\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7657\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7347\ : std_logic;
signal \N__7344\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7275\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6996\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \bfn_6_7_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_3\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_7\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_a2_1_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_165_i_i_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \U712_CHIP_RAM.N_90_i_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_298_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_300_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_310\ : std_logic;
signal \U712_CHIP_RAM.N_310_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_313\ : std_logic;
signal \U712_CHIP_RAM.N_389\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3_cascade_\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\ : std_logic;
signal \DBR_SYNC_i_1\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a3_0_a2_0\ : std_logic;
signal \N_178_i\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0\ : std_logic;
signal \N_176_i\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER19\ : std_logic;
signal \U712_CHIP_RAM.N_464_cascade_\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0\ : std_logic;
signal \U712_CHIP_RAM.N_390\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_o2_0_0\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.N_90_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \N_188_i\ : std_logic;
signal \U712_CHIP_RAM.N_302\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3\ : std_logic;
signal \U712_CHIP_RAM.N_455\ : std_logic;
signal \U712_CHIP_RAM.N_417_cascade_\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto7_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lt7\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_419\ : std_logic;
signal \U712_BYTE_ENABLE.N_326\ : std_logic;
signal \U712_BYTE_ENABLE.N_323\ : std_logic;
signal \U712_BYTE_ENABLE.N_324\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U712_CHIP_RAM.N_463_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.N_385_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_384\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_461\ : std_logic;
signal \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERlde_0_a3_0_0_a2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERlde_0_a3_0_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_533_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_370\ : std_logic;
signal \U712_CHIP_RAM.N_391_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.N_295_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_546\ : std_logic;
signal \U712_CHIP_RAM.N_464\ : std_logic;
signal \U712_CHIP_RAM.N_465\ : std_logic;
signal \U712_CHIP_RAM.N_465_cascade_\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0\ : std_logic;
signal \U712_CHIP_RAM.DBENn_8_0_0\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \CLK40_PLL_i_i\ : std_logic;
signal \N_167_i\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\ : std_logic;
signal \LATCH_CLK_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_a2_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_533\ : std_logic;
signal \U712_CHIP_RAM.N_296_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_550\ : std_logic;
signal \U712_CHIP_RAM.N_463\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.N_442_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_441\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_8_iv_i_a2_1\ : std_logic;
signal \U712_CHIP_RAM.N_295\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_551\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_458\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_0_0_0_a2_1\ : std_logic;
signal \U712_CHIP_RAM.N_428\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_300\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_438\ : std_logic;
signal \U712_CHIP_RAM.N_469\ : std_logic;
signal \U712_CHIP_RAM.N_438_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_a2_1\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_a2_2\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \U712_CYCLE_TERM.N_321\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \A_c_9\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_305_cascade_\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0Z0Z_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_325\ : std_logic;
signal \N_186_i\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CYCLE_TERM.N_450_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ1Z_2\ : std_logic;
signal \CLK40_PLL_i\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_5\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_6\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_4\ : std_logic;
signal \U712_REG_SM.N_320_cascade_\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA25_0_i\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_346\ : std_logic;
signal \U712_CHIP_RAM.N_352\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\ : std_logic;
signal \N_169_i\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_REG_SM.N_397_cascade_\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_3\ : std_logic;
signal \U712_REG_SM.N_548\ : std_logic;
signal \U712_REG_SM.N_319_cascade_\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_5_iv_0_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_409\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \U712_REG_SM.STATE_COUNTsr_0\ : std_logic;
signal \U712_REG_SM.N_328\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_412_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_3\ : std_logic;
signal \U712_REG_SM.N_360_cascade_\ : std_logic;
signal \U712_REG_SM.N_320\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\ : std_logic;
signal \U712_REG_SM.START_RSTZ0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_7\ : std_logic;
signal \U712_REG_SM.N_319\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_318_cascade_\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \BLSn_c\ : std_logic;
signal \U712_REG_SM.REGENn_e_1\ : std_logic;
signal \N_326_i\ : std_logic;
signal \N_325_i\ : std_logic;
signal \N_323_i\ : std_logic;
signal \A_c_1\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \N_324_i\ : std_logic;
signal \WEn_c\ : std_logic;
signal \U712_CHIP_RAM.N_305\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA25_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_i_0_9\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_8\ : std_logic;
signal \U712_REG_SM.N_400\ : std_logic;
signal \UDSn_c\ : std_logic;
signal \U712_REG_SM.WRITE_CYCLEZ0\ : std_logic;
signal \PRnW_c\ : std_logic;
signal \U712_REG_SM.N_398\ : std_logic;
signal \LDSn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \RASn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_152\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.N_152_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_0\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \RnW_c\ : std_logic;
signal \DMA_WRITE_CYCLE\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \N_362\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \DA_wire\ : std_logic_vector(2 downto 0);
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \PRnW_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \BLSn_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    TBIn <= \TBIn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    ASn <= \ASn_wire\;
    DA <= \DA_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    TCIn <= \TCIn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    PRnW <= \PRnW_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    \C3_wire\ <= C3;
    BLSn <= \BLSn_wire\;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL_i\,
            REFERENCECLK => \N__4445\,
            RESETB => \N__6377\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13257\,
            DIN => \N__13256\,
            DOUT => \N__13255\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13257\,
            PADOUT => \N__13256\,
            PADIN => \N__13255\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7040\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13248\,
            DIN => \N__13247\,
            DOUT => \N__13246\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13248\,
            PADOUT => \N__13247\,
            PADIN => \N__13246\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13239\,
            DIN => \N__13238\,
            DOUT => \N__13237\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13239\,
            PADOUT => \N__13238\,
            PADIN => \N__13237\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10454\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13230\,
            DIN => \N__13229\,
            DOUT => \N__13228\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13230\,
            PADOUT => \N__13229\,
            PADIN => \N__13228\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12374\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13221\,
            DIN => \N__13220\,
            DOUT => \N__13219\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13221\,
            PADOUT => \N__13220\,
            PADIN => \N__13219\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13212\,
            DIN => \N__13211\,
            DOUT => \N__13210\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13212\,
            PADOUT => \N__13211\,
            PADIN => \N__13210\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13203\,
            DIN => \N__13202\,
            DOUT => \N__13201\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13203\,
            PADOUT => \N__13202\,
            PADIN => \N__13201\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13194\,
            DIN => \N__13193\,
            DOUT => \N__13192\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13194\,
            PADOUT => \N__13193\,
            PADIN => \N__13192\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13185\,
            DIN => \N__13184\,
            DOUT => \N__13183\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13185\,
            PADOUT => \N__13184\,
            PADIN => \N__13183\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13176\,
            DIN => \N__13175\,
            DOUT => \N__13174\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13176\,
            PADOUT => \N__13175\,
            PADIN => \N__13174\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13167\,
            DIN => \N__13166\,
            DOUT => \N__13165\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13167\,
            PADOUT => \N__13166\,
            PADIN => \N__13165\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13158\,
            DIN => \N__13157\,
            DOUT => \N__13156\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13158\,
            PADOUT => \N__13157\,
            PADIN => \N__13156\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8420\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13149\,
            DIN => \N__13148\,
            DOUT => \N__13147\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13149\,
            PADOUT => \N__13148\,
            PADIN => \N__13147\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8786\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13140\,
            DIN => \N__13139\,
            DOUT => \N__13138\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13140\,
            PADOUT => \N__13139\,
            PADIN => \N__13138\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13131\,
            DIN => \N__13130\,
            DOUT => \N__13129\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13131\,
            PADOUT => \N__13130\,
            PADIN => \N__13129\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13122\,
            DIN => \N__13121\,
            DOUT => \N__13120\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13122\,
            PADOUT => \N__13121\,
            PADIN => \N__13120\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13113\,
            DIN => \N__13112\,
            DOUT => \N__13111\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13113\,
            PADOUT => \N__13112\,
            PADIN => \N__13111\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4691\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13104\,
            DIN => \N__13103\,
            DOUT => \N__13102\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13104\,
            PADOUT => \N__13103\,
            PADIN => \N__13102\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13095\,
            DIN => \N__13094\,
            DOUT => \N__13093\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13095\,
            PADOUT => \N__13094\,
            PADIN => \N__13093\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13086\,
            DIN => \N__13085\,
            DOUT => \N__13084\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13086\,
            PADOUT => \N__13085\,
            PADIN => \N__13084\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8549\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13077\,
            DIN => \N__13076\,
            DOUT => \N__13075\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13077\,
            PADOUT => \N__13076\,
            PADIN => \N__13075\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13068\,
            DIN => \N__13067\,
            DOUT => \N__13066\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13068\,
            PADOUT => \N__13067\,
            PADIN => \N__13066\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12140\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13059\,
            DIN => \N__13058\,
            DOUT => \N__13057\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13059\,
            PADOUT => \N__13058\,
            PADIN => \N__13057\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13050\,
            DIN => \N__13049\,
            DOUT => \N__13048\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13050\,
            PADOUT => \N__13049\,
            PADIN => \N__13048\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9782\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13041\,
            DIN => \N__13040\,
            DOUT => \N__13039\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13041\,
            PADOUT => \N__13040\,
            PADIN => \N__13039\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6921\,
            DIN0 => OPEN,
            DOUT0 => \N__7647\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13032\,
            DIN => \N__13031\,
            DOUT => \N__13030\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13032\,
            PADOUT => \N__13031\,
            PADIN => \N__13030\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13023\,
            DIN => \N__13022\,
            DOUT => \N__13021\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13023\,
            PADOUT => \N__13022\,
            PADIN => \N__13021\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13014\,
            DIN => \N__13013\,
            DOUT => \N__13012\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13014\,
            PADOUT => \N__13013\,
            PADIN => \N__13012\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13005\,
            DIN => \N__13004\,
            DOUT => \N__13003\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13005\,
            PADOUT => \N__13004\,
            PADIN => \N__13003\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12996\,
            DIN => \N__12995\,
            DOUT => \N__12994\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12996\,
            PADOUT => \N__12995\,
            PADIN => \N__12994\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12987\,
            DIN => \N__12986\,
            DOUT => \N__12985\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12987\,
            PADOUT => \N__12986\,
            PADIN => \N__12985\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5924\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12978\,
            DIN => \N__12977\,
            DOUT => \N__12976\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12978\,
            PADOUT => \N__12977\,
            PADIN => \N__12976\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12969\,
            DIN => \N__12968\,
            DOUT => \N__12967\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12969\,
            PADOUT => \N__12968\,
            PADIN => \N__12967\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12960\,
            DIN => \N__12959\,
            DOUT => \N__12958\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12960\,
            PADOUT => \N__12959\,
            PADIN => \N__12958\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12951\,
            DIN => \N__12950\,
            DOUT => \N__12949\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12951\,
            PADOUT => \N__12950\,
            PADIN => \N__12949\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12942\,
            DIN => \N__12941\,
            DOUT => \N__12940\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12942\,
            PADOUT => \N__12941\,
            PADIN => \N__12940\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12933\,
            DIN => \N__12932\,
            DOUT => \N__12931\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12933\,
            PADOUT => \N__12932\,
            PADIN => \N__12931\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10388\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12924\,
            DIN => \N__12923\,
            DOUT => \N__12922\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12924\,
            PADOUT => \N__12923\,
            PADIN => \N__12922\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12915\,
            DIN => \N__12914\,
            DOUT => \N__12913\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12915\,
            PADOUT => \N__12914\,
            PADIN => \N__12913\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12906\,
            DIN => \N__12905\,
            DOUT => \N__12904\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12906\,
            PADOUT => \N__12905\,
            PADIN => \N__12904\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12218\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12897\,
            DIN => \N__12896\,
            DOUT => \N__12895\,
            PACKAGEPIN => \DA_wire\(0)
        );

    \DA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12897\,
            PADOUT => \N__12896\,
            PADIN => \N__12895\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7532\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12888\,
            DIN => \N__12887\,
            DOUT => \N__12886\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12888\,
            PADOUT => \N__12887\,
            PADIN => \N__12886\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12879\,
            DIN => \N__12878\,
            DOUT => \N__12877\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12879\,
            PADOUT => \N__12878\,
            PADIN => \N__12877\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8531\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12870\,
            DIN => \N__12869\,
            DOUT => \N__12868\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12870\,
            PADOUT => \N__12869\,
            PADIN => \N__12868\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8447\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12861\,
            DIN => \N__12860\,
            DOUT => \N__12859\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12861\,
            PADOUT => \N__12860\,
            PADIN => \N__12859\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8840\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12852\,
            DIN => \N__12851\,
            DOUT => \N__12850\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12852\,
            PADOUT => \N__12851\,
            PADIN => \N__12850\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12843\,
            DIN => \N__12842\,
            DOUT => \N__12841\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12843\,
            PADOUT => \N__12842\,
            PADIN => \N__12841\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7769\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12834\,
            DIN => \N__12833\,
            DOUT => \N__12832\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12834\,
            PADOUT => \N__12833\,
            PADIN => \N__12832\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6928\,
            DIN0 => OPEN,
            DOUT0 => \N__7651\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12825\,
            DIN => \N__12824\,
            DOUT => \N__12823\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12825\,
            PADOUT => \N__12824\,
            PADIN => \N__12823\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9413\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12816\,
            DIN => \N__12815\,
            DOUT => \N__12814\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12816\,
            PADOUT => \N__12815\,
            PADIN => \N__12814\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6002\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12807\,
            DIN => \N__12806\,
            DOUT => \N__12805\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12807\,
            PADOUT => \N__12806\,
            PADIN => \N__12805\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4952\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12798\,
            DIN => \N__12797\,
            DOUT => \N__12796\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12798\,
            PADOUT => \N__12797\,
            PADIN => \N__12796\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12789\,
            DIN => \N__12788\,
            DOUT => \N__12787\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12789\,
            PADOUT => \N__12788\,
            PADIN => \N__12787\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12780\,
            DIN => \N__12779\,
            DOUT => \N__12778\,
            PACKAGEPIN => \DA_wire\(2)
        );

    \DA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12780\,
            PADOUT => \N__12779\,
            PADIN => \N__12778\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6347\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12771\,
            DIN => \N__12770\,
            DOUT => \N__12769\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12771\,
            PADOUT => \N__12770\,
            PADIN => \N__12769\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12762\,
            DIN => \N__12761\,
            DOUT => \N__12760\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12762\,
            PADOUT => \N__12761\,
            PADIN => \N__12760\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12753\,
            DIN => \N__12752\,
            DOUT => \N__12751\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12753\,
            PADOUT => \N__12752\,
            PADIN => \N__12751\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7934\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12744\,
            DIN => \N__12743\,
            DOUT => \N__12742\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12744\,
            PADOUT => \N__12743\,
            PADIN => \N__12742\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9800\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12735\,
            DIN => \N__12734\,
            DOUT => \N__12733\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12735\,
            PADOUT => \N__12734\,
            PADIN => \N__12733\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12726\,
            DIN => \N__12725\,
            DOUT => \N__12724\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12726\,
            PADOUT => \N__12725\,
            PADIN => \N__12724\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5177\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12717\,
            DIN => \N__12716\,
            DOUT => \N__12715\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12717\,
            PADOUT => \N__12716\,
            PADIN => \N__12715\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6929\,
            DIN0 => OPEN,
            DOUT0 => \N__7652\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12708\,
            DIN => \N__12707\,
            DOUT => \N__12706\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12708\,
            PADOUT => \N__12707\,
            PADIN => \N__12706\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6860\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12699\,
            DIN => \N__12698\,
            DOUT => \N__12697\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12699\,
            PADOUT => \N__12698\,
            PADIN => \N__12697\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12690\,
            DIN => \N__12689\,
            DOUT => \N__12688\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12690\,
            PADOUT => \N__12689\,
            PADIN => \N__12688\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12681\,
            DIN => \N__12680\,
            DOUT => \N__12679\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12681\,
            PADOUT => \N__12680\,
            PADIN => \N__12679\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8480\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12672\,
            DIN => \N__12671\,
            DOUT => \N__12670\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12672\,
            PADOUT => \N__12671\,
            PADIN => \N__12670\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12663\,
            DIN => \N__12662\,
            DOUT => \N__12661\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12663\,
            PADOUT => \N__12662\,
            PADIN => \N__12661\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12654\,
            DIN => \N__12653\,
            DOUT => \N__12652\,
            PACKAGEPIN => \DA_wire\(1)
        );

    \DA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12654\,
            PADOUT => \N__12653\,
            PADIN => \N__12652\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7493\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12645\,
            DIN => \N__12644\,
            DOUT => \N__12643\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12645\,
            PADOUT => \N__12644\,
            PADIN => \N__12643\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12636\,
            DIN => \N__12635\,
            DOUT => \N__12634\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12636\,
            PADOUT => \N__12635\,
            PADIN => \N__12634\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12627\,
            DIN => \N__12626\,
            DOUT => \N__12625\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12627\,
            PADOUT => \N__12626\,
            PADIN => \N__12625\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8177\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12618\,
            DIN => \N__12617\,
            DOUT => \N__12616\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12618\,
            PADOUT => \N__12617\,
            PADIN => \N__12616\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9914\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12609\,
            DIN => \N__12608\,
            DOUT => \N__12607\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12609\,
            PADOUT => \N__12608\,
            PADIN => \N__12607\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9431\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12600\,
            DIN => \N__12599\,
            DOUT => \N__12598\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12600\,
            PADOUT => \N__12599\,
            PADIN => \N__12598\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5885\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12591\,
            DIN => \N__12590\,
            DOUT => \N__12589\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12591\,
            PADOUT => \N__12590\,
            PADIN => \N__12589\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12582\,
            DIN => \N__12581\,
            DOUT => \N__12580\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12582\,
            PADOUT => \N__12581\,
            PADIN => \N__12580\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12573\,
            DIN => \N__12572\,
            DOUT => \N__12571\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12573\,
            PADOUT => \N__12572\,
            PADIN => \N__12571\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8507\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12564\,
            DIN => \N__12563\,
            DOUT => \N__12562\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12564\,
            PADOUT => \N__12563\,
            PADIN => \N__12562\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12555\,
            DIN => \N__12554\,
            DOUT => \N__12553\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12555\,
            PADOUT => \N__12554\,
            PADIN => \N__12553\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12546\,
            DIN => \N__12545\,
            DOUT => \N__12544\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12546\,
            PADOUT => \N__12545\,
            PADIN => \N__12544\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6287\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12537\,
            DIN => \N__12536\,
            DOUT => \N__12535\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12537\,
            PADOUT => \N__12536\,
            PADIN => \N__12535\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9827\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12528\,
            DIN => \N__12527\,
            DOUT => \N__12526\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12528\,
            PADOUT => \N__12527\,
            PADIN => \N__12526\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5975\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PRnW_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12519\,
            DIN => \N__12518\,
            DOUT => \N__12517\,
            PACKAGEPIN => \PRnW_wire\
        );

    \PRnW_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12519\,
            PADOUT => \N__12518\,
            PADIN => \N__12517\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9857\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12510\,
            DIN => \N__12509\,
            DOUT => \N__12508\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12510\,
            PADOUT => \N__12509\,
            PADIN => \N__12508\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12501\,
            DIN => \N__12500\,
            DOUT => \N__12499\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12501\,
            PADOUT => \N__12500\,
            PADIN => \N__12499\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5974\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12492\,
            DIN => \N__12491\,
            DOUT => \N__12490\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12492\,
            PADOUT => \N__12491\,
            PADIN => \N__12490\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4484\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12483\,
            DIN => \N__12482\,
            DOUT => \N__12481\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12483\,
            PADOUT => \N__12482\,
            PADIN => \N__12481\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9272\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12474\,
            DIN => \N__12473\,
            DOUT => \N__12472\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12474\,
            PADOUT => \N__12473\,
            PADIN => \N__12472\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12465\,
            DIN => \N__12464\,
            DOUT => \N__12463\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12465\,
            PADOUT => \N__12464\,
            PADIN => \N__12463\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12456\,
            DIN => \N__12455\,
            DOUT => \N__12454\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12456\,
            PADOUT => \N__12455\,
            PADIN => \N__12454\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BLSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12447\,
            DIN => \N__12446\,
            DOUT => \N__12445\,
            PACKAGEPIN => \BLSn_wire\
        );

    \BLSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12447\,
            PADOUT => \N__12446\,
            PADIN => \N__12445\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8830\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12438\,
            DIN => \N__12437\,
            DOUT => \N__12436\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12438\,
            PADOUT => \N__12437\,
            PADIN => \N__12436\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12429\,
            DIN => \N__12428\,
            DOUT => \N__12427\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12429\,
            PADOUT => \N__12428\,
            PADIN => \N__12427\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5949\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12420\,
            DIN => \N__12419\,
            DOUT => \N__12418\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12420\,
            PADOUT => \N__12419\,
            PADIN => \N__12418\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8111\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12411\,
            DIN => \N__12410\,
            DOUT => \N__12409\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12411\,
            PADOUT => \N__12410\,
            PADIN => \N__12409\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5372\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12402\,
            DIN => \N__12401\,
            DOUT => \N__12400\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12402\,
            PADOUT => \N__12401\,
            PADIN => \N__12400\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8750\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12393\,
            DIN => \N__12392\,
            DOUT => \N__12391\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12393\,
            PADOUT => \N__12392\,
            PADIN => \N__12391\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__3032\ : IoInMux
    port map (
            O => \N__12374\,
            I => \N__12371\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__12371\,
            I => \N__12368\
        );

    \I__3030\ : Span4Mux_s3_h
    port map (
            O => \N__12368\,
            I => \N__12365\
        );

    \I__3029\ : Span4Mux_v
    port map (
            O => \N__12365\,
            I => \N__12362\
        );

    \I__3028\ : Odrv4
    port map (
            O => \N__12362\,
            I => \N_362\
        );

    \I__3027\ : CascadeMux
    port map (
            O => \N__12359\,
            I => \N__12354\
        );

    \I__3026\ : InMux
    port map (
            O => \N__12358\,
            I => \N__12351\
        );

    \I__3025\ : InMux
    port map (
            O => \N__12357\,
            I => \N__12345\
        );

    \I__3024\ : InMux
    port map (
            O => \N__12354\,
            I => \N__12345\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__12351\,
            I => \N__12342\
        );

    \I__3022\ : InMux
    port map (
            O => \N__12350\,
            I => \N__12339\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__12345\,
            I => \U712_REG_SM.N_152\
        );

    \I__3020\ : Odrv4
    port map (
            O => \N__12342\,
            I => \U712_REG_SM.N_152\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__12339\,
            I => \U712_REG_SM.N_152\
        );

    \I__3018\ : CascadeMux
    port map (
            O => \N__12332\,
            I => \N__12326\
        );

    \I__3017\ : InMux
    port map (
            O => \N__12331\,
            I => \N__12321\
        );

    \I__3016\ : InMux
    port map (
            O => \N__12330\,
            I => \N__12315\
        );

    \I__3015\ : CascadeMux
    port map (
            O => \N__12329\,
            I => \N__12311\
        );

    \I__3014\ : InMux
    port map (
            O => \N__12326\,
            I => \N__12308\
        );

    \I__3013\ : CascadeMux
    port map (
            O => \N__12325\,
            I => \N__12301\
        );

    \I__3012\ : CascadeMux
    port map (
            O => \N__12324\,
            I => \N__12298\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__12321\,
            I => \N__12294\
        );

    \I__3010\ : InMux
    port map (
            O => \N__12320\,
            I => \N__12291\
        );

    \I__3009\ : InMux
    port map (
            O => \N__12319\,
            I => \N__12286\
        );

    \I__3008\ : InMux
    port map (
            O => \N__12318\,
            I => \N__12286\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__12315\,
            I => \N__12283\
        );

    \I__3006\ : InMux
    port map (
            O => \N__12314\,
            I => \N__12278\
        );

    \I__3005\ : InMux
    port map (
            O => \N__12311\,
            I => \N__12278\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__12308\,
            I => \N__12275\
        );

    \I__3003\ : InMux
    port map (
            O => \N__12307\,
            I => \N__12268\
        );

    \I__3002\ : InMux
    port map (
            O => \N__12306\,
            I => \N__12268\
        );

    \I__3001\ : InMux
    port map (
            O => \N__12305\,
            I => \N__12268\
        );

    \I__3000\ : InMux
    port map (
            O => \N__12304\,
            I => \N__12265\
        );

    \I__2999\ : InMux
    port map (
            O => \N__12301\,
            I => \N__12262\
        );

    \I__2998\ : InMux
    port map (
            O => \N__12298\,
            I => \N__12257\
        );

    \I__2997\ : InMux
    port map (
            O => \N__12297\,
            I => \N__12257\
        );

    \I__2996\ : Span4Mux_v
    port map (
            O => \N__12294\,
            I => \N__12252\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__12291\,
            I => \N__12252\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__12286\,
            I => \N__12249\
        );

    \I__2993\ : Span4Mux_v
    port map (
            O => \N__12283\,
            I => \N__12246\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__12278\,
            I => \N__12243\
        );

    \I__2991\ : Span4Mux_h
    port map (
            O => \N__12275\,
            I => \N__12232\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__12268\,
            I => \N__12232\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__12265\,
            I => \N__12232\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__12262\,
            I => \N__12232\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__12257\,
            I => \N__12232\
        );

    \I__2986\ : Span4Mux_h
    port map (
            O => \N__12252\,
            I => \N__12229\
        );

    \I__2985\ : Odrv4
    port map (
            O => \N__12249\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2984\ : Odrv4
    port map (
            O => \N__12246\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2983\ : Odrv4
    port map (
            O => \N__12243\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2982\ : Odrv4
    port map (
            O => \N__12232\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2981\ : Odrv4
    port map (
            O => \N__12229\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__2980\ : IoInMux
    port map (
            O => \N__12218\,
            I => \N__12215\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__12215\,
            I => \N__12212\
        );

    \I__2978\ : Span4Mux_s3_v
    port map (
            O => \N__12212\,
            I => \N__12209\
        );

    \I__2977\ : Span4Mux_v
    port map (
            O => \N__12209\,
            I => \N__12206\
        );

    \I__2976\ : Span4Mux_v
    port map (
            O => \N__12206\,
            I => \N__12203\
        );

    \I__2975\ : Sp12to4
    port map (
            O => \N__12203\,
            I => \N__12200\
        );

    \I__2974\ : Odrv12
    port map (
            O => \N__12200\,
            I => \ASn_c\
        );

    \I__2973\ : CEMux
    port map (
            O => \N__12197\,
            I => \N__12194\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__12194\,
            I => \N__12191\
        );

    \I__2971\ : Span4Mux_h
    port map (
            O => \N__12191\,
            I => \N__12188\
        );

    \I__2970\ : Odrv4
    port map (
            O => \N__12188\,
            I => \U712_REG_SM.N_152_0\
        );

    \I__2969\ : InMux
    port map (
            O => \N__12185\,
            I => \N__12181\
        );

    \I__2968\ : InMux
    port map (
            O => \N__12184\,
            I => \N__12178\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__12181\,
            I => \N__12175\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__12178\,
            I => \N__12170\
        );

    \I__2965\ : Span4Mux_h
    port map (
            O => \N__12175\,
            I => \N__12167\
        );

    \I__2964\ : CascadeMux
    port map (
            O => \N__12174\,
            I => \N__12163\
        );

    \I__2963\ : InMux
    port map (
            O => \N__12173\,
            I => \N__12160\
        );

    \I__2962\ : Span4Mux_h
    port map (
            O => \N__12170\,
            I => \N__12155\
        );

    \I__2961\ : Span4Mux_h
    port map (
            O => \N__12167\,
            I => \N__12155\
        );

    \I__2960\ : InMux
    port map (
            O => \N__12166\,
            I => \N__12152\
        );

    \I__2959\ : InMux
    port map (
            O => \N__12163\,
            I => \N__12149\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__12160\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2957\ : Odrv4
    port map (
            O => \N__12155\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__12152\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__12149\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2954\ : IoInMux
    port map (
            O => \N__12140\,
            I => \N__12137\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__12137\,
            I => \N__12134\
        );

    \I__2952\ : Span4Mux_s1_v
    port map (
            O => \N__12134\,
            I => \N__12131\
        );

    \I__2951\ : Span4Mux_v
    port map (
            O => \N__12131\,
            I => \N__12128\
        );

    \I__2950\ : Span4Mux_v
    port map (
            O => \N__12128\,
            I => \N__12125\
        );

    \I__2949\ : Odrv4
    port map (
            O => \N__12125\,
            I => \CRCSn_c\
        );

    \I__2948\ : InMux
    port map (
            O => \N__12122\,
            I => \N__12116\
        );

    \I__2947\ : InMux
    port map (
            O => \N__12121\,
            I => \N__12113\
        );

    \I__2946\ : InMux
    port map (
            O => \N__12120\,
            I => \N__12110\
        );

    \I__2945\ : InMux
    port map (
            O => \N__12119\,
            I => \N__12107\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__12116\,
            I => \N__12102\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__12113\,
            I => \N__12102\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__12110\,
            I => \N__12099\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__12107\,
            I => \N__12096\
        );

    \I__2940\ : Span4Mux_v
    port map (
            O => \N__12102\,
            I => \N__12093\
        );

    \I__2939\ : Span4Mux_h
    port map (
            O => \N__12099\,
            I => \N__12090\
        );

    \I__2938\ : Span12Mux_v
    port map (
            O => \N__12096\,
            I => \N__12085\
        );

    \I__2937\ : Sp12to4
    port map (
            O => \N__12093\,
            I => \N__12085\
        );

    \I__2936\ : Span4Mux_v
    port map (
            O => \N__12090\,
            I => \N__12082\
        );

    \I__2935\ : Span12Mux_h
    port map (
            O => \N__12085\,
            I => \N__12079\
        );

    \I__2934\ : Span4Mux_h
    port map (
            O => \N__12082\,
            I => \N__12076\
        );

    \I__2933\ : Odrv12
    port map (
            O => \N__12079\,
            I => \DRA_c_7\
        );

    \I__2932\ : Odrv4
    port map (
            O => \N__12076\,
            I => \DRA_c_7\
        );

    \I__2931\ : InMux
    port map (
            O => \N__12071\,
            I => \N__12065\
        );

    \I__2930\ : InMux
    port map (
            O => \N__12070\,
            I => \N__12062\
        );

    \I__2929\ : InMux
    port map (
            O => \N__12069\,
            I => \N__12059\
        );

    \I__2928\ : InMux
    port map (
            O => \N__12068\,
            I => \N__12056\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__12065\,
            I => \N__12051\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__12062\,
            I => \N__12051\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__12059\,
            I => \N__12046\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__12056\,
            I => \N__12046\
        );

    \I__2923\ : Span4Mux_v
    port map (
            O => \N__12051\,
            I => \N__12043\
        );

    \I__2922\ : Span4Mux_v
    port map (
            O => \N__12046\,
            I => \N__12040\
        );

    \I__2921\ : Sp12to4
    port map (
            O => \N__12043\,
            I => \N__12037\
        );

    \I__2920\ : Sp12to4
    port map (
            O => \N__12040\,
            I => \N__12034\
        );

    \I__2919\ : Span12Mux_h
    port map (
            O => \N__12037\,
            I => \N__12031\
        );

    \I__2918\ : Odrv12
    port map (
            O => \N__12034\,
            I => \DRA_c_8\
        );

    \I__2917\ : Odrv12
    port map (
            O => \N__12031\,
            I => \DRA_c_8\
        );

    \I__2916\ : InMux
    port map (
            O => \N__12026\,
            I => \N__12023\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__12023\,
            I => \N__12020\
        );

    \I__2914\ : Span4Mux_h
    port map (
            O => \N__12020\,
            I => \N__12017\
        );

    \I__2913\ : Odrv4
    port map (
            O => \N__12017\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2912\ : InMux
    port map (
            O => \N__12014\,
            I => \N__12010\
        );

    \I__2911\ : InMux
    port map (
            O => \N__12013\,
            I => \N__12007\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__12010\,
            I => \N__12000\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__12007\,
            I => \N__12000\
        );

    \I__2908\ : InMux
    port map (
            O => \N__12006\,
            I => \N__11995\
        );

    \I__2907\ : InMux
    port map (
            O => \N__12005\,
            I => \N__11995\
        );

    \I__2906\ : Span4Mux_v
    port map (
            O => \N__12000\,
            I => \N__11992\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__11995\,
            I => \N__11989\
        );

    \I__2904\ : Sp12to4
    port map (
            O => \N__11992\,
            I => \N__11986\
        );

    \I__2903\ : Span12Mux_v
    port map (
            O => \N__11989\,
            I => \N__11983\
        );

    \I__2902\ : Span12Mux_h
    port map (
            O => \N__11986\,
            I => \N__11980\
        );

    \I__2901\ : Span12Mux_h
    port map (
            O => \N__11983\,
            I => \N__11977\
        );

    \I__2900\ : Span12Mux_v
    port map (
            O => \N__11980\,
            I => \N__11974\
        );

    \I__2899\ : Odrv12
    port map (
            O => \N__11977\,
            I => \DRA_c_2\
        );

    \I__2898\ : Odrv12
    port map (
            O => \N__11974\,
            I => \DRA_c_2\
        );

    \I__2897\ : InMux
    port map (
            O => \N__11969\,
            I => \N__11966\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__11966\,
            I => \N__11961\
        );

    \I__2895\ : InMux
    port map (
            O => \N__11965\,
            I => \N__11958\
        );

    \I__2894\ : InMux
    port map (
            O => \N__11964\,
            I => \N__11955\
        );

    \I__2893\ : Span4Mux_h
    port map (
            O => \N__11961\,
            I => \N__11948\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__11958\,
            I => \N__11948\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__11955\,
            I => \N__11948\
        );

    \I__2890\ : Span4Mux_v
    port map (
            O => \N__11948\,
            I => \N__11944\
        );

    \I__2889\ : InMux
    port map (
            O => \N__11947\,
            I => \N__11941\
        );

    \I__2888\ : Span4Mux_v
    port map (
            O => \N__11944\,
            I => \N__11938\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__11941\,
            I => \N__11935\
        );

    \I__2886\ : Span4Mux_h
    port map (
            O => \N__11938\,
            I => \N__11932\
        );

    \I__2885\ : Sp12to4
    port map (
            O => \N__11935\,
            I => \N__11929\
        );

    \I__2884\ : Sp12to4
    port map (
            O => \N__11932\,
            I => \N__11924\
        );

    \I__2883\ : Span12Mux_v
    port map (
            O => \N__11929\,
            I => \N__11924\
        );

    \I__2882\ : Odrv12
    port map (
            O => \N__11924\,
            I => \DRA_c_3\
        );

    \I__2881\ : InMux
    port map (
            O => \N__11921\,
            I => \N__11918\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__11918\,
            I => \N__11915\
        );

    \I__2879\ : Span4Mux_h
    port map (
            O => \N__11915\,
            I => \N__11912\
        );

    \I__2878\ : Span4Mux_h
    port map (
            O => \N__11912\,
            I => \N__11909\
        );

    \I__2877\ : Odrv4
    port map (
            O => \N__11909\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__2876\ : CascadeMux
    port map (
            O => \N__11906\,
            I => \N__11903\
        );

    \I__2875\ : InMux
    port map (
            O => \N__11903\,
            I => \N__11899\
        );

    \I__2874\ : InMux
    port map (
            O => \N__11902\,
            I => \N__11896\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__11899\,
            I => \N__11892\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__11896\,
            I => \N__11889\
        );

    \I__2871\ : InMux
    port map (
            O => \N__11895\,
            I => \N__11886\
        );

    \I__2870\ : Span4Mux_h
    port map (
            O => \N__11892\,
            I => \N__11880\
        );

    \I__2869\ : Span4Mux_v
    port map (
            O => \N__11889\,
            I => \N__11880\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__11886\,
            I => \N__11877\
        );

    \I__2867\ : InMux
    port map (
            O => \N__11885\,
            I => \N__11874\
        );

    \I__2866\ : Span4Mux_v
    port map (
            O => \N__11880\,
            I => \N__11871\
        );

    \I__2865\ : Span4Mux_h
    port map (
            O => \N__11877\,
            I => \N__11868\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__11874\,
            I => \N__11865\
        );

    \I__2863\ : Sp12to4
    port map (
            O => \N__11871\,
            I => \N__11862\
        );

    \I__2862\ : Span4Mux_v
    port map (
            O => \N__11868\,
            I => \N__11859\
        );

    \I__2861\ : Span4Mux_v
    port map (
            O => \N__11865\,
            I => \N__11856\
        );

    \I__2860\ : Span12Mux_h
    port map (
            O => \N__11862\,
            I => \N__11853\
        );

    \I__2859\ : Sp12to4
    port map (
            O => \N__11859\,
            I => \N__11848\
        );

    \I__2858\ : Sp12to4
    port map (
            O => \N__11856\,
            I => \N__11848\
        );

    \I__2857\ : Span12Mux_v
    port map (
            O => \N__11853\,
            I => \N__11845\
        );

    \I__2856\ : Span12Mux_v
    port map (
            O => \N__11848\,
            I => \N__11842\
        );

    \I__2855\ : Odrv12
    port map (
            O => \N__11845\,
            I => \DRA_c_9\
        );

    \I__2854\ : Odrv12
    port map (
            O => \N__11842\,
            I => \DRA_c_9\
        );

    \I__2853\ : CascadeMux
    port map (
            O => \N__11837\,
            I => \N__11832\
        );

    \I__2852\ : CascadeMux
    port map (
            O => \N__11836\,
            I => \N__11824\
        );

    \I__2851\ : InMux
    port map (
            O => \N__11835\,
            I => \N__11820\
        );

    \I__2850\ : InMux
    port map (
            O => \N__11832\,
            I => \N__11816\
        );

    \I__2849\ : InMux
    port map (
            O => \N__11831\,
            I => \N__11813\
        );

    \I__2848\ : InMux
    port map (
            O => \N__11830\,
            I => \N__11808\
        );

    \I__2847\ : InMux
    port map (
            O => \N__11829\,
            I => \N__11805\
        );

    \I__2846\ : InMux
    port map (
            O => \N__11828\,
            I => \N__11802\
        );

    \I__2845\ : InMux
    port map (
            O => \N__11827\,
            I => \N__11795\
        );

    \I__2844\ : InMux
    port map (
            O => \N__11824\,
            I => \N__11790\
        );

    \I__2843\ : InMux
    port map (
            O => \N__11823\,
            I => \N__11790\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__11820\,
            I => \N__11787\
        );

    \I__2841\ : InMux
    port map (
            O => \N__11819\,
            I => \N__11784\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__11816\,
            I => \N__11781\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__11813\,
            I => \N__11778\
        );

    \I__2838\ : InMux
    port map (
            O => \N__11812\,
            I => \N__11775\
        );

    \I__2837\ : InMux
    port map (
            O => \N__11811\,
            I => \N__11772\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__11808\,
            I => \N__11765\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__11805\,
            I => \N__11765\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__11802\,
            I => \N__11765\
        );

    \I__2833\ : InMux
    port map (
            O => \N__11801\,
            I => \N__11762\
        );

    \I__2832\ : InMux
    port map (
            O => \N__11800\,
            I => \N__11754\
        );

    \I__2831\ : InMux
    port map (
            O => \N__11799\,
            I => \N__11751\
        );

    \I__2830\ : InMux
    port map (
            O => \N__11798\,
            I => \N__11748\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__11795\,
            I => \N__11743\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__11790\,
            I => \N__11743\
        );

    \I__2827\ : Span4Mux_v
    port map (
            O => \N__11787\,
            I => \N__11738\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__11784\,
            I => \N__11738\
        );

    \I__2825\ : Span4Mux_h
    port map (
            O => \N__11781\,
            I => \N__11725\
        );

    \I__2824\ : Span4Mux_v
    port map (
            O => \N__11778\,
            I => \N__11725\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__11775\,
            I => \N__11725\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__11772\,
            I => \N__11725\
        );

    \I__2821\ : Span4Mux_v
    port map (
            O => \N__11765\,
            I => \N__11725\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__11762\,
            I => \N__11725\
        );

    \I__2819\ : InMux
    port map (
            O => \N__11761\,
            I => \N__11720\
        );

    \I__2818\ : InMux
    port map (
            O => \N__11760\,
            I => \N__11720\
        );

    \I__2817\ : InMux
    port map (
            O => \N__11759\,
            I => \N__11717\
        );

    \I__2816\ : InMux
    port map (
            O => \N__11758\,
            I => \N__11712\
        );

    \I__2815\ : InMux
    port map (
            O => \N__11757\,
            I => \N__11712\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__11754\,
            I => \N__11703\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__11751\,
            I => \N__11703\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__11748\,
            I => \N__11703\
        );

    \I__2811\ : Span4Mux_v
    port map (
            O => \N__11743\,
            I => \N__11703\
        );

    \I__2810\ : Span4Mux_v
    port map (
            O => \N__11738\,
            I => \N__11700\
        );

    \I__2809\ : Span4Mux_h
    port map (
            O => \N__11725\,
            I => \N__11697\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__11720\,
            I => \N__11694\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__11717\,
            I => \N__11685\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__11712\,
            I => \N__11685\
        );

    \I__2805\ : Sp12to4
    port map (
            O => \N__11703\,
            I => \N__11685\
        );

    \I__2804\ : Sp12to4
    port map (
            O => \N__11700\,
            I => \N__11685\
        );

    \I__2803\ : Sp12to4
    port map (
            O => \N__11697\,
            I => \N__11682\
        );

    \I__2802\ : Span12Mux_v
    port map (
            O => \N__11694\,
            I => \N__11679\
        );

    \I__2801\ : Span12Mux_h
    port map (
            O => \N__11685\,
            I => \N__11676\
        );

    \I__2800\ : Span12Mux_v
    port map (
            O => \N__11682\,
            I => \N__11673\
        );

    \I__2799\ : Span12Mux_h
    port map (
            O => \N__11679\,
            I => \N__11668\
        );

    \I__2798\ : Span12Mux_v
    port map (
            O => \N__11676\,
            I => \N__11668\
        );

    \I__2797\ : Span12Mux_h
    port map (
            O => \N__11673\,
            I => \N__11665\
        );

    \I__2796\ : Odrv12
    port map (
            O => \N__11668\,
            I => \AGNUS_REV_c\
        );

    \I__2795\ : Odrv12
    port map (
            O => \N__11665\,
            I => \AGNUS_REV_c\
        );

    \I__2794\ : InMux
    port map (
            O => \N__11660\,
            I => \N__11657\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__11657\,
            I => \N__11654\
        );

    \I__2792\ : Span4Mux_h
    port map (
            O => \N__11654\,
            I => \N__11651\
        );

    \I__2791\ : Odrv4
    port map (
            O => \N__11651\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2790\ : ClkMux
    port map (
            O => \N__11648\,
            I => \N__11627\
        );

    \I__2789\ : ClkMux
    port map (
            O => \N__11647\,
            I => \N__11627\
        );

    \I__2788\ : ClkMux
    port map (
            O => \N__11646\,
            I => \N__11627\
        );

    \I__2787\ : ClkMux
    port map (
            O => \N__11645\,
            I => \N__11627\
        );

    \I__2786\ : ClkMux
    port map (
            O => \N__11644\,
            I => \N__11627\
        );

    \I__2785\ : ClkMux
    port map (
            O => \N__11643\,
            I => \N__11627\
        );

    \I__2784\ : ClkMux
    port map (
            O => \N__11642\,
            I => \N__11627\
        );

    \I__2783\ : GlobalMux
    port map (
            O => \N__11627\,
            I => \N__11624\
        );

    \I__2782\ : gio2CtrlBuf
    port map (
            O => \N__11624\,
            I => \C3_c_g\
        );

    \I__2781\ : CEMux
    port map (
            O => \N__11621\,
            I => \N__11582\
        );

    \I__2780\ : CEMux
    port map (
            O => \N__11620\,
            I => \N__11582\
        );

    \I__2779\ : CEMux
    port map (
            O => \N__11619\,
            I => \N__11582\
        );

    \I__2778\ : CEMux
    port map (
            O => \N__11618\,
            I => \N__11582\
        );

    \I__2777\ : CEMux
    port map (
            O => \N__11617\,
            I => \N__11582\
        );

    \I__2776\ : CEMux
    port map (
            O => \N__11616\,
            I => \N__11582\
        );

    \I__2775\ : CEMux
    port map (
            O => \N__11615\,
            I => \N__11582\
        );

    \I__2774\ : CEMux
    port map (
            O => \N__11614\,
            I => \N__11582\
        );

    \I__2773\ : CEMux
    port map (
            O => \N__11613\,
            I => \N__11582\
        );

    \I__2772\ : CEMux
    port map (
            O => \N__11612\,
            I => \N__11582\
        );

    \I__2771\ : CEMux
    port map (
            O => \N__11611\,
            I => \N__11582\
        );

    \I__2770\ : CEMux
    port map (
            O => \N__11610\,
            I => \N__11582\
        );

    \I__2769\ : CEMux
    port map (
            O => \N__11609\,
            I => \N__11582\
        );

    \I__2768\ : GlobalMux
    port map (
            O => \N__11582\,
            I => \N__11579\
        );

    \I__2767\ : gio2CtrlBuf
    port map (
            O => \N__11579\,
            I => \DBRn_c_i_0_g\
        );

    \I__2766\ : InMux
    port map (
            O => \N__11576\,
            I => \N__11566\
        );

    \I__2765\ : InMux
    port map (
            O => \N__11575\,
            I => \N__11563\
        );

    \I__2764\ : InMux
    port map (
            O => \N__11574\,
            I => \N__11558\
        );

    \I__2763\ : InMux
    port map (
            O => \N__11573\,
            I => \N__11558\
        );

    \I__2762\ : InMux
    port map (
            O => \N__11572\,
            I => \N__11555\
        );

    \I__2761\ : InMux
    port map (
            O => \N__11571\,
            I => \N__11552\
        );

    \I__2760\ : InMux
    port map (
            O => \N__11570\,
            I => \N__11549\
        );

    \I__2759\ : InMux
    port map (
            O => \N__11569\,
            I => \N__11546\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__11566\,
            I => \N__11541\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__11563\,
            I => \N__11526\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__11558\,
            I => \N__11523\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__11555\,
            I => \N__11515\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__11552\,
            I => \N__11502\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__11549\,
            I => \N__11496\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__11546\,
            I => \N__11485\
        );

    \I__2751\ : SRMux
    port map (
            O => \N__11545\,
            I => \N__11366\
        );

    \I__2750\ : SRMux
    port map (
            O => \N__11544\,
            I => \N__11366\
        );

    \I__2749\ : Glb2LocalMux
    port map (
            O => \N__11541\,
            I => \N__11366\
        );

    \I__2748\ : SRMux
    port map (
            O => \N__11540\,
            I => \N__11366\
        );

    \I__2747\ : SRMux
    port map (
            O => \N__11539\,
            I => \N__11366\
        );

    \I__2746\ : SRMux
    port map (
            O => \N__11538\,
            I => \N__11366\
        );

    \I__2745\ : SRMux
    port map (
            O => \N__11537\,
            I => \N__11366\
        );

    \I__2744\ : SRMux
    port map (
            O => \N__11536\,
            I => \N__11366\
        );

    \I__2743\ : SRMux
    port map (
            O => \N__11535\,
            I => \N__11366\
        );

    \I__2742\ : SRMux
    port map (
            O => \N__11534\,
            I => \N__11366\
        );

    \I__2741\ : SRMux
    port map (
            O => \N__11533\,
            I => \N__11366\
        );

    \I__2740\ : SRMux
    port map (
            O => \N__11532\,
            I => \N__11366\
        );

    \I__2739\ : SRMux
    port map (
            O => \N__11531\,
            I => \N__11366\
        );

    \I__2738\ : SRMux
    port map (
            O => \N__11530\,
            I => \N__11366\
        );

    \I__2737\ : SRMux
    port map (
            O => \N__11529\,
            I => \N__11366\
        );

    \I__2736\ : Glb2LocalMux
    port map (
            O => \N__11526\,
            I => \N__11366\
        );

    \I__2735\ : Glb2LocalMux
    port map (
            O => \N__11523\,
            I => \N__11366\
        );

    \I__2734\ : SRMux
    port map (
            O => \N__11522\,
            I => \N__11366\
        );

    \I__2733\ : SRMux
    port map (
            O => \N__11521\,
            I => \N__11366\
        );

    \I__2732\ : SRMux
    port map (
            O => \N__11520\,
            I => \N__11366\
        );

    \I__2731\ : SRMux
    port map (
            O => \N__11519\,
            I => \N__11366\
        );

    \I__2730\ : SRMux
    port map (
            O => \N__11518\,
            I => \N__11366\
        );

    \I__2729\ : Glb2LocalMux
    port map (
            O => \N__11515\,
            I => \N__11366\
        );

    \I__2728\ : SRMux
    port map (
            O => \N__11514\,
            I => \N__11366\
        );

    \I__2727\ : SRMux
    port map (
            O => \N__11513\,
            I => \N__11366\
        );

    \I__2726\ : SRMux
    port map (
            O => \N__11512\,
            I => \N__11366\
        );

    \I__2725\ : SRMux
    port map (
            O => \N__11511\,
            I => \N__11366\
        );

    \I__2724\ : SRMux
    port map (
            O => \N__11510\,
            I => \N__11366\
        );

    \I__2723\ : SRMux
    port map (
            O => \N__11509\,
            I => \N__11366\
        );

    \I__2722\ : SRMux
    port map (
            O => \N__11508\,
            I => \N__11366\
        );

    \I__2721\ : SRMux
    port map (
            O => \N__11507\,
            I => \N__11366\
        );

    \I__2720\ : SRMux
    port map (
            O => \N__11506\,
            I => \N__11366\
        );

    \I__2719\ : SRMux
    port map (
            O => \N__11505\,
            I => \N__11366\
        );

    \I__2718\ : Glb2LocalMux
    port map (
            O => \N__11502\,
            I => \N__11366\
        );

    \I__2717\ : SRMux
    port map (
            O => \N__11501\,
            I => \N__11366\
        );

    \I__2716\ : SRMux
    port map (
            O => \N__11500\,
            I => \N__11366\
        );

    \I__2715\ : SRMux
    port map (
            O => \N__11499\,
            I => \N__11366\
        );

    \I__2714\ : Glb2LocalMux
    port map (
            O => \N__11496\,
            I => \N__11366\
        );

    \I__2713\ : SRMux
    port map (
            O => \N__11495\,
            I => \N__11366\
        );

    \I__2712\ : SRMux
    port map (
            O => \N__11494\,
            I => \N__11366\
        );

    \I__2711\ : SRMux
    port map (
            O => \N__11493\,
            I => \N__11366\
        );

    \I__2710\ : SRMux
    port map (
            O => \N__11492\,
            I => \N__11366\
        );

    \I__2709\ : SRMux
    port map (
            O => \N__11491\,
            I => \N__11366\
        );

    \I__2708\ : SRMux
    port map (
            O => \N__11490\,
            I => \N__11366\
        );

    \I__2707\ : SRMux
    port map (
            O => \N__11489\,
            I => \N__11366\
        );

    \I__2706\ : SRMux
    port map (
            O => \N__11488\,
            I => \N__11366\
        );

    \I__2705\ : Glb2LocalMux
    port map (
            O => \N__11485\,
            I => \N__11366\
        );

    \I__2704\ : SRMux
    port map (
            O => \N__11484\,
            I => \N__11366\
        );

    \I__2703\ : SRMux
    port map (
            O => \N__11483\,
            I => \N__11366\
        );

    \I__2702\ : SRMux
    port map (
            O => \N__11482\,
            I => \N__11366\
        );

    \I__2701\ : SRMux
    port map (
            O => \N__11481\,
            I => \N__11366\
        );

    \I__2700\ : SRMux
    port map (
            O => \N__11480\,
            I => \N__11366\
        );

    \I__2699\ : SRMux
    port map (
            O => \N__11479\,
            I => \N__11366\
        );

    \I__2698\ : SRMux
    port map (
            O => \N__11478\,
            I => \N__11366\
        );

    \I__2697\ : SRMux
    port map (
            O => \N__11477\,
            I => \N__11366\
        );

    \I__2696\ : GlobalMux
    port map (
            O => \N__11366\,
            I => \N__11363\
        );

    \I__2695\ : gio2CtrlBuf
    port map (
            O => \N__11363\,
            I => \RESETn_c_i_g\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__11360\,
            I => \N__11353\
        );

    \I__2693\ : InMux
    port map (
            O => \N__11359\,
            I => \N__11345\
        );

    \I__2692\ : InMux
    port map (
            O => \N__11358\,
            I => \N__11342\
        );

    \I__2691\ : InMux
    port map (
            O => \N__11357\,
            I => \N__11339\
        );

    \I__2690\ : CascadeMux
    port map (
            O => \N__11356\,
            I => \N__11335\
        );

    \I__2689\ : InMux
    port map (
            O => \N__11353\,
            I => \N__11325\
        );

    \I__2688\ : InMux
    port map (
            O => \N__11352\,
            I => \N__11325\
        );

    \I__2687\ : InMux
    port map (
            O => \N__11351\,
            I => \N__11325\
        );

    \I__2686\ : InMux
    port map (
            O => \N__11350\,
            I => \N__11318\
        );

    \I__2685\ : InMux
    port map (
            O => \N__11349\,
            I => \N__11318\
        );

    \I__2684\ : InMux
    port map (
            O => \N__11348\,
            I => \N__11318\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__11345\,
            I => \N__11313\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__11342\,
            I => \N__11308\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__11339\,
            I => \N__11308\
        );

    \I__2680\ : InMux
    port map (
            O => \N__11338\,
            I => \N__11305\
        );

    \I__2679\ : InMux
    port map (
            O => \N__11335\,
            I => \N__11302\
        );

    \I__2678\ : InMux
    port map (
            O => \N__11334\,
            I => \N__11295\
        );

    \I__2677\ : InMux
    port map (
            O => \N__11333\,
            I => \N__11295\
        );

    \I__2676\ : InMux
    port map (
            O => \N__11332\,
            I => \N__11292\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__11325\,
            I => \N__11285\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__11318\,
            I => \N__11285\
        );

    \I__2673\ : InMux
    port map (
            O => \N__11317\,
            I => \N__11280\
        );

    \I__2672\ : InMux
    port map (
            O => \N__11316\,
            I => \N__11280\
        );

    \I__2671\ : Span4Mux_v
    port map (
            O => \N__11313\,
            I => \N__11271\
        );

    \I__2670\ : Span4Mux_v
    port map (
            O => \N__11308\,
            I => \N__11271\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__11305\,
            I => \N__11271\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__11302\,
            I => \N__11271\
        );

    \I__2667\ : InMux
    port map (
            O => \N__11301\,
            I => \N__11266\
        );

    \I__2666\ : InMux
    port map (
            O => \N__11300\,
            I => \N__11266\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__11295\,
            I => \N__11258\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__11292\,
            I => \N__11258\
        );

    \I__2663\ : InMux
    port map (
            O => \N__11291\,
            I => \N__11253\
        );

    \I__2662\ : InMux
    port map (
            O => \N__11290\,
            I => \N__11253\
        );

    \I__2661\ : Span4Mux_v
    port map (
            O => \N__11285\,
            I => \N__11239\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__11280\,
            I => \N__11236\
        );

    \I__2659\ : Span4Mux_h
    port map (
            O => \N__11271\,
            I => \N__11231\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__11266\,
            I => \N__11231\
        );

    \I__2657\ : InMux
    port map (
            O => \N__11265\,
            I => \N__11226\
        );

    \I__2656\ : InMux
    port map (
            O => \N__11264\,
            I => \N__11226\
        );

    \I__2655\ : InMux
    port map (
            O => \N__11263\,
            I => \N__11223\
        );

    \I__2654\ : Span4Mux_v
    port map (
            O => \N__11258\,
            I => \N__11218\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__11253\,
            I => \N__11218\
        );

    \I__2652\ : InMux
    port map (
            O => \N__11252\,
            I => \N__11209\
        );

    \I__2651\ : InMux
    port map (
            O => \N__11251\,
            I => \N__11209\
        );

    \I__2650\ : InMux
    port map (
            O => \N__11250\,
            I => \N__11209\
        );

    \I__2649\ : InMux
    port map (
            O => \N__11249\,
            I => \N__11209\
        );

    \I__2648\ : InMux
    port map (
            O => \N__11248\,
            I => \N__11206\
        );

    \I__2647\ : InMux
    port map (
            O => \N__11247\,
            I => \N__11197\
        );

    \I__2646\ : InMux
    port map (
            O => \N__11246\,
            I => \N__11197\
        );

    \I__2645\ : InMux
    port map (
            O => \N__11245\,
            I => \N__11197\
        );

    \I__2644\ : InMux
    port map (
            O => \N__11244\,
            I => \N__11197\
        );

    \I__2643\ : InMux
    port map (
            O => \N__11243\,
            I => \N__11187\
        );

    \I__2642\ : InMux
    port map (
            O => \N__11242\,
            I => \N__11187\
        );

    \I__2641\ : Span4Mux_h
    port map (
            O => \N__11239\,
            I => \N__11178\
        );

    \I__2640\ : Span4Mux_v
    port map (
            O => \N__11236\,
            I => \N__11178\
        );

    \I__2639\ : Span4Mux_v
    port map (
            O => \N__11231\,
            I => \N__11178\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__11226\,
            I => \N__11178\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__11223\,
            I => \N__11175\
        );

    \I__2636\ : Sp12to4
    port map (
            O => \N__11218\,
            I => \N__11170\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__11209\,
            I => \N__11170\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__11206\,
            I => \N__11167\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__11197\,
            I => \N__11164\
        );

    \I__2632\ : InMux
    port map (
            O => \N__11196\,
            I => \N__11155\
        );

    \I__2631\ : InMux
    port map (
            O => \N__11195\,
            I => \N__11155\
        );

    \I__2630\ : InMux
    port map (
            O => \N__11194\,
            I => \N__11155\
        );

    \I__2629\ : InMux
    port map (
            O => \N__11193\,
            I => \N__11155\
        );

    \I__2628\ : InMux
    port map (
            O => \N__11192\,
            I => \N__11152\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__11187\,
            I => \N__11149\
        );

    \I__2626\ : Span4Mux_h
    port map (
            O => \N__11178\,
            I => \N__11144\
        );

    \I__2625\ : Span4Mux_v
    port map (
            O => \N__11175\,
            I => \N__11144\
        );

    \I__2624\ : Span12Mux_v
    port map (
            O => \N__11170\,
            I => \N__11141\
        );

    \I__2623\ : Span12Mux_v
    port map (
            O => \N__11167\,
            I => \N__11132\
        );

    \I__2622\ : Span12Mux_v
    port map (
            O => \N__11164\,
            I => \N__11132\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__11155\,
            I => \N__11132\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__11152\,
            I => \N__11132\
        );

    \I__2619\ : Span12Mux_v
    port map (
            O => \N__11149\,
            I => \N__11129\
        );

    \I__2618\ : Span4Mux_h
    port map (
            O => \N__11144\,
            I => \N__11126\
        );

    \I__2617\ : Span12Mux_h
    port map (
            O => \N__11141\,
            I => \N__11123\
        );

    \I__2616\ : Span12Mux_h
    port map (
            O => \N__11132\,
            I => \N__11120\
        );

    \I__2615\ : Span12Mux_h
    port map (
            O => \N__11129\,
            I => \N__11117\
        );

    \I__2614\ : Span4Mux_h
    port map (
            O => \N__11126\,
            I => \N__11114\
        );

    \I__2613\ : Odrv12
    port map (
            O => \N__11123\,
            I => \RESETn_c\
        );

    \I__2612\ : Odrv12
    port map (
            O => \N__11120\,
            I => \RESETn_c\
        );

    \I__2611\ : Odrv12
    port map (
            O => \N__11117\,
            I => \RESETn_c\
        );

    \I__2610\ : Odrv4
    port map (
            O => \N__11114\,
            I => \RESETn_c\
        );

    \I__2609\ : InMux
    port map (
            O => \N__11105\,
            I => \N__11102\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__11102\,
            I => \N__11099\
        );

    \I__2607\ : Span12Mux_h
    port map (
            O => \N__11099\,
            I => \N__11096\
        );

    \I__2606\ : Odrv12
    port map (
            O => \N__11096\,
            I => \RAS1n_c\
        );

    \I__2605\ : InMux
    port map (
            O => \N__11093\,
            I => \N__11090\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__11090\,
            I => \N__11086\
        );

    \I__2603\ : InMux
    port map (
            O => \N__11089\,
            I => \N__11083\
        );

    \I__2602\ : Sp12to4
    port map (
            O => \N__11086\,
            I => \N__11080\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__11083\,
            I => \N__11077\
        );

    \I__2600\ : Span12Mux_v
    port map (
            O => \N__11080\,
            I => \N__11074\
        );

    \I__2599\ : Span12Mux_h
    port map (
            O => \N__11077\,
            I => \N__11071\
        );

    \I__2598\ : Odrv12
    port map (
            O => \N__11074\,
            I => \RAS0n_c\
        );

    \I__2597\ : Odrv12
    port map (
            O => \N__11071\,
            I => \RAS0n_c\
        );

    \I__2596\ : InMux
    port map (
            O => \N__11066\,
            I => \N__11063\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__11063\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2594\ : InMux
    port map (
            O => \N__11060\,
            I => \N__11057\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__11057\,
            I => \N__11026\
        );

    \I__2592\ : ClkMux
    port map (
            O => \N__11056\,
            I => \N__10892\
        );

    \I__2591\ : ClkMux
    port map (
            O => \N__11055\,
            I => \N__10892\
        );

    \I__2590\ : ClkMux
    port map (
            O => \N__11054\,
            I => \N__10892\
        );

    \I__2589\ : ClkMux
    port map (
            O => \N__11053\,
            I => \N__10892\
        );

    \I__2588\ : ClkMux
    port map (
            O => \N__11052\,
            I => \N__10892\
        );

    \I__2587\ : ClkMux
    port map (
            O => \N__11051\,
            I => \N__10892\
        );

    \I__2586\ : ClkMux
    port map (
            O => \N__11050\,
            I => \N__10892\
        );

    \I__2585\ : ClkMux
    port map (
            O => \N__11049\,
            I => \N__10892\
        );

    \I__2584\ : ClkMux
    port map (
            O => \N__11048\,
            I => \N__10892\
        );

    \I__2583\ : ClkMux
    port map (
            O => \N__11047\,
            I => \N__10892\
        );

    \I__2582\ : ClkMux
    port map (
            O => \N__11046\,
            I => \N__10892\
        );

    \I__2581\ : ClkMux
    port map (
            O => \N__11045\,
            I => \N__10892\
        );

    \I__2580\ : ClkMux
    port map (
            O => \N__11044\,
            I => \N__10892\
        );

    \I__2579\ : ClkMux
    port map (
            O => \N__11043\,
            I => \N__10892\
        );

    \I__2578\ : ClkMux
    port map (
            O => \N__11042\,
            I => \N__10892\
        );

    \I__2577\ : ClkMux
    port map (
            O => \N__11041\,
            I => \N__10892\
        );

    \I__2576\ : ClkMux
    port map (
            O => \N__11040\,
            I => \N__10892\
        );

    \I__2575\ : ClkMux
    port map (
            O => \N__11039\,
            I => \N__10892\
        );

    \I__2574\ : ClkMux
    port map (
            O => \N__11038\,
            I => \N__10892\
        );

    \I__2573\ : ClkMux
    port map (
            O => \N__11037\,
            I => \N__10892\
        );

    \I__2572\ : ClkMux
    port map (
            O => \N__11036\,
            I => \N__10892\
        );

    \I__2571\ : ClkMux
    port map (
            O => \N__11035\,
            I => \N__10892\
        );

    \I__2570\ : ClkMux
    port map (
            O => \N__11034\,
            I => \N__10892\
        );

    \I__2569\ : ClkMux
    port map (
            O => \N__11033\,
            I => \N__10892\
        );

    \I__2568\ : ClkMux
    port map (
            O => \N__11032\,
            I => \N__10892\
        );

    \I__2567\ : ClkMux
    port map (
            O => \N__11031\,
            I => \N__10892\
        );

    \I__2566\ : ClkMux
    port map (
            O => \N__11030\,
            I => \N__10892\
        );

    \I__2565\ : ClkMux
    port map (
            O => \N__11029\,
            I => \N__10892\
        );

    \I__2564\ : Glb2LocalMux
    port map (
            O => \N__11026\,
            I => \N__10892\
        );

    \I__2563\ : ClkMux
    port map (
            O => \N__11025\,
            I => \N__10892\
        );

    \I__2562\ : ClkMux
    port map (
            O => \N__11024\,
            I => \N__10892\
        );

    \I__2561\ : ClkMux
    port map (
            O => \N__11023\,
            I => \N__10892\
        );

    \I__2560\ : ClkMux
    port map (
            O => \N__11022\,
            I => \N__10892\
        );

    \I__2559\ : ClkMux
    port map (
            O => \N__11021\,
            I => \N__10892\
        );

    \I__2558\ : ClkMux
    port map (
            O => \N__11020\,
            I => \N__10892\
        );

    \I__2557\ : ClkMux
    port map (
            O => \N__11019\,
            I => \N__10892\
        );

    \I__2556\ : ClkMux
    port map (
            O => \N__11018\,
            I => \N__10892\
        );

    \I__2555\ : ClkMux
    port map (
            O => \N__11017\,
            I => \N__10892\
        );

    \I__2554\ : ClkMux
    port map (
            O => \N__11016\,
            I => \N__10892\
        );

    \I__2553\ : ClkMux
    port map (
            O => \N__11015\,
            I => \N__10892\
        );

    \I__2552\ : ClkMux
    port map (
            O => \N__11014\,
            I => \N__10892\
        );

    \I__2551\ : ClkMux
    port map (
            O => \N__11013\,
            I => \N__10892\
        );

    \I__2550\ : ClkMux
    port map (
            O => \N__11012\,
            I => \N__10892\
        );

    \I__2549\ : ClkMux
    port map (
            O => \N__11011\,
            I => \N__10892\
        );

    \I__2548\ : ClkMux
    port map (
            O => \N__11010\,
            I => \N__10892\
        );

    \I__2547\ : ClkMux
    port map (
            O => \N__11009\,
            I => \N__10892\
        );

    \I__2546\ : ClkMux
    port map (
            O => \N__11008\,
            I => \N__10892\
        );

    \I__2545\ : ClkMux
    port map (
            O => \N__11007\,
            I => \N__10892\
        );

    \I__2544\ : ClkMux
    port map (
            O => \N__11006\,
            I => \N__10892\
        );

    \I__2543\ : ClkMux
    port map (
            O => \N__11005\,
            I => \N__10892\
        );

    \I__2542\ : ClkMux
    port map (
            O => \N__11004\,
            I => \N__10892\
        );

    \I__2541\ : ClkMux
    port map (
            O => \N__11003\,
            I => \N__10892\
        );

    \I__2540\ : ClkMux
    port map (
            O => \N__11002\,
            I => \N__10892\
        );

    \I__2539\ : ClkMux
    port map (
            O => \N__11001\,
            I => \N__10892\
        );

    \I__2538\ : GlobalMux
    port map (
            O => \N__10892\,
            I => \CLK80_PLL\
        );

    \I__2537\ : InMux
    port map (
            O => \N__10889\,
            I => \N__10884\
        );

    \I__2536\ : CascadeMux
    port map (
            O => \N__10888\,
            I => \N__10881\
        );

    \I__2535\ : InMux
    port map (
            O => \N__10887\,
            I => \N__10877\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__10884\,
            I => \N__10874\
        );

    \I__2533\ : InMux
    port map (
            O => \N__10881\,
            I => \N__10871\
        );

    \I__2532\ : InMux
    port map (
            O => \N__10880\,
            I => \N__10867\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__10877\,
            I => \N__10864\
        );

    \I__2530\ : Span4Mux_h
    port map (
            O => \N__10874\,
            I => \N__10859\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__10871\,
            I => \N__10859\
        );

    \I__2528\ : InMux
    port map (
            O => \N__10870\,
            I => \N__10856\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__10867\,
            I => \N__10853\
        );

    \I__2526\ : Span4Mux_v
    port map (
            O => \N__10864\,
            I => \N__10850\
        );

    \I__2525\ : Span4Mux_v
    port map (
            O => \N__10859\,
            I => \N__10845\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__10856\,
            I => \N__10845\
        );

    \I__2523\ : Span4Mux_v
    port map (
            O => \N__10853\,
            I => \N__10842\
        );

    \I__2522\ : Span4Mux_v
    port map (
            O => \N__10850\,
            I => \N__10839\
        );

    \I__2521\ : Span4Mux_h
    port map (
            O => \N__10845\,
            I => \N__10836\
        );

    \I__2520\ : Sp12to4
    port map (
            O => \N__10842\,
            I => \N__10833\
        );

    \I__2519\ : Sp12to4
    port map (
            O => \N__10839\,
            I => \N__10830\
        );

    \I__2518\ : Sp12to4
    port map (
            O => \N__10836\,
            I => \N__10827\
        );

    \I__2517\ : Span12Mux_h
    port map (
            O => \N__10833\,
            I => \N__10824\
        );

    \I__2516\ : Span12Mux_h
    port map (
            O => \N__10830\,
            I => \N__10819\
        );

    \I__2515\ : Span12Mux_v
    port map (
            O => \N__10827\,
            I => \N__10819\
        );

    \I__2514\ : Span12Mux_v
    port map (
            O => \N__10824\,
            I => \N__10816\
        );

    \I__2513\ : Span12Mux_h
    port map (
            O => \N__10819\,
            I => \N__10813\
        );

    \I__2512\ : Odrv12
    port map (
            O => \N__10816\,
            I => \RnW_c\
        );

    \I__2511\ : Odrv12
    port map (
            O => \N__10813\,
            I => \RnW_c\
        );

    \I__2510\ : InMux
    port map (
            O => \N__10808\,
            I => \N__10804\
        );

    \I__2509\ : InMux
    port map (
            O => \N__10807\,
            I => \N__10801\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__10804\,
            I => \N__10798\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__10801\,
            I => \N__10795\
        );

    \I__2506\ : Span12Mux_s8_h
    port map (
            O => \N__10798\,
            I => \N__10792\
        );

    \I__2505\ : Span12Mux_h
    port map (
            O => \N__10795\,
            I => \N__10789\
        );

    \I__2504\ : Span12Mux_v
    port map (
            O => \N__10792\,
            I => \N__10783\
        );

    \I__2503\ : Span12Mux_v
    port map (
            O => \N__10789\,
            I => \N__10783\
        );

    \I__2502\ : InMux
    port map (
            O => \N__10788\,
            I => \N__10780\
        );

    \I__2501\ : Odrv12
    port map (
            O => \N__10783\,
            I => \DMA_WRITE_CYCLE\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__10780\,
            I => \DMA_WRITE_CYCLE\
        );

    \I__2499\ : CascadeMux
    port map (
            O => \N__10775\,
            I => \N__10772\
        );

    \I__2498\ : InMux
    port map (
            O => \N__10772\,
            I => \N__10768\
        );

    \I__2497\ : CascadeMux
    port map (
            O => \N__10771\,
            I => \N__10765\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__10768\,
            I => \N__10759\
        );

    \I__2495\ : InMux
    port map (
            O => \N__10765\,
            I => \N__10756\
        );

    \I__2494\ : InMux
    port map (
            O => \N__10764\,
            I => \N__10753\
        );

    \I__2493\ : CascadeMux
    port map (
            O => \N__10763\,
            I => \N__10750\
        );

    \I__2492\ : InMux
    port map (
            O => \N__10762\,
            I => \N__10747\
        );

    \I__2491\ : Span4Mux_v
    port map (
            O => \N__10759\,
            I => \N__10740\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__10756\,
            I => \N__10740\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__10753\,
            I => \N__10740\
        );

    \I__2488\ : InMux
    port map (
            O => \N__10750\,
            I => \N__10737\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__10747\,
            I => \N__10734\
        );

    \I__2486\ : Span4Mux_v
    port map (
            O => \N__10740\,
            I => \N__10731\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__10737\,
            I => \N__10728\
        );

    \I__2484\ : Span4Mux_v
    port map (
            O => \N__10734\,
            I => \N__10724\
        );

    \I__2483\ : Span4Mux_h
    port map (
            O => \N__10731\,
            I => \N__10719\
        );

    \I__2482\ : Span4Mux_v
    port map (
            O => \N__10728\,
            I => \N__10719\
        );

    \I__2481\ : CascadeMux
    port map (
            O => \N__10727\,
            I => \N__10716\
        );

    \I__2480\ : Span4Mux_v
    port map (
            O => \N__10724\,
            I => \N__10713\
        );

    \I__2479\ : Sp12to4
    port map (
            O => \N__10719\,
            I => \N__10710\
        );

    \I__2478\ : InMux
    port map (
            O => \N__10716\,
            I => \N__10707\
        );

    \I__2477\ : Sp12to4
    port map (
            O => \N__10713\,
            I => \N__10704\
        );

    \I__2476\ : Span12Mux_h
    port map (
            O => \N__10710\,
            I => \N__10699\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__10707\,
            I => \N__10699\
        );

    \I__2474\ : Span12Mux_h
    port map (
            O => \N__10704\,
            I => \N__10694\
        );

    \I__2473\ : Span12Mux_v
    port map (
            O => \N__10699\,
            I => \N__10694\
        );

    \I__2472\ : Odrv12
    port map (
            O => \N__10694\,
            I => \CASLn_c\
        );

    \I__2471\ : InMux
    port map (
            O => \N__10691\,
            I => \N__10686\
        );

    \I__2470\ : InMux
    port map (
            O => \N__10690\,
            I => \N__10683\
        );

    \I__2469\ : InMux
    port map (
            O => \N__10689\,
            I => \N__10680\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__10686\,
            I => \N__10674\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__10683\,
            I => \N__10674\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__10680\,
            I => \N__10671\
        );

    \I__2465\ : InMux
    port map (
            O => \N__10679\,
            I => \N__10668\
        );

    \I__2464\ : Span4Mux_v
    port map (
            O => \N__10674\,
            I => \N__10663\
        );

    \I__2463\ : Span4Mux_v
    port map (
            O => \N__10671\,
            I => \N__10658\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__10668\,
            I => \N__10658\
        );

    \I__2461\ : InMux
    port map (
            O => \N__10667\,
            I => \N__10655\
        );

    \I__2460\ : InMux
    port map (
            O => \N__10666\,
            I => \N__10652\
        );

    \I__2459\ : Sp12to4
    port map (
            O => \N__10663\,
            I => \N__10649\
        );

    \I__2458\ : Sp12to4
    port map (
            O => \N__10658\,
            I => \N__10644\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__10655\,
            I => \N__10644\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__10652\,
            I => \N__10641\
        );

    \I__2455\ : Span12Mux_h
    port map (
            O => \N__10649\,
            I => \N__10638\
        );

    \I__2454\ : Span12Mux_v
    port map (
            O => \N__10644\,
            I => \N__10635\
        );

    \I__2453\ : Span4Mux_h
    port map (
            O => \N__10641\,
            I => \N__10632\
        );

    \I__2452\ : Span12Mux_v
    port map (
            O => \N__10638\,
            I => \N__10629\
        );

    \I__2451\ : Span12Mux_h
    port map (
            O => \N__10635\,
            I => \N__10626\
        );

    \I__2450\ : Span4Mux_v
    port map (
            O => \N__10632\,
            I => \N__10623\
        );

    \I__2449\ : Odrv12
    port map (
            O => \N__10629\,
            I => \CASUn_c\
        );

    \I__2448\ : Odrv12
    port map (
            O => \N__10626\,
            I => \CASUn_c\
        );

    \I__2447\ : Odrv4
    port map (
            O => \N__10623\,
            I => \CASUn_c\
        );

    \I__2446\ : CascadeMux
    port map (
            O => \N__10616\,
            I => \N__10613\
        );

    \I__2445\ : InMux
    port map (
            O => \N__10613\,
            I => \N__10606\
        );

    \I__2444\ : CascadeMux
    port map (
            O => \N__10612\,
            I => \N__10602\
        );

    \I__2443\ : InMux
    port map (
            O => \N__10611\,
            I => \N__10594\
        );

    \I__2442\ : InMux
    port map (
            O => \N__10610\,
            I => \N__10591\
        );

    \I__2441\ : InMux
    port map (
            O => \N__10609\,
            I => \N__10588\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__10606\,
            I => \N__10583\
        );

    \I__2439\ : InMux
    port map (
            O => \N__10605\,
            I => \N__10576\
        );

    \I__2438\ : InMux
    port map (
            O => \N__10602\,
            I => \N__10576\
        );

    \I__2437\ : InMux
    port map (
            O => \N__10601\,
            I => \N__10576\
        );

    \I__2436\ : InMux
    port map (
            O => \N__10600\,
            I => \N__10569\
        );

    \I__2435\ : InMux
    port map (
            O => \N__10599\,
            I => \N__10569\
        );

    \I__2434\ : InMux
    port map (
            O => \N__10598\,
            I => \N__10569\
        );

    \I__2433\ : CascadeMux
    port map (
            O => \N__10597\,
            I => \N__10566\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__10594\,
            I => \N__10563\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__10591\,
            I => \N__10555\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__10588\,
            I => \N__10555\
        );

    \I__2429\ : InMux
    port map (
            O => \N__10587\,
            I => \N__10543\
        );

    \I__2428\ : InMux
    port map (
            O => \N__10586\,
            I => \N__10543\
        );

    \I__2427\ : Span4Mux_v
    port map (
            O => \N__10583\,
            I => \N__10534\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__10576\,
            I => \N__10534\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__10569\,
            I => \N__10534\
        );

    \I__2424\ : InMux
    port map (
            O => \N__10566\,
            I => \N__10531\
        );

    \I__2423\ : Span4Mux_v
    port map (
            O => \N__10563\,
            I => \N__10528\
        );

    \I__2422\ : InMux
    port map (
            O => \N__10562\,
            I => \N__10525\
        );

    \I__2421\ : InMux
    port map (
            O => \N__10561\,
            I => \N__10520\
        );

    \I__2420\ : InMux
    port map (
            O => \N__10560\,
            I => \N__10520\
        );

    \I__2419\ : Span4Mux_v
    port map (
            O => \N__10555\,
            I => \N__10517\
        );

    \I__2418\ : InMux
    port map (
            O => \N__10554\,
            I => \N__10514\
        );

    \I__2417\ : InMux
    port map (
            O => \N__10553\,
            I => \N__10503\
        );

    \I__2416\ : InMux
    port map (
            O => \N__10552\,
            I => \N__10503\
        );

    \I__2415\ : InMux
    port map (
            O => \N__10551\,
            I => \N__10503\
        );

    \I__2414\ : InMux
    port map (
            O => \N__10550\,
            I => \N__10503\
        );

    \I__2413\ : InMux
    port map (
            O => \N__10549\,
            I => \N__10503\
        );

    \I__2412\ : InMux
    port map (
            O => \N__10548\,
            I => \N__10499\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__10543\,
            I => \N__10496\
        );

    \I__2410\ : InMux
    port map (
            O => \N__10542\,
            I => \N__10493\
        );

    \I__2409\ : InMux
    port map (
            O => \N__10541\,
            I => \N__10490\
        );

    \I__2408\ : Span4Mux_h
    port map (
            O => \N__10534\,
            I => \N__10487\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__10531\,
            I => \N__10472\
        );

    \I__2406\ : Sp12to4
    port map (
            O => \N__10528\,
            I => \N__10472\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__10525\,
            I => \N__10472\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__10520\,
            I => \N__10472\
        );

    \I__2403\ : Sp12to4
    port map (
            O => \N__10517\,
            I => \N__10472\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__10514\,
            I => \N__10472\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__10503\,
            I => \N__10472\
        );

    \I__2400\ : InMux
    port map (
            O => \N__10502\,
            I => \N__10469\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__10499\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2398\ : Odrv4
    port map (
            O => \N__10496\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__10493\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__10490\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2395\ : Odrv4
    port map (
            O => \N__10487\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2394\ : Odrv12
    port map (
            O => \N__10472\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__10469\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2392\ : IoInMux
    port map (
            O => \N__10454\,
            I => \N__10451\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__10451\,
            I => \N__10448\
        );

    \I__2390\ : Span4Mux_s3_v
    port map (
            O => \N__10448\,
            I => \N__10445\
        );

    \I__2389\ : Span4Mux_v
    port map (
            O => \N__10445\,
            I => \N__10442\
        );

    \I__2388\ : Sp12to4
    port map (
            O => \N__10442\,
            I => \N__10439\
        );

    \I__2387\ : Span12Mux_h
    port map (
            O => \N__10439\,
            I => \N__10436\
        );

    \I__2386\ : Odrv12
    port map (
            O => \N__10436\,
            I => \CASn_c\
        );

    \I__2385\ : InMux
    port map (
            O => \N__10433\,
            I => \N__10430\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__10430\,
            I => \N__10426\
        );

    \I__2383\ : InMux
    port map (
            O => \N__10429\,
            I => \N__10423\
        );

    \I__2382\ : Span4Mux_v
    port map (
            O => \N__10426\,
            I => \N__10416\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__10423\,
            I => \N__10416\
        );

    \I__2380\ : CascadeMux
    port map (
            O => \N__10422\,
            I => \N__10412\
        );

    \I__2379\ : InMux
    port map (
            O => \N__10421\,
            I => \N__10408\
        );

    \I__2378\ : Span4Mux_h
    port map (
            O => \N__10416\,
            I => \N__10405\
        );

    \I__2377\ : InMux
    port map (
            O => \N__10415\,
            I => \N__10400\
        );

    \I__2376\ : InMux
    port map (
            O => \N__10412\,
            I => \N__10400\
        );

    \I__2375\ : InMux
    port map (
            O => \N__10411\,
            I => \N__10397\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__10408\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2373\ : Odrv4
    port map (
            O => \N__10405\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__10400\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__10397\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2370\ : IoInMux
    port map (
            O => \N__10388\,
            I => \N__10385\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__10385\,
            I => \N__10382\
        );

    \I__2368\ : Span4Mux_s3_v
    port map (
            O => \N__10382\,
            I => \N__10379\
        );

    \I__2367\ : Span4Mux_v
    port map (
            O => \N__10379\,
            I => \N__10376\
        );

    \I__2366\ : Span4Mux_h
    port map (
            O => \N__10376\,
            I => \N__10373\
        );

    \I__2365\ : Odrv4
    port map (
            O => \N__10373\,
            I => \RASn_c\
        );

    \I__2364\ : CascadeMux
    port map (
            O => \N__10370\,
            I => \N__10367\
        );

    \I__2363\ : InMux
    port map (
            O => \N__10367\,
            I => \N__10364\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__10364\,
            I => \N__10361\
        );

    \I__2361\ : Span4Mux_h
    port map (
            O => \N__10361\,
            I => \N__10358\
        );

    \I__2360\ : Odrv4
    port map (
            O => \N__10358\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__2359\ : InMux
    port map (
            O => \N__10355\,
            I => \N__10349\
        );

    \I__2358\ : InMux
    port map (
            O => \N__10354\,
            I => \N__10344\
        );

    \I__2357\ : InMux
    port map (
            O => \N__10353\,
            I => \N__10344\
        );

    \I__2356\ : InMux
    port map (
            O => \N__10352\,
            I => \N__10341\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__10349\,
            I => \N__10338\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__10344\,
            I => \N__10333\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__10341\,
            I => \N__10333\
        );

    \I__2352\ : Span4Mux_v
    port map (
            O => \N__10338\,
            I => \N__10330\
        );

    \I__2351\ : Span12Mux_v
    port map (
            O => \N__10333\,
            I => \N__10327\
        );

    \I__2350\ : Span4Mux_v
    port map (
            O => \N__10330\,
            I => \N__10324\
        );

    \I__2349\ : Span12Mux_h
    port map (
            O => \N__10327\,
            I => \N__10321\
        );

    \I__2348\ : Sp12to4
    port map (
            O => \N__10324\,
            I => \N__10318\
        );

    \I__2347\ : Odrv12
    port map (
            O => \N__10321\,
            I => \DRA_c_5\
        );

    \I__2346\ : Odrv12
    port map (
            O => \N__10318\,
            I => \DRA_c_5\
        );

    \I__2345\ : InMux
    port map (
            O => \N__10313\,
            I => \N__10309\
        );

    \I__2344\ : InMux
    port map (
            O => \N__10312\,
            I => \N__10306\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__10309\,
            I => \N__10299\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__10306\,
            I => \N__10299\
        );

    \I__2341\ : InMux
    port map (
            O => \N__10305\,
            I => \N__10296\
        );

    \I__2340\ : InMux
    port map (
            O => \N__10304\,
            I => \N__10293\
        );

    \I__2339\ : Span4Mux_h
    port map (
            O => \N__10299\,
            I => \N__10288\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__10296\,
            I => \N__10288\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__10293\,
            I => \N__10283\
        );

    \I__2336\ : Sp12to4
    port map (
            O => \N__10288\,
            I => \N__10283\
        );

    \I__2335\ : Span12Mux_v
    port map (
            O => \N__10283\,
            I => \N__10280\
        );

    \I__2334\ : Span12Mux_h
    port map (
            O => \N__10280\,
            I => \N__10277\
        );

    \I__2333\ : Odrv12
    port map (
            O => \N__10277\,
            I => \DRA_c_4\
        );

    \I__2332\ : InMux
    port map (
            O => \N__10274\,
            I => \N__10271\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__10271\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__2330\ : InMux
    port map (
            O => \N__10268\,
            I => \N__10264\
        );

    \I__2329\ : InMux
    port map (
            O => \N__10267\,
            I => \N__10261\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__10264\,
            I => \N__10256\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__10261\,
            I => \N__10256\
        );

    \I__2326\ : Span4Mux_h
    port map (
            O => \N__10256\,
            I => \N__10253\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__10253\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__2324\ : InMux
    port map (
            O => \N__10250\,
            I => \N__10246\
        );

    \I__2323\ : InMux
    port map (
            O => \N__10249\,
            I => \N__10243\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__10246\,
            I => \N__10240\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__10243\,
            I => \N__10235\
        );

    \I__2320\ : Span4Mux_v
    port map (
            O => \N__10240\,
            I => \N__10232\
        );

    \I__2319\ : InMux
    port map (
            O => \N__10239\,
            I => \N__10229\
        );

    \I__2318\ : InMux
    port map (
            O => \N__10238\,
            I => \N__10226\
        );

    \I__2317\ : Sp12to4
    port map (
            O => \N__10235\,
            I => \N__10223\
        );

    \I__2316\ : Sp12to4
    port map (
            O => \N__10232\,
            I => \N__10216\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__10229\,
            I => \N__10216\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__10226\,
            I => \N__10216\
        );

    \I__2313\ : Span12Mux_v
    port map (
            O => \N__10223\,
            I => \N__10213\
        );

    \I__2312\ : Span12Mux_h
    port map (
            O => \N__10216\,
            I => \N__10210\
        );

    \I__2311\ : Span12Mux_h
    port map (
            O => \N__10213\,
            I => \N__10205\
        );

    \I__2310\ : Span12Mux_v
    port map (
            O => \N__10210\,
            I => \N__10205\
        );

    \I__2309\ : Odrv12
    port map (
            O => \N__10205\,
            I => \DRA_c_1\
        );

    \I__2308\ : InMux
    port map (
            O => \N__10202\,
            I => \N__10198\
        );

    \I__2307\ : InMux
    port map (
            O => \N__10201\,
            I => \N__10195\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__10198\,
            I => \N__10190\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__10195\,
            I => \N__10190\
        );

    \I__2304\ : Sp12to4
    port map (
            O => \N__10190\,
            I => \N__10187\
        );

    \I__2303\ : Span12Mux_v
    port map (
            O => \N__10187\,
            I => \N__10184\
        );

    \I__2302\ : Span12Mux_h
    port map (
            O => \N__10184\,
            I => \N__10181\
        );

    \I__2301\ : Odrv12
    port map (
            O => \N__10181\,
            I => \DRA_c_0\
        );

    \I__2300\ : InMux
    port map (
            O => \N__10178\,
            I => \N__10175\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__10175\,
            I => \N__10172\
        );

    \I__2298\ : Span4Mux_h
    port map (
            O => \N__10172\,
            I => \N__10169\
        );

    \I__2297\ : Odrv4
    port map (
            O => \N__10169\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__2296\ : InMux
    port map (
            O => \N__10166\,
            I => \N__10163\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__10163\,
            I => \N__10160\
        );

    \I__2294\ : Odrv12
    port map (
            O => \N__10160\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_2\
        );

    \I__2293\ : InMux
    port map (
            O => \N__10157\,
            I => \N__10154\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__10154\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\
        );

    \I__2291\ : InMux
    port map (
            O => \N__10151\,
            I => \N__10148\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__10148\,
            I => \N__10145\
        );

    \I__2289\ : Span4Mux_h
    port map (
            O => \N__10145\,
            I => \N__10142\
        );

    \I__2288\ : Odrv4
    port map (
            O => \N__10142\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__2287\ : InMux
    port map (
            O => \N__10139\,
            I => \N__10136\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__10136\,
            I => \N__10133\
        );

    \I__2285\ : Span4Mux_h
    port map (
            O => \N__10133\,
            I => \N__10130\
        );

    \I__2284\ : Odrv4
    port map (
            O => \N__10130\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__2283\ : InMux
    port map (
            O => \N__10127\,
            I => \N__10124\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__10124\,
            I => \N__10121\
        );

    \I__2281\ : Span4Mux_h
    port map (
            O => \N__10121\,
            I => \N__10118\
        );

    \I__2280\ : Odrv4
    port map (
            O => \N__10118\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__2279\ : CascadeMux
    port map (
            O => \N__10115\,
            I => \N__10112\
        );

    \I__2278\ : InMux
    port map (
            O => \N__10112\,
            I => \N__10109\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__10109\,
            I => \N__10106\
        );

    \I__2276\ : Span4Mux_v
    port map (
            O => \N__10106\,
            I => \N__10103\
        );

    \I__2275\ : Odrv4
    port map (
            O => \N__10103\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2274\ : InMux
    port map (
            O => \N__10100\,
            I => \N__10095\
        );

    \I__2273\ : InMux
    port map (
            O => \N__10099\,
            I => \N__10092\
        );

    \I__2272\ : InMux
    port map (
            O => \N__10098\,
            I => \N__10089\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__10095\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__10092\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__10089\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__2268\ : CascadeMux
    port map (
            O => \N__10082\,
            I => \N__10075\
        );

    \I__2267\ : CascadeMux
    port map (
            O => \N__10081\,
            I => \N__10072\
        );

    \I__2266\ : InMux
    port map (
            O => \N__10080\,
            I => \N__10069\
        );

    \I__2265\ : InMux
    port map (
            O => \N__10079\,
            I => \N__10066\
        );

    \I__2264\ : InMux
    port map (
            O => \N__10078\,
            I => \N__10063\
        );

    \I__2263\ : InMux
    port map (
            O => \N__10075\,
            I => \N__10060\
        );

    \I__2262\ : InMux
    port map (
            O => \N__10072\,
            I => \N__10057\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__10069\,
            I => \N__10054\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__10066\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__10063\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__10060\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__10057\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__2256\ : Odrv4
    port map (
            O => \N__10054\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__2255\ : CascadeMux
    port map (
            O => \N__10043\,
            I => \N__10034\
        );

    \I__2254\ : InMux
    port map (
            O => \N__10042\,
            I => \N__10023\
        );

    \I__2253\ : InMux
    port map (
            O => \N__10041\,
            I => \N__10023\
        );

    \I__2252\ : InMux
    port map (
            O => \N__10040\,
            I => \N__10023\
        );

    \I__2251\ : InMux
    port map (
            O => \N__10039\,
            I => \N__10016\
        );

    \I__2250\ : InMux
    port map (
            O => \N__10038\,
            I => \N__10016\
        );

    \I__2249\ : InMux
    port map (
            O => \N__10037\,
            I => \N__10016\
        );

    \I__2248\ : InMux
    port map (
            O => \N__10034\,
            I => \N__10013\
        );

    \I__2247\ : InMux
    port map (
            O => \N__10033\,
            I => \N__10006\
        );

    \I__2246\ : InMux
    port map (
            O => \N__10032\,
            I => \N__10006\
        );

    \I__2245\ : InMux
    port map (
            O => \N__10031\,
            I => \N__10006\
        );

    \I__2244\ : InMux
    port map (
            O => \N__10030\,
            I => \N__10003\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__10023\,
            I => \N__10000\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__10016\,
            I => \N__9997\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__10013\,
            I => \N__9994\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__10006\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__10003\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__2238\ : Odrv4
    port map (
            O => \N__10000\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__2237\ : Odrv4
    port map (
            O => \N__9997\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__2236\ : Odrv4
    port map (
            O => \N__9994\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__2235\ : InMux
    port map (
            O => \N__9983\,
            I => \N__9980\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__9980\,
            I => \N__9974\
        );

    \I__2233\ : CascadeMux
    port map (
            O => \N__9979\,
            I => \N__9971\
        );

    \I__2232\ : InMux
    port map (
            O => \N__9978\,
            I => \N__9968\
        );

    \I__2231\ : CascadeMux
    port map (
            O => \N__9977\,
            I => \N__9964\
        );

    \I__2230\ : Span4Mux_v
    port map (
            O => \N__9974\,
            I => \N__9959\
        );

    \I__2229\ : InMux
    port map (
            O => \N__9971\,
            I => \N__9956\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__9968\,
            I => \N__9953\
        );

    \I__2227\ : InMux
    port map (
            O => \N__9967\,
            I => \N__9950\
        );

    \I__2226\ : InMux
    port map (
            O => \N__9964\,
            I => \N__9947\
        );

    \I__2225\ : InMux
    port map (
            O => \N__9963\,
            I => \N__9942\
        );

    \I__2224\ : InMux
    port map (
            O => \N__9962\,
            I => \N__9942\
        );

    \I__2223\ : Span4Mux_h
    port map (
            O => \N__9959\,
            I => \N__9937\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__9956\,
            I => \N__9937\
        );

    \I__2221\ : Span4Mux_h
    port map (
            O => \N__9953\,
            I => \N__9934\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__9950\,
            I => \N__9931\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__9947\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_8\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__9942\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_8\
        );

    \I__2217\ : Odrv4
    port map (
            O => \N__9937\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_8\
        );

    \I__2216\ : Odrv4
    port map (
            O => \N__9934\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_8\
        );

    \I__2215\ : Odrv4
    port map (
            O => \N__9931\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_8\
        );

    \I__2214\ : InMux
    port map (
            O => \N__9920\,
            I => \N__9917\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__9917\,
            I => \U712_REG_SM.N_400\
        );

    \I__2212\ : IoInMux
    port map (
            O => \N__9914\,
            I => \N__9911\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__9911\,
            I => \N__9908\
        );

    \I__2210\ : Span4Mux_s2_v
    port map (
            O => \N__9908\,
            I => \N__9905\
        );

    \I__2209\ : Span4Mux_h
    port map (
            O => \N__9905\,
            I => \N__9902\
        );

    \I__2208\ : Span4Mux_h
    port map (
            O => \N__9902\,
            I => \N__9898\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__9901\,
            I => \N__9895\
        );

    \I__2206\ : Sp12to4
    port map (
            O => \N__9898\,
            I => \N__9892\
        );

    \I__2205\ : InMux
    port map (
            O => \N__9895\,
            I => \N__9889\
        );

    \I__2204\ : Odrv12
    port map (
            O => \N__9892\,
            I => \UDSn_c\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__9889\,
            I => \UDSn_c\
        );

    \I__2202\ : InMux
    port map (
            O => \N__9884\,
            I => \N__9879\
        );

    \I__2201\ : InMux
    port map (
            O => \N__9883\,
            I => \N__9873\
        );

    \I__2200\ : InMux
    port map (
            O => \N__9882\,
            I => \N__9873\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__9879\,
            I => \N__9870\
        );

    \I__2198\ : InMux
    port map (
            O => \N__9878\,
            I => \N__9867\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__9873\,
            I => \N__9864\
        );

    \I__2196\ : Odrv4
    port map (
            O => \N__9870\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__9867\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__2194\ : Odrv4
    port map (
            O => \N__9864\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__2193\ : IoInMux
    port map (
            O => \N__9857\,
            I => \N__9854\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__9854\,
            I => \N__9851\
        );

    \I__2191\ : IoSpan4Mux
    port map (
            O => \N__9851\,
            I => \N__9848\
        );

    \I__2190\ : Sp12to4
    port map (
            O => \N__9848\,
            I => \N__9845\
        );

    \I__2189\ : Span12Mux_v
    port map (
            O => \N__9845\,
            I => \N__9841\
        );

    \I__2188\ : InMux
    port map (
            O => \N__9844\,
            I => \N__9838\
        );

    \I__2187\ : Odrv12
    port map (
            O => \N__9841\,
            I => \PRnW_c\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__9838\,
            I => \PRnW_c\
        );

    \I__2185\ : InMux
    port map (
            O => \N__9833\,
            I => \N__9830\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__9830\,
            I => \U712_REG_SM.N_398\
        );

    \I__2183\ : IoInMux
    port map (
            O => \N__9827\,
            I => \N__9824\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__9824\,
            I => \N__9821\
        );

    \I__2181\ : Span4Mux_s3_v
    port map (
            O => \N__9821\,
            I => \N__9818\
        );

    \I__2180\ : Sp12to4
    port map (
            O => \N__9818\,
            I => \N__9814\
        );

    \I__2179\ : CascadeMux
    port map (
            O => \N__9817\,
            I => \N__9811\
        );

    \I__2178\ : Span12Mux_h
    port map (
            O => \N__9814\,
            I => \N__9808\
        );

    \I__2177\ : InMux
    port map (
            O => \N__9811\,
            I => \N__9805\
        );

    \I__2176\ : Odrv12
    port map (
            O => \N__9808\,
            I => \LDSn_c\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__9805\,
            I => \LDSn_c\
        );

    \I__2174\ : IoInMux
    port map (
            O => \N__9800\,
            I => \N__9797\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__9797\,
            I => \N__9794\
        );

    \I__2172\ : IoSpan4Mux
    port map (
            O => \N__9794\,
            I => \N__9791\
        );

    \I__2171\ : Span4Mux_s2_v
    port map (
            O => \N__9791\,
            I => \N__9788\
        );

    \I__2170\ : Span4Mux_v
    port map (
            O => \N__9788\,
            I => \N__9785\
        );

    \I__2169\ : Odrv4
    port map (
            O => \N__9785\,
            I => \N_325_i\
        );

    \I__2168\ : IoInMux
    port map (
            O => \N__9782\,
            I => \N__9779\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__9779\,
            I => \N__9776\
        );

    \I__2166\ : Span4Mux_s2_v
    port map (
            O => \N__9776\,
            I => \N__9773\
        );

    \I__2165\ : Span4Mux_v
    port map (
            O => \N__9773\,
            I => \N__9770\
        );

    \I__2164\ : Odrv4
    port map (
            O => \N__9770\,
            I => \N_323_i\
        );

    \I__2163\ : InMux
    port map (
            O => \N__9767\,
            I => \N__9762\
        );

    \I__2162\ : InMux
    port map (
            O => \N__9766\,
            I => \N__9757\
        );

    \I__2161\ : InMux
    port map (
            O => \N__9765\,
            I => \N__9757\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__9762\,
            I => \N__9747\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__9757\,
            I => \N__9747\
        );

    \I__2158\ : InMux
    port map (
            O => \N__9756\,
            I => \N__9744\
        );

    \I__2157\ : InMux
    port map (
            O => \N__9755\,
            I => \N__9735\
        );

    \I__2156\ : InMux
    port map (
            O => \N__9754\,
            I => \N__9735\
        );

    \I__2155\ : InMux
    port map (
            O => \N__9753\,
            I => \N__9735\
        );

    \I__2154\ : InMux
    port map (
            O => \N__9752\,
            I => \N__9735\
        );

    \I__2153\ : Span4Mux_h
    port map (
            O => \N__9747\,
            I => \N__9730\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__9744\,
            I => \N__9730\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__9735\,
            I => \N__9727\
        );

    \I__2150\ : Span4Mux_v
    port map (
            O => \N__9730\,
            I => \N__9724\
        );

    \I__2149\ : Span4Mux_v
    port map (
            O => \N__9727\,
            I => \N__9721\
        );

    \I__2148\ : Span4Mux_v
    port map (
            O => \N__9724\,
            I => \N__9718\
        );

    \I__2147\ : Sp12to4
    port map (
            O => \N__9721\,
            I => \N__9715\
        );

    \I__2146\ : Sp12to4
    port map (
            O => \N__9718\,
            I => \N__9710\
        );

    \I__2145\ : Span12Mux_h
    port map (
            O => \N__9715\,
            I => \N__9710\
        );

    \I__2144\ : Odrv12
    port map (
            O => \N__9710\,
            I => \A_c_1\
        );

    \I__2143\ : CascadeMux
    port map (
            O => \N__9707\,
            I => \N__9703\
        );

    \I__2142\ : CascadeMux
    port map (
            O => \N__9706\,
            I => \N__9699\
        );

    \I__2141\ : InMux
    port map (
            O => \N__9703\,
            I => \N__9696\
        );

    \I__2140\ : InMux
    port map (
            O => \N__9702\,
            I => \N__9691\
        );

    \I__2139\ : InMux
    port map (
            O => \N__9699\,
            I => \N__9691\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__9696\,
            I => \N__9688\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__9691\,
            I => \N__9685\
        );

    \I__2136\ : Span4Mux_v
    port map (
            O => \N__9688\,
            I => \N__9675\
        );

    \I__2135\ : Span4Mux_v
    port map (
            O => \N__9685\,
            I => \N__9672\
        );

    \I__2134\ : InMux
    port map (
            O => \N__9684\,
            I => \N__9669\
        );

    \I__2133\ : InMux
    port map (
            O => \N__9683\,
            I => \N__9666\
        );

    \I__2132\ : InMux
    port map (
            O => \N__9682\,
            I => \N__9663\
        );

    \I__2131\ : InMux
    port map (
            O => \N__9681\,
            I => \N__9654\
        );

    \I__2130\ : InMux
    port map (
            O => \N__9680\,
            I => \N__9654\
        );

    \I__2129\ : InMux
    port map (
            O => \N__9679\,
            I => \N__9654\
        );

    \I__2128\ : InMux
    port map (
            O => \N__9678\,
            I => \N__9654\
        );

    \I__2127\ : Sp12to4
    port map (
            O => \N__9675\,
            I => \N__9647\
        );

    \I__2126\ : Sp12to4
    port map (
            O => \N__9672\,
            I => \N__9647\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__9669\,
            I => \N__9647\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__9666\,
            I => \N__9640\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__9663\,
            I => \N__9640\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__9654\,
            I => \N__9640\
        );

    \I__2121\ : Span12Mux_h
    port map (
            O => \N__9647\,
            I => \N__9637\
        );

    \I__2120\ : Span12Mux_v
    port map (
            O => \N__9640\,
            I => \N__9634\
        );

    \I__2119\ : Span12Mux_v
    port map (
            O => \N__9637\,
            I => \N__9629\
        );

    \I__2118\ : Span12Mux_h
    port map (
            O => \N__9634\,
            I => \N__9629\
        );

    \I__2117\ : Odrv12
    port map (
            O => \N__9629\,
            I => \SIZ_c_1\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__9626\,
            I => \N__9618\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__9625\,
            I => \N__9615\
        );

    \I__2114\ : InMux
    port map (
            O => \N__9624\,
            I => \N__9608\
        );

    \I__2113\ : CascadeMux
    port map (
            O => \N__9623\,
            I => \N__9605\
        );

    \I__2112\ : InMux
    port map (
            O => \N__9622\,
            I => \N__9596\
        );

    \I__2111\ : InMux
    port map (
            O => \N__9621\,
            I => \N__9596\
        );

    \I__2110\ : InMux
    port map (
            O => \N__9618\,
            I => \N__9596\
        );

    \I__2109\ : InMux
    port map (
            O => \N__9615\,
            I => \N__9596\
        );

    \I__2108\ : InMux
    port map (
            O => \N__9614\,
            I => \N__9593\
        );

    \I__2107\ : InMux
    port map (
            O => \N__9613\,
            I => \N__9590\
        );

    \I__2106\ : InMux
    port map (
            O => \N__9612\,
            I => \N__9585\
        );

    \I__2105\ : InMux
    port map (
            O => \N__9611\,
            I => \N__9585\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__9608\,
            I => \N__9582\
        );

    \I__2103\ : InMux
    port map (
            O => \N__9605\,
            I => \N__9579\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__9596\,
            I => \N__9576\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__9593\,
            I => \N__9571\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__9590\,
            I => \N__9571\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__9585\,
            I => \N__9568\
        );

    \I__2098\ : Span4Mux_v
    port map (
            O => \N__9582\,
            I => \N__9563\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__9579\,
            I => \N__9563\
        );

    \I__2096\ : Span4Mux_v
    port map (
            O => \N__9576\,
            I => \N__9558\
        );

    \I__2095\ : Span4Mux_v
    port map (
            O => \N__9571\,
            I => \N__9558\
        );

    \I__2094\ : Span4Mux_v
    port map (
            O => \N__9568\,
            I => \N__9555\
        );

    \I__2093\ : Span4Mux_h
    port map (
            O => \N__9563\,
            I => \N__9552\
        );

    \I__2092\ : Sp12to4
    port map (
            O => \N__9558\,
            I => \N__9549\
        );

    \I__2091\ : Span4Mux_v
    port map (
            O => \N__9555\,
            I => \N__9546\
        );

    \I__2090\ : Span4Mux_v
    port map (
            O => \N__9552\,
            I => \N__9543\
        );

    \I__2089\ : Span12Mux_h
    port map (
            O => \N__9549\,
            I => \N__9536\
        );

    \I__2088\ : Sp12to4
    port map (
            O => \N__9546\,
            I => \N__9536\
        );

    \I__2087\ : Sp12to4
    port map (
            O => \N__9543\,
            I => \N__9536\
        );

    \I__2086\ : Odrv12
    port map (
            O => \N__9536\,
            I => \A_c_0\
        );

    \I__2085\ : CascadeMux
    port map (
            O => \N__9533\,
            I => \N__9529\
        );

    \I__2084\ : InMux
    port map (
            O => \N__9532\,
            I => \N__9525\
        );

    \I__2083\ : InMux
    port map (
            O => \N__9529\,
            I => \N__9522\
        );

    \I__2082\ : CascadeMux
    port map (
            O => \N__9528\,
            I => \N__9516\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__9525\,
            I => \N__9510\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__9522\,
            I => \N__9510\
        );

    \I__2079\ : CascadeMux
    port map (
            O => \N__9521\,
            I => \N__9507\
        );

    \I__2078\ : CascadeMux
    port map (
            O => \N__9520\,
            I => \N__9504\
        );

    \I__2077\ : InMux
    port map (
            O => \N__9519\,
            I => \N__9499\
        );

    \I__2076\ : InMux
    port map (
            O => \N__9516\,
            I => \N__9494\
        );

    \I__2075\ : InMux
    port map (
            O => \N__9515\,
            I => \N__9494\
        );

    \I__2074\ : Span4Mux_v
    port map (
            O => \N__9510\,
            I => \N__9491\
        );

    \I__2073\ : InMux
    port map (
            O => \N__9507\,
            I => \N__9482\
        );

    \I__2072\ : InMux
    port map (
            O => \N__9504\,
            I => \N__9482\
        );

    \I__2071\ : InMux
    port map (
            O => \N__9503\,
            I => \N__9482\
        );

    \I__2070\ : InMux
    port map (
            O => \N__9502\,
            I => \N__9482\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__9499\,
            I => \N__9479\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__9494\,
            I => \N__9476\
        );

    \I__2067\ : Span4Mux_v
    port map (
            O => \N__9491\,
            I => \N__9470\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__9482\,
            I => \N__9470\
        );

    \I__2065\ : Span4Mux_v
    port map (
            O => \N__9479\,
            I => \N__9467\
        );

    \I__2064\ : Span4Mux_v
    port map (
            O => \N__9476\,
            I => \N__9464\
        );

    \I__2063\ : InMux
    port map (
            O => \N__9475\,
            I => \N__9461\
        );

    \I__2062\ : Span4Mux_h
    port map (
            O => \N__9470\,
            I => \N__9458\
        );

    \I__2061\ : Sp12to4
    port map (
            O => \N__9467\,
            I => \N__9451\
        );

    \I__2060\ : Sp12to4
    port map (
            O => \N__9464\,
            I => \N__9451\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__9461\,
            I => \N__9451\
        );

    \I__2058\ : Span4Mux_v
    port map (
            O => \N__9458\,
            I => \N__9448\
        );

    \I__2057\ : Span12Mux_h
    port map (
            O => \N__9451\,
            I => \N__9445\
        );

    \I__2056\ : Span4Mux_h
    port map (
            O => \N__9448\,
            I => \N__9442\
        );

    \I__2055\ : Span12Mux_v
    port map (
            O => \N__9445\,
            I => \N__9439\
        );

    \I__2054\ : Sp12to4
    port map (
            O => \N__9442\,
            I => \N__9436\
        );

    \I__2053\ : Odrv12
    port map (
            O => \N__9439\,
            I => \SIZ_c_0\
        );

    \I__2052\ : Odrv12
    port map (
            O => \N__9436\,
            I => \SIZ_c_0\
        );

    \I__2051\ : IoInMux
    port map (
            O => \N__9431\,
            I => \N__9428\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__9428\,
            I => \N__9425\
        );

    \I__2049\ : Span4Mux_s2_v
    port map (
            O => \N__9425\,
            I => \N__9422\
        );

    \I__2048\ : Span4Mux_h
    port map (
            O => \N__9422\,
            I => \N__9419\
        );

    \I__2047\ : Span4Mux_v
    port map (
            O => \N__9419\,
            I => \N__9416\
        );

    \I__2046\ : Odrv4
    port map (
            O => \N__9416\,
            I => \N_324_i\
        );

    \I__2045\ : IoInMux
    port map (
            O => \N__9413\,
            I => \N__9410\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__9410\,
            I => \N__9407\
        );

    \I__2043\ : Span4Mux_s2_h
    port map (
            O => \N__9407\,
            I => \N__9404\
        );

    \I__2042\ : Span4Mux_v
    port map (
            O => \N__9404\,
            I => \N__9401\
        );

    \I__2041\ : Sp12to4
    port map (
            O => \N__9401\,
            I => \N__9398\
        );

    \I__2040\ : Span12Mux_h
    port map (
            O => \N__9398\,
            I => \N__9395\
        );

    \I__2039\ : Odrv12
    port map (
            O => \N__9395\,
            I => \WEn_c\
        );

    \I__2038\ : InMux
    port map (
            O => \N__9392\,
            I => \N__9379\
        );

    \I__2037\ : InMux
    port map (
            O => \N__9391\,
            I => \N__9379\
        );

    \I__2036\ : InMux
    port map (
            O => \N__9390\,
            I => \N__9379\
        );

    \I__2035\ : InMux
    port map (
            O => \N__9389\,
            I => \N__9376\
        );

    \I__2034\ : InMux
    port map (
            O => \N__9388\,
            I => \N__9369\
        );

    \I__2033\ : InMux
    port map (
            O => \N__9387\,
            I => \N__9369\
        );

    \I__2032\ : InMux
    port map (
            O => \N__9386\,
            I => \N__9369\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__9379\,
            I => \N__9365\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__9376\,
            I => \N__9360\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__9369\,
            I => \N__9360\
        );

    \I__2028\ : InMux
    port map (
            O => \N__9368\,
            I => \N__9356\
        );

    \I__2027\ : Span4Mux_h
    port map (
            O => \N__9365\,
            I => \N__9352\
        );

    \I__2026\ : Span4Mux_h
    port map (
            O => \N__9360\,
            I => \N__9349\
        );

    \I__2025\ : InMux
    port map (
            O => \N__9359\,
            I => \N__9346\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__9356\,
            I => \N__9343\
        );

    \I__2023\ : InMux
    port map (
            O => \N__9355\,
            I => \N__9340\
        );

    \I__2022\ : Odrv4
    port map (
            O => \N__9352\,
            I => \U712_CHIP_RAM.N_305\
        );

    \I__2021\ : Odrv4
    port map (
            O => \N__9349\,
            I => \U712_CHIP_RAM.N_305\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__9346\,
            I => \U712_CHIP_RAM.N_305\
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__9343\,
            I => \U712_CHIP_RAM.N_305\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__9340\,
            I => \U712_CHIP_RAM.N_305\
        );

    \I__2017\ : CascadeMux
    port map (
            O => \N__9329\,
            I => \N__9321\
        );

    \I__2016\ : CascadeMux
    port map (
            O => \N__9328\,
            I => \N__9318\
        );

    \I__2015\ : CascadeMux
    port map (
            O => \N__9327\,
            I => \N__9315\
        );

    \I__2014\ : CascadeMux
    port map (
            O => \N__9326\,
            I => \N__9312\
        );

    \I__2013\ : CascadeMux
    port map (
            O => \N__9325\,
            I => \N__9308\
        );

    \I__2012\ : CascadeMux
    port map (
            O => \N__9324\,
            I => \N__9305\
        );

    \I__2011\ : InMux
    port map (
            O => \N__9321\,
            I => \N__9302\
        );

    \I__2010\ : InMux
    port map (
            O => \N__9318\,
            I => \N__9297\
        );

    \I__2009\ : InMux
    port map (
            O => \N__9315\,
            I => \N__9297\
        );

    \I__2008\ : InMux
    port map (
            O => \N__9312\,
            I => \N__9292\
        );

    \I__2007\ : InMux
    port map (
            O => \N__9311\,
            I => \N__9292\
        );

    \I__2006\ : InMux
    port map (
            O => \N__9308\,
            I => \N__9289\
        );

    \I__2005\ : InMux
    port map (
            O => \N__9305\,
            I => \N__9286\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__9302\,
            I => \N__9283\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__9297\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__9292\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__9289\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__9286\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__1999\ : Odrv4
    port map (
            O => \N__9283\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__1998\ : IoInMux
    port map (
            O => \N__9272\,
            I => \N__9269\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__9269\,
            I => \N__9266\
        );

    \I__1996\ : IoSpan4Mux
    port map (
            O => \N__9266\,
            I => \N__9263\
        );

    \I__1995\ : Sp12to4
    port map (
            O => \N__9263\,
            I => \N__9260\
        );

    \I__1994\ : Span12Mux_s1_h
    port map (
            O => \N__9260\,
            I => \N__9257\
        );

    \I__1993\ : Span12Mux_h
    port map (
            O => \N__9257\,
            I => \N__9254\
        );

    \I__1992\ : Odrv12
    port map (
            O => \N__9254\,
            I => \CMA_c_3\
        );

    \I__1991\ : CEMux
    port map (
            O => \N__9251\,
            I => \N__9246\
        );

    \I__1990\ : CEMux
    port map (
            O => \N__9250\,
            I => \N__9241\
        );

    \I__1989\ : CEMux
    port map (
            O => \N__9249\,
            I => \N__9237\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__9246\,
            I => \N__9234\
        );

    \I__1987\ : CEMux
    port map (
            O => \N__9245\,
            I => \N__9230\
        );

    \I__1986\ : CEMux
    port map (
            O => \N__9244\,
            I => \N__9227\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__9241\,
            I => \N__9224\
        );

    \I__1984\ : CEMux
    port map (
            O => \N__9240\,
            I => \N__9221\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__9237\,
            I => \N__9216\
        );

    \I__1982\ : Span4Mux_v
    port map (
            O => \N__9234\,
            I => \N__9216\
        );

    \I__1981\ : CEMux
    port map (
            O => \N__9233\,
            I => \N__9213\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__9230\,
            I => \N__9210\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__9227\,
            I => \N__9207\
        );

    \I__1978\ : Span4Mux_v
    port map (
            O => \N__9224\,
            I => \N__9204\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__9221\,
            I => \N__9199\
        );

    \I__1976\ : Span4Mux_h
    port map (
            O => \N__9216\,
            I => \N__9199\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__9213\,
            I => \N__9196\
        );

    \I__1974\ : Sp12to4
    port map (
            O => \N__9210\,
            I => \N__9193\
        );

    \I__1973\ : Span4Mux_h
    port map (
            O => \N__9207\,
            I => \N__9190\
        );

    \I__1972\ : Odrv4
    port map (
            O => \N__9204\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__1971\ : Odrv4
    port map (
            O => \N__9199\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__1970\ : Odrv4
    port map (
            O => \N__9196\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__1969\ : Odrv12
    port map (
            O => \N__9193\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__1968\ : Odrv4
    port map (
            O => \N__9190\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__1967\ : InMux
    port map (
            O => \N__9179\,
            I => \N__9175\
        );

    \I__1966\ : InMux
    port map (
            O => \N__9178\,
            I => \N__9172\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__9175\,
            I => \N__9169\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__9172\,
            I => \N__9166\
        );

    \I__1963\ : Span4Mux_h
    port map (
            O => \N__9169\,
            I => \N__9160\
        );

    \I__1962\ : Span4Mux_h
    port map (
            O => \N__9166\,
            I => \N__9157\
        );

    \I__1961\ : InMux
    port map (
            O => \N__9165\,
            I => \N__9154\
        );

    \I__1960\ : InMux
    port map (
            O => \N__9164\,
            I => \N__9149\
        );

    \I__1959\ : InMux
    port map (
            O => \N__9163\,
            I => \N__9149\
        );

    \I__1958\ : Odrv4
    port map (
            O => \N__9160\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__9157\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__9154\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__9149\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1954\ : InMux
    port map (
            O => \N__9140\,
            I => \N__9137\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__9137\,
            I => \U712_CHIP_RAM.CMA_5_i_0_9\
        );

    \I__1952\ : InMux
    port map (
            O => \N__9134\,
            I => \N__9131\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__9131\,
            I => \N__9128\
        );

    \I__1950\ : Odrv12
    port map (
            O => \N__9128\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\
        );

    \I__1949\ : CascadeMux
    port map (
            O => \N__9125\,
            I => \N__9116\
        );

    \I__1948\ : CascadeMux
    port map (
            O => \N__9124\,
            I => \N__9112\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__9123\,
            I => \N__9109\
        );

    \I__1946\ : InMux
    port map (
            O => \N__9122\,
            I => \N__9105\
        );

    \I__1945\ : InMux
    port map (
            O => \N__9121\,
            I => \N__9098\
        );

    \I__1944\ : InMux
    port map (
            O => \N__9120\,
            I => \N__9098\
        );

    \I__1943\ : InMux
    port map (
            O => \N__9119\,
            I => \N__9098\
        );

    \I__1942\ : InMux
    port map (
            O => \N__9116\,
            I => \N__9095\
        );

    \I__1941\ : InMux
    port map (
            O => \N__9115\,
            I => \N__9092\
        );

    \I__1940\ : InMux
    port map (
            O => \N__9112\,
            I => \N__9089\
        );

    \I__1939\ : InMux
    port map (
            O => \N__9109\,
            I => \N__9086\
        );

    \I__1938\ : InMux
    port map (
            O => \N__9108\,
            I => \N__9076\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__9105\,
            I => \N__9070\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__9098\,
            I => \N__9067\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__9095\,
            I => \N__9058\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__9092\,
            I => \N__9058\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__9089\,
            I => \N__9058\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__9086\,
            I => \N__9058\
        );

    \I__1931\ : InMux
    port map (
            O => \N__9085\,
            I => \N__9055\
        );

    \I__1930\ : InMux
    port map (
            O => \N__9084\,
            I => \N__9052\
        );

    \I__1929\ : InMux
    port map (
            O => \N__9083\,
            I => \N__9049\
        );

    \I__1928\ : InMux
    port map (
            O => \N__9082\,
            I => \N__9044\
        );

    \I__1927\ : InMux
    port map (
            O => \N__9081\,
            I => \N__9044\
        );

    \I__1926\ : InMux
    port map (
            O => \N__9080\,
            I => \N__9039\
        );

    \I__1925\ : InMux
    port map (
            O => \N__9079\,
            I => \N__9039\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__9076\,
            I => \N__9036\
        );

    \I__1923\ : InMux
    port map (
            O => \N__9075\,
            I => \N__9032\
        );

    \I__1922\ : InMux
    port map (
            O => \N__9074\,
            I => \N__9027\
        );

    \I__1921\ : InMux
    port map (
            O => \N__9073\,
            I => \N__9027\
        );

    \I__1920\ : Span4Mux_h
    port map (
            O => \N__9070\,
            I => \N__9024\
        );

    \I__1919\ : Span4Mux_h
    port map (
            O => \N__9067\,
            I => \N__9021\
        );

    \I__1918\ : Span4Mux_h
    port map (
            O => \N__9058\,
            I => \N__9018\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__9055\,
            I => \N__9015\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__9052\,
            I => \N__9008\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__9049\,
            I => \N__9008\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__9044\,
            I => \N__9008\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__9039\,
            I => \N__9003\
        );

    \I__1912\ : Span4Mux_v
    port map (
            O => \N__9036\,
            I => \N__9003\
        );

    \I__1911\ : CascadeMux
    port map (
            O => \N__9035\,
            I => \N__8999\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__9032\,
            I => \N__8994\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__9027\,
            I => \N__8991\
        );

    \I__1908\ : Span4Mux_h
    port map (
            O => \N__9024\,
            I => \N__8986\
        );

    \I__1907\ : Span4Mux_h
    port map (
            O => \N__9021\,
            I => \N__8986\
        );

    \I__1906\ : Span4Mux_h
    port map (
            O => \N__9018\,
            I => \N__8983\
        );

    \I__1905\ : Span4Mux_v
    port map (
            O => \N__9015\,
            I => \N__8976\
        );

    \I__1904\ : Span4Mux_v
    port map (
            O => \N__9008\,
            I => \N__8976\
        );

    \I__1903\ : Span4Mux_h
    port map (
            O => \N__9003\,
            I => \N__8976\
        );

    \I__1902\ : InMux
    port map (
            O => \N__9002\,
            I => \N__8969\
        );

    \I__1901\ : InMux
    port map (
            O => \N__8999\,
            I => \N__8969\
        );

    \I__1900\ : InMux
    port map (
            O => \N__8998\,
            I => \N__8969\
        );

    \I__1899\ : InMux
    port map (
            O => \N__8997\,
            I => \N__8966\
        );

    \I__1898\ : Odrv4
    port map (
            O => \N__8994\,
            I => \CPU_CYCLEm\
        );

    \I__1897\ : Odrv4
    port map (
            O => \N__8991\,
            I => \CPU_CYCLEm\
        );

    \I__1896\ : Odrv4
    port map (
            O => \N__8986\,
            I => \CPU_CYCLEm\
        );

    \I__1895\ : Odrv4
    port map (
            O => \N__8983\,
            I => \CPU_CYCLEm\
        );

    \I__1894\ : Odrv4
    port map (
            O => \N__8976\,
            I => \CPU_CYCLEm\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__8969\,
            I => \CPU_CYCLEm\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__8966\,
            I => \CPU_CYCLEm\
        );

    \I__1891\ : InMux
    port map (
            O => \N__8951\,
            I => \N__8948\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__8948\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__1889\ : InMux
    port map (
            O => \N__8945\,
            I => \N__8942\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__8942\,
            I => \N__8939\
        );

    \I__1887\ : Odrv4
    port map (
            O => \N__8939\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__1886\ : InMux
    port map (
            O => \N__8936\,
            I => \N__8932\
        );

    \I__1885\ : InMux
    port map (
            O => \N__8935\,
            I => \N__8929\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__8932\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__8929\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__1882\ : InMux
    port map (
            O => \N__8924\,
            I => \N__8921\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__8921\,
            I => \N__8918\
        );

    \I__1880\ : Odrv12
    port map (
            O => \N__8918\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_7\
        );

    \I__1879\ : InMux
    port map (
            O => \N__8915\,
            I => \N__8910\
        );

    \I__1878\ : InMux
    port map (
            O => \N__8914\,
            I => \N__8907\
        );

    \I__1877\ : InMux
    port map (
            O => \N__8913\,
            I => \N__8904\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__8910\,
            I => \U712_REG_SM.N_319\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__8907\,
            I => \U712_REG_SM.N_319\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__8904\,
            I => \U712_REG_SM.N_319\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8897\,
            I => \N__8893\
        );

    \I__1872\ : InMux
    port map (
            O => \N__8896\,
            I => \N__8890\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__8893\,
            I => \N__8885\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__8890\,
            I => \N__8882\
        );

    \I__1869\ : InMux
    port map (
            O => \N__8889\,
            I => \N__8879\
        );

    \I__1868\ : InMux
    port map (
            O => \N__8888\,
            I => \N__8876\
        );

    \I__1867\ : Span4Mux_h
    port map (
            O => \N__8885\,
            I => \N__8873\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__8882\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__8879\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__8876\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__1863\ : Odrv4
    port map (
            O => \N__8873\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__8864\,
            I => \U712_REG_SM.N_318_cascade_\
        );

    \I__1861\ : InMux
    port map (
            O => \N__8861\,
            I => \N__8855\
        );

    \I__1860\ : InMux
    port map (
            O => \N__8860\,
            I => \N__8850\
        );

    \I__1859\ : InMux
    port map (
            O => \N__8859\,
            I => \N__8850\
        );

    \I__1858\ : InMux
    port map (
            O => \N__8858\,
            I => \N__8847\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__8855\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__8850\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__8847\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1854\ : IoInMux
    port map (
            O => \N__8840\,
            I => \N__8837\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__8837\,
            I => \N__8834\
        );

    \I__1852\ : Span4Mux_s0_v
    port map (
            O => \N__8834\,
            I => \N__8831\
        );

    \I__1851\ : Span4Mux_v
    port map (
            O => \N__8831\,
            I => \N__8827\
        );

    \I__1850\ : IoInMux
    port map (
            O => \N__8830\,
            I => \N__8824\
        );

    \I__1849\ : Span4Mux_v
    port map (
            O => \N__8827\,
            I => \N__8821\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__8824\,
            I => \N__8818\
        );

    \I__1847\ : Sp12to4
    port map (
            O => \N__8821\,
            I => \N__8815\
        );

    \I__1846\ : Span12Mux_s8_v
    port map (
            O => \N__8818\,
            I => \N__8812\
        );

    \I__1845\ : Span12Mux_h
    port map (
            O => \N__8815\,
            I => \N__8805\
        );

    \I__1844\ : Span12Mux_h
    port map (
            O => \N__8812\,
            I => \N__8805\
        );

    \I__1843\ : InMux
    port map (
            O => \N__8811\,
            I => \N__8802\
        );

    \I__1842\ : InMux
    port map (
            O => \N__8810\,
            I => \N__8799\
        );

    \I__1841\ : Odrv12
    port map (
            O => \N__8805\,
            I => \BLSn_c\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__8802\,
            I => \BLSn_c\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__8799\,
            I => \BLSn_c\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8792\,
            I => \N__8789\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__8789\,
            I => \U712_REG_SM.REGENn_e_1\
        );

    \I__1836\ : IoInMux
    port map (
            O => \N__8786\,
            I => \N__8783\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__8783\,
            I => \N__8780\
        );

    \I__1834\ : Span4Mux_s0_v
    port map (
            O => \N__8780\,
            I => \N__8777\
        );

    \I__1833\ : Span4Mux_v
    port map (
            O => \N__8777\,
            I => \N__8774\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__8774\,
            I => \N_326_i\
        );

    \I__1831\ : InMux
    port map (
            O => \N__8771\,
            I => \N__8768\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8768\,
            I => \N__8765\
        );

    \I__1829\ : Span4Mux_v
    port map (
            O => \N__8765\,
            I => \N__8762\
        );

    \I__1828\ : Span4Mux_v
    port map (
            O => \N__8762\,
            I => \N__8759\
        );

    \I__1827\ : Sp12to4
    port map (
            O => \N__8759\,
            I => \N__8756\
        );

    \I__1826\ : Span12Mux_h
    port map (
            O => \N__8756\,
            I => \N__8753\
        );

    \I__1825\ : Odrv12
    port map (
            O => \N__8753\,
            I => \A_c_19\
        );

    \I__1824\ : IoInMux
    port map (
            O => \N__8750\,
            I => \N__8747\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__8747\,
            I => \N__8744\
        );

    \I__1822\ : IoSpan4Mux
    port map (
            O => \N__8744\,
            I => \N__8741\
        );

    \I__1821\ : Span4Mux_s0_h
    port map (
            O => \N__8741\,
            I => \N__8738\
        );

    \I__1820\ : Sp12to4
    port map (
            O => \N__8738\,
            I => \N__8735\
        );

    \I__1819\ : Span12Mux_h
    port map (
            O => \N__8735\,
            I => \N__8732\
        );

    \I__1818\ : Odrv12
    port map (
            O => \N__8732\,
            I => \CMA_c_9\
        );

    \I__1817\ : InMux
    port map (
            O => \N__8729\,
            I => \N__8726\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__8726\,
            I => \N__8723\
        );

    \I__1815\ : Odrv4
    port map (
            O => \N__8723\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__1814\ : InMux
    port map (
            O => \N__8720\,
            I => \N__8717\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__8717\,
            I => \N__8714\
        );

    \I__1812\ : Odrv4
    port map (
            O => \N__8714\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__1811\ : InMux
    port map (
            O => \N__8711\,
            I => \N__8708\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__8708\,
            I => \N__8705\
        );

    \I__1809\ : Odrv12
    port map (
            O => \N__8705\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__1808\ : InMux
    port map (
            O => \N__8702\,
            I => \N__8699\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__8699\,
            I => \N__8696\
        );

    \I__1806\ : Span4Mux_h
    port map (
            O => \N__8696\,
            I => \N__8693\
        );

    \I__1805\ : Odrv4
    port map (
            O => \N__8693\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__1804\ : InMux
    port map (
            O => \N__8690\,
            I => \N__8687\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__8687\,
            I => \N__8684\
        );

    \I__1802\ : Odrv4
    port map (
            O => \N__8684\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8681\,
            I => \N__8678\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__8678\,
            I => \N__8675\
        );

    \I__1799\ : Span4Mux_h
    port map (
            O => \N__8675\,
            I => \N__8672\
        );

    \I__1798\ : Odrv4
    port map (
            O => \N__8672\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__1797\ : InMux
    port map (
            O => \N__8669\,
            I => \N__8661\
        );

    \I__1796\ : InMux
    port map (
            O => \N__8668\,
            I => \N__8661\
        );

    \I__1795\ : InMux
    port map (
            O => \N__8667\,
            I => \N__8658\
        );

    \I__1794\ : InMux
    port map (
            O => \N__8666\,
            I => \N__8655\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__8661\,
            I => \N__8652\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__8658\,
            I => \N__8649\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__8655\,
            I => \N__8646\
        );

    \I__1790\ : Span4Mux_h
    port map (
            O => \N__8652\,
            I => \N__8643\
        );

    \I__1789\ : Span4Mux_h
    port map (
            O => \N__8649\,
            I => \N__8640\
        );

    \I__1788\ : Span12Mux_v
    port map (
            O => \N__8646\,
            I => \N__8637\
        );

    \I__1787\ : Sp12to4
    port map (
            O => \N__8643\,
            I => \N__8634\
        );

    \I__1786\ : Span4Mux_v
    port map (
            O => \N__8640\,
            I => \N__8631\
        );

    \I__1785\ : Span12Mux_h
    port map (
            O => \N__8637\,
            I => \N__8628\
        );

    \I__1784\ : Span12Mux_v
    port map (
            O => \N__8634\,
            I => \N__8623\
        );

    \I__1783\ : Sp12to4
    port map (
            O => \N__8631\,
            I => \N__8623\
        );

    \I__1782\ : Odrv12
    port map (
            O => \N__8628\,
            I => \DRA_c_6\
        );

    \I__1781\ : Odrv12
    port map (
            O => \N__8623\,
            I => \DRA_c_6\
        );

    \I__1780\ : InMux
    port map (
            O => \N__8618\,
            I => \N__8615\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__8615\,
            I => \N__8612\
        );

    \I__1778\ : Span4Mux_h
    port map (
            O => \N__8612\,
            I => \N__8609\
        );

    \I__1777\ : Span4Mux_v
    port map (
            O => \N__8609\,
            I => \N__8606\
        );

    \I__1776\ : Odrv4
    port map (
            O => \N__8606\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__1775\ : InMux
    port map (
            O => \N__8603\,
            I => \N__8599\
        );

    \I__1774\ : IoInMux
    port map (
            O => \N__8602\,
            I => \N__8596\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__8599\,
            I => \N__8593\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__8596\,
            I => \N__8590\
        );

    \I__1771\ : Span4Mux_v
    port map (
            O => \N__8593\,
            I => \N__8587\
        );

    \I__1770\ : IoSpan4Mux
    port map (
            O => \N__8590\,
            I => \N__8584\
        );

    \I__1769\ : Sp12to4
    port map (
            O => \N__8587\,
            I => \N__8581\
        );

    \I__1768\ : IoSpan4Mux
    port map (
            O => \N__8584\,
            I => \N__8578\
        );

    \I__1767\ : Span12Mux_h
    port map (
            O => \N__8581\,
            I => \N__8575\
        );

    \I__1766\ : IoSpan4Mux
    port map (
            O => \N__8578\,
            I => \N__8572\
        );

    \I__1765\ : Odrv12
    port map (
            O => \N__8575\,
            I => \C1_c\
        );

    \I__1764\ : Odrv4
    port map (
            O => \N__8572\,
            I => \C1_c\
        );

    \I__1763\ : InMux
    port map (
            O => \N__8567\,
            I => \N__8564\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__8564\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1761\ : InMux
    port map (
            O => \N__8561\,
            I => \N__8558\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__8558\,
            I => \N__8555\
        );

    \I__1759\ : Span4Mux_v
    port map (
            O => \N__8555\,
            I => \N__8552\
        );

    \I__1758\ : Odrv4
    port map (
            O => \N__8552\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__1757\ : IoInMux
    port map (
            O => \N__8549\,
            I => \N__8546\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__8546\,
            I => \N__8543\
        );

    \I__1755\ : Span4Mux_s1_v
    port map (
            O => \N__8543\,
            I => \N__8540\
        );

    \I__1754\ : Span4Mux_v
    port map (
            O => \N__8540\,
            I => \N__8537\
        );

    \I__1753\ : Span4Mux_v
    port map (
            O => \N__8537\,
            I => \N__8534\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__8534\,
            I => \CMA_c_0\
        );

    \I__1751\ : IoInMux
    port map (
            O => \N__8531\,
            I => \N__8528\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__8528\,
            I => \N__8525\
        );

    \I__1749\ : Span4Mux_s0_v
    port map (
            O => \N__8525\,
            I => \N__8522\
        );

    \I__1748\ : Sp12to4
    port map (
            O => \N__8522\,
            I => \N__8519\
        );

    \I__1747\ : Span12Mux_h
    port map (
            O => \N__8519\,
            I => \N__8516\
        );

    \I__1746\ : Odrv12
    port map (
            O => \N__8516\,
            I => \CMA_c_10\
        );

    \I__1745\ : InMux
    port map (
            O => \N__8513\,
            I => \N__8510\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__8510\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__1743\ : IoInMux
    port map (
            O => \N__8507\,
            I => \N__8504\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__8504\,
            I => \N__8501\
        );

    \I__1741\ : IoSpan4Mux
    port map (
            O => \N__8501\,
            I => \N__8498\
        );

    \I__1740\ : IoSpan4Mux
    port map (
            O => \N__8498\,
            I => \N__8495\
        );

    \I__1739\ : Span4Mux_s3_h
    port map (
            O => \N__8495\,
            I => \N__8492\
        );

    \I__1738\ : Sp12to4
    port map (
            O => \N__8492\,
            I => \N__8489\
        );

    \I__1737\ : Odrv12
    port map (
            O => \N__8489\,
            I => \CMA_c_6\
        );

    \I__1736\ : InMux
    port map (
            O => \N__8486\,
            I => \N__8483\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__8483\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\
        );

    \I__1734\ : IoInMux
    port map (
            O => \N__8480\,
            I => \N__8477\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__8477\,
            I => \N__8474\
        );

    \I__1732\ : IoSpan4Mux
    port map (
            O => \N__8474\,
            I => \N__8471\
        );

    \I__1731\ : Span4Mux_s2_h
    port map (
            O => \N__8471\,
            I => \N__8468\
        );

    \I__1730\ : Span4Mux_v
    port map (
            O => \N__8468\,
            I => \N__8465\
        );

    \I__1729\ : Span4Mux_h
    port map (
            O => \N__8465\,
            I => \N__8462\
        );

    \I__1728\ : Span4Mux_h
    port map (
            O => \N__8462\,
            I => \N__8459\
        );

    \I__1727\ : Odrv4
    port map (
            O => \N__8459\,
            I => \CMA_c_8\
        );

    \I__1726\ : InMux
    port map (
            O => \N__8456\,
            I => \N__8453\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__8453\,
            I => \N__8450\
        );

    \I__1724\ : Odrv4
    port map (
            O => \N__8450\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__1723\ : IoInMux
    port map (
            O => \N__8447\,
            I => \N__8444\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__8444\,
            I => \N__8441\
        );

    \I__1721\ : Span4Mux_s2_h
    port map (
            O => \N__8441\,
            I => \N__8438\
        );

    \I__1720\ : Sp12to4
    port map (
            O => \N__8438\,
            I => \N__8435\
        );

    \I__1719\ : Span12Mux_s11_v
    port map (
            O => \N__8435\,
            I => \N__8432\
        );

    \I__1718\ : Span12Mux_h
    port map (
            O => \N__8432\,
            I => \N__8429\
        );

    \I__1717\ : Odrv12
    port map (
            O => \N__8429\,
            I => \CMA_c_4\
        );

    \I__1716\ : InMux
    port map (
            O => \N__8426\,
            I => \N__8423\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__8423\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__1714\ : IoInMux
    port map (
            O => \N__8420\,
            I => \N__8417\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__8417\,
            I => \N__8414\
        );

    \I__1712\ : Span4Mux_s2_h
    port map (
            O => \N__8414\,
            I => \N__8411\
        );

    \I__1711\ : Sp12to4
    port map (
            O => \N__8411\,
            I => \N__8408\
        );

    \I__1710\ : Span12Mux_s10_v
    port map (
            O => \N__8408\,
            I => \N__8405\
        );

    \I__1709\ : Odrv12
    port map (
            O => \N__8405\,
            I => \CMA_c_7\
        );

    \I__1708\ : CascadeMux
    port map (
            O => \N__8402\,
            I => \U712_REG_SM.REG_CYCLE_5_iv_0_0_cascade_\
        );

    \I__1707\ : InMux
    port map (
            O => \N__8399\,
            I => \N__8396\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__8396\,
            I => \U712_REG_SM.N_409\
        );

    \I__1705\ : InMux
    port map (
            O => \N__8393\,
            I => \N__8390\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__8390\,
            I => \N__8387\
        );

    \I__1703\ : Span4Mux_v
    port map (
            O => \N__8387\,
            I => \N__8383\
        );

    \I__1702\ : InMux
    port map (
            O => \N__8386\,
            I => \N__8380\
        );

    \I__1701\ : Span4Mux_h
    port map (
            O => \N__8383\,
            I => \N__8375\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8380\,
            I => \N__8372\
        );

    \I__1699\ : InMux
    port map (
            O => \N__8379\,
            I => \N__8367\
        );

    \I__1698\ : InMux
    port map (
            O => \N__8378\,
            I => \N__8367\
        );

    \I__1697\ : Odrv4
    port map (
            O => \N__8375\,
            I => \REG_CYCLEm\
        );

    \I__1696\ : Odrv4
    port map (
            O => \N__8372\,
            I => \REG_CYCLEm\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__8367\,
            I => \REG_CYCLEm\
        );

    \I__1694\ : InMux
    port map (
            O => \N__8360\,
            I => \N__8357\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__8357\,
            I => \U712_REG_SM.STATE_COUNTsr_0\
        );

    \I__1692\ : CascadeMux
    port map (
            O => \N__8354\,
            I => \N__8351\
        );

    \I__1691\ : InMux
    port map (
            O => \N__8351\,
            I => \N__8348\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__8348\,
            I => \U712_REG_SM.N_328\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__8345\,
            I => \N__8341\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__8344\,
            I => \N__8338\
        );

    \I__1687\ : InMux
    port map (
            O => \N__8341\,
            I => \N__8335\
        );

    \I__1686\ : InMux
    port map (
            O => \N__8338\,
            I => \N__8326\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__8335\,
            I => \N__8323\
        );

    \I__1684\ : InMux
    port map (
            O => \N__8334\,
            I => \N__8320\
        );

    \I__1683\ : InMux
    port map (
            O => \N__8333\,
            I => \N__8311\
        );

    \I__1682\ : InMux
    port map (
            O => \N__8332\,
            I => \N__8311\
        );

    \I__1681\ : InMux
    port map (
            O => \N__8331\,
            I => \N__8311\
        );

    \I__1680\ : InMux
    port map (
            O => \N__8330\,
            I => \N__8311\
        );

    \I__1679\ : InMux
    port map (
            O => \N__8329\,
            I => \N__8308\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__8326\,
            I => \N__8305\
        );

    \I__1677\ : Span4Mux_h
    port map (
            O => \N__8323\,
            I => \N__8300\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__8320\,
            I => \N__8300\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__8311\,
            I => \N__8294\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__8308\,
            I => \N__8294\
        );

    \I__1673\ : Span4Mux_v
    port map (
            O => \N__8305\,
            I => \N__8289\
        );

    \I__1672\ : Span4Mux_h
    port map (
            O => \N__8300\,
            I => \N__8289\
        );

    \I__1671\ : InMux
    port map (
            O => \N__8299\,
            I => \N__8286\
        );

    \I__1670\ : Odrv4
    port map (
            O => \N__8294\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1669\ : Odrv4
    port map (
            O => \N__8289\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__8286\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1667\ : CascadeMux
    port map (
            O => \N__8279\,
            I => \U712_REG_SM.N_412_cascade_\
        );

    \I__1666\ : InMux
    port map (
            O => \N__8276\,
            I => \N__8271\
        );

    \I__1665\ : InMux
    port map (
            O => \N__8275\,
            I => \N__8266\
        );

    \I__1664\ : InMux
    port map (
            O => \N__8274\,
            I => \N__8266\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__8271\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_3\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__8266\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_3\
        );

    \I__1661\ : CascadeMux
    port map (
            O => \N__8261\,
            I => \U712_REG_SM.N_360_cascade_\
        );

    \I__1660\ : InMux
    port map (
            O => \N__8258\,
            I => \N__8255\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__8255\,
            I => \U712_REG_SM.N_320\
        );

    \I__1658\ : InMux
    port map (
            O => \N__8252\,
            I => \N__8245\
        );

    \I__1657\ : InMux
    port map (
            O => \N__8251\,
            I => \N__8245\
        );

    \I__1656\ : InMux
    port map (
            O => \N__8250\,
            I => \N__8242\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__8245\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__8242\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1653\ : IoInMux
    port map (
            O => \N__8237\,
            I => \N__8234\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__8234\,
            I => \N__8231\
        );

    \I__1651\ : IoSpan4Mux
    port map (
            O => \N__8231\,
            I => \N__8228\
        );

    \I__1650\ : Span4Mux_s3_h
    port map (
            O => \N__8228\,
            I => \N__8225\
        );

    \I__1649\ : Span4Mux_v
    port map (
            O => \N__8225\,
            I => \N__8221\
        );

    \I__1648\ : InMux
    port map (
            O => \N__8224\,
            I => \N__8218\
        );

    \I__1647\ : Span4Mux_h
    port map (
            O => \N__8221\,
            I => \N__8215\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__8218\,
            I => \N__8212\
        );

    \I__1645\ : Sp12to4
    port map (
            O => \N__8215\,
            I => \N__8209\
        );

    \I__1644\ : Span4Mux_v
    port map (
            O => \N__8212\,
            I => \N__8206\
        );

    \I__1643\ : Span12Mux_h
    port map (
            O => \N__8209\,
            I => \N__8201\
        );

    \I__1642\ : Sp12to4
    port map (
            O => \N__8206\,
            I => \N__8201\
        );

    \I__1641\ : Span12Mux_h
    port map (
            O => \N__8201\,
            I => \N__8198\
        );

    \I__1640\ : Odrv12
    port map (
            O => \N__8198\,
            I => \C3_c\
        );

    \I__1639\ : InMux
    port map (
            O => \N__8195\,
            I => \N__8192\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__8192\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1637\ : InMux
    port map (
            O => \N__8189\,
            I => \N__8186\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__8186\,
            I => \U712_CHIP_RAM.N_346\
        );

    \I__1635\ : InMux
    port map (
            O => \N__8183\,
            I => \N__8180\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__8180\,
            I => \U712_CHIP_RAM.N_352\
        );

    \I__1633\ : IoInMux
    port map (
            O => \N__8177\,
            I => \N__8174\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__8174\,
            I => \N__8171\
        );

    \I__1631\ : IoSpan4Mux
    port map (
            O => \N__8171\,
            I => \N__8168\
        );

    \I__1630\ : Sp12to4
    port map (
            O => \N__8168\,
            I => \N__8165\
        );

    \I__1629\ : Span12Mux_s7_h
    port map (
            O => \N__8165\,
            I => \N__8162\
        );

    \I__1628\ : Span12Mux_v
    port map (
            O => \N__8162\,
            I => \N__8159\
        );

    \I__1627\ : Odrv12
    port map (
            O => \N__8159\,
            I => \CMA_c_5\
        );

    \I__1626\ : InMux
    port map (
            O => \N__8156\,
            I => \N__8152\
        );

    \I__1625\ : InMux
    port map (
            O => \N__8155\,
            I => \N__8149\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__8152\,
            I => \N__8146\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__8149\,
            I => \N__8143\
        );

    \I__1622\ : Span4Mux_h
    port map (
            O => \N__8146\,
            I => \N__8140\
        );

    \I__1621\ : Span4Mux_v
    port map (
            O => \N__8143\,
            I => \N__8137\
        );

    \I__1620\ : Span4Mux_v
    port map (
            O => \N__8140\,
            I => \N__8134\
        );

    \I__1619\ : Span4Mux_h
    port map (
            O => \N__8137\,
            I => \N__8131\
        );

    \I__1618\ : Odrv4
    port map (
            O => \N__8134\,
            I => \DBRn_c_i\
        );

    \I__1617\ : Odrv4
    port map (
            O => \N__8131\,
            I => \DBRn_c_i\
        );

    \I__1616\ : InMux
    port map (
            O => \N__8126\,
            I => \N__8122\
        );

    \I__1615\ : InMux
    port map (
            O => \N__8125\,
            I => \N__8119\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__8122\,
            I => \N__8116\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__8119\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__1612\ : Odrv4
    port map (
            O => \N__8116\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__1611\ : IoInMux
    port map (
            O => \N__8111\,
            I => \N__8108\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__8108\,
            I => \N__8105\
        );

    \I__1609\ : Span4Mux_s0_v
    port map (
            O => \N__8105\,
            I => \N__8102\
        );

    \I__1608\ : Span4Mux_v
    port map (
            O => \N__8102\,
            I => \N__8099\
        );

    \I__1607\ : Span4Mux_v
    port map (
            O => \N__8099\,
            I => \N__8096\
        );

    \I__1606\ : Sp12to4
    port map (
            O => \N__8096\,
            I => \N__8093\
        );

    \I__1605\ : Span12Mux_h
    port map (
            O => \N__8093\,
            I => \N__8090\
        );

    \I__1604\ : Odrv12
    port map (
            O => \N__8090\,
            I => \N_169_i\
        );

    \I__1603\ : InMux
    port map (
            O => \N__8087\,
            I => \N__8084\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__8084\,
            I => \N__8081\
        );

    \I__1601\ : Span4Mux_v
    port map (
            O => \N__8081\,
            I => \N__8078\
        );

    \I__1600\ : Span4Mux_v
    port map (
            O => \N__8078\,
            I => \N__8075\
        );

    \I__1599\ : Span4Mux_v
    port map (
            O => \N__8075\,
            I => \N__8072\
        );

    \I__1598\ : Sp12to4
    port map (
            O => \N__8072\,
            I => \N__8069\
        );

    \I__1597\ : Span12Mux_h
    port map (
            O => \N__8069\,
            I => \N__8066\
        );

    \I__1596\ : Odrv12
    port map (
            O => \N__8066\,
            I => \REGSPACEn_c\
        );

    \I__1595\ : CascadeMux
    port map (
            O => \N__8063\,
            I => \U712_REG_SM.N_397_cascade_\
        );

    \I__1594\ : InMux
    port map (
            O => \N__8060\,
            I => \N__8057\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__8057\,
            I => \N__8054\
        );

    \I__1592\ : Span4Mux_v
    port map (
            O => \N__8054\,
            I => \N__8050\
        );

    \I__1591\ : InMux
    port map (
            O => \N__8053\,
            I => \N__8047\
        );

    \I__1590\ : Sp12to4
    port map (
            O => \N__8050\,
            I => \N__8044\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__8047\,
            I => \N__8041\
        );

    \I__1588\ : Span12Mux_h
    port map (
            O => \N__8044\,
            I => \N__8038\
        );

    \I__1587\ : Span12Mux_h
    port map (
            O => \N__8041\,
            I => \N__8035\
        );

    \I__1586\ : Span12Mux_v
    port map (
            O => \N__8038\,
            I => \N__8032\
        );

    \I__1585\ : Span12Mux_v
    port map (
            O => \N__8035\,
            I => \N__8029\
        );

    \I__1584\ : Odrv12
    port map (
            O => \N__8032\,
            I => \TSn_c\
        );

    \I__1583\ : Odrv12
    port map (
            O => \N__8029\,
            I => \TSn_c\
        );

    \I__1582\ : InMux
    port map (
            O => \N__8024\,
            I => \N__8021\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__8021\,
            I => \N__8018\
        );

    \I__1580\ : Odrv12
    port map (
            O => \N__8018\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_3\
        );

    \I__1579\ : InMux
    port map (
            O => \N__8015\,
            I => \N__8011\
        );

    \I__1578\ : InMux
    port map (
            O => \N__8014\,
            I => \N__8008\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__8011\,
            I => \U712_REG_SM.N_548\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__8008\,
            I => \U712_REG_SM.N_548\
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__8003\,
            I => \U712_REG_SM.N_319_cascade_\
        );

    \I__1574\ : CascadeMux
    port map (
            O => \N__8000\,
            I => \U712_REG_SM.N_320_cascade_\
        );

    \I__1573\ : IoInMux
    port map (
            O => \N__7997\,
            I => \N__7994\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__7994\,
            I => \N__7991\
        );

    \I__1571\ : Span12Mux_s1_v
    port map (
            O => \N__7991\,
            I => \N__7988\
        );

    \I__1570\ : Odrv12
    port map (
            O => \N__7988\,
            I => \RESETn_c_i\
        );

    \I__1569\ : InMux
    port map (
            O => \N__7985\,
            I => \N__7982\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__7982\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\
        );

    \I__1567\ : CascadeMux
    port map (
            O => \N__7979\,
            I => \N__7976\
        );

    \I__1566\ : InMux
    port map (
            O => \N__7976\,
            I => \N__7973\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__7973\,
            I => \N__7970\
        );

    \I__1564\ : Span4Mux_h
    port map (
            O => \N__7970\,
            I => \N__7967\
        );

    \I__1563\ : Odrv4
    port map (
            O => \N__7967\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__1562\ : InMux
    port map (
            O => \N__7964\,
            I => \N__7961\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__7961\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i\
        );

    \I__1560\ : InMux
    port map (
            O => \N__7958\,
            I => \N__7955\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__7955\,
            I => \N__7952\
        );

    \I__1558\ : Odrv4
    port map (
            O => \N__7952\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8\
        );

    \I__1557\ : InMux
    port map (
            O => \N__7949\,
            I => \N__7946\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__7946\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__7943\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_\
        );

    \I__1554\ : InMux
    port map (
            O => \N__7940\,
            I => \N__7937\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__7937\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__1552\ : IoInMux
    port map (
            O => \N__7934\,
            I => \N__7931\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__7931\,
            I => \N__7928\
        );

    \I__1550\ : Span4Mux_s3_v
    port map (
            O => \N__7928\,
            I => \N__7925\
        );

    \I__1549\ : Span4Mux_v
    port map (
            O => \N__7925\,
            I => \N__7922\
        );

    \I__1548\ : Span4Mux_v
    port map (
            O => \N__7922\,
            I => \N__7919\
        );

    \I__1547\ : Odrv4
    port map (
            O => \N__7919\,
            I => \CMA_c_1\
        );

    \I__1546\ : InMux
    port map (
            O => \N__7916\,
            I => \N__7913\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__7913\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__1544\ : InMux
    port map (
            O => \N__7910\,
            I => \N__7902\
        );

    \I__1543\ : InMux
    port map (
            O => \N__7909\,
            I => \N__7902\
        );

    \I__1542\ : InMux
    port map (
            O => \N__7908\,
            I => \N__7897\
        );

    \I__1541\ : InMux
    port map (
            O => \N__7907\,
            I => \N__7897\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__7902\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__7897\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1538\ : InMux
    port map (
            O => \N__7892\,
            I => \N__7889\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__7889\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\
        );

    \I__1536\ : CascadeMux
    port map (
            O => \N__7886\,
            I => \N__7883\
        );

    \I__1535\ : InMux
    port map (
            O => \N__7883\,
            I => \N__7880\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__7880\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1533\ : InMux
    port map (
            O => \N__7877\,
            I => \N__7873\
        );

    \I__1532\ : InMux
    port map (
            O => \N__7876\,
            I => \N__7870\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__7873\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__7870\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1529\ : CascadeMux
    port map (
            O => \N__7865\,
            I => \N__7861\
        );

    \I__1528\ : InMux
    port map (
            O => \N__7864\,
            I => \N__7855\
        );

    \I__1527\ : InMux
    port map (
            O => \N__7861\,
            I => \N__7855\
        );

    \I__1526\ : InMux
    port map (
            O => \N__7860\,
            I => \N__7852\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__7855\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__7852\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1523\ : InMux
    port map (
            O => \N__7847\,
            I => \N__7841\
        );

    \I__1522\ : InMux
    port map (
            O => \N__7846\,
            I => \N__7836\
        );

    \I__1521\ : InMux
    port map (
            O => \N__7845\,
            I => \N__7836\
        );

    \I__1520\ : InMux
    port map (
            O => \N__7844\,
            I => \N__7833\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__7841\,
            I => \REG_TACK\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__7836\,
            I => \REG_TACK\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__7833\,
            I => \REG_TACK\
        );

    \I__1516\ : InMux
    port map (
            O => \N__7826\,
            I => \N__7823\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__7823\,
            I => \U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7820\,
            I => \N__7814\
        );

    \I__1513\ : InMux
    port map (
            O => \N__7819\,
            I => \N__7814\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__7814\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_5\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7811\,
            I => \N__7808\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__7808\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_6\
        );

    \I__1509\ : InMux
    port map (
            O => \N__7805\,
            I => \N__7802\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__7802\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_4\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7799\,
            I => \N__7795\
        );

    \I__1506\ : InMux
    port map (
            O => \N__7798\,
            I => \N__7792\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__7795\,
            I => \N__7789\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__7792\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0Z0Z_0\
        );

    \I__1503\ : Odrv12
    port map (
            O => \N__7789\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0Z0Z_0\
        );

    \I__1502\ : CascadeMux
    port map (
            O => \N__7784\,
            I => \N__7781\
        );

    \I__1501\ : InMux
    port map (
            O => \N__7781\,
            I => \N__7778\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__7778\,
            I => \N__7775\
        );

    \I__1499\ : Span4Mux_v
    port map (
            O => \N__7775\,
            I => \N__7772\
        );

    \I__1498\ : Odrv4
    port map (
            O => \N__7772\,
            I => \U712_BYTE_ENABLE.N_325\
        );

    \I__1497\ : IoInMux
    port map (
            O => \N__7769\,
            I => \N__7766\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__7766\,
            I => \N__7763\
        );

    \I__1495\ : Span12Mux_s10_h
    port map (
            O => \N__7763\,
            I => \N__7760\
        );

    \I__1494\ : Span12Mux_v
    port map (
            O => \N__7760\,
            I => \N__7757\
        );

    \I__1493\ : Odrv12
    port map (
            O => \N__7757\,
            I => \N_186_i\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7754\,
            I => \N__7748\
        );

    \I__1491\ : InMux
    port map (
            O => \N__7753\,
            I => \N__7745\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7752\,
            I => \N__7740\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7751\,
            I => \N__7740\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__7748\,
            I => \CPU_TACKm\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__7745\,
            I => \CPU_TACKm\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__7740\,
            I => \CPU_TACKm\
        );

    \I__1485\ : CascadeMux
    port map (
            O => \N__7733\,
            I => \U712_CYCLE_TERM.N_450_cascade_\
        );

    \I__1484\ : CascadeMux
    port map (
            O => \N__7730\,
            I => \N__7727\
        );

    \I__1483\ : InMux
    port map (
            O => \N__7727\,
            I => \N__7721\
        );

    \I__1482\ : InMux
    port map (
            O => \N__7726\,
            I => \N__7721\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__7721\,
            I => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7718\,
            I => \N__7715\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__7715\,
            I => \N__7711\
        );

    \I__1478\ : CascadeMux
    port map (
            O => \N__7714\,
            I => \N__7706\
        );

    \I__1477\ : Span4Mux_v
    port map (
            O => \N__7711\,
            I => \N__7703\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7710\,
            I => \N__7698\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7709\,
            I => \N__7698\
        );

    \I__1474\ : InMux
    port map (
            O => \N__7706\,
            I => \N__7695\
        );

    \I__1473\ : Span4Mux_v
    port map (
            O => \N__7703\,
            I => \N__7692\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__7698\,
            I => \N__7689\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__7695\,
            I => \N__7686\
        );

    \I__1470\ : Sp12to4
    port map (
            O => \N__7692\,
            I => \N__7683\
        );

    \I__1469\ : Sp12to4
    port map (
            O => \N__7689\,
            I => \N__7678\
        );

    \I__1468\ : Sp12to4
    port map (
            O => \N__7686\,
            I => \N__7678\
        );

    \I__1467\ : Span12Mux_h
    port map (
            O => \N__7683\,
            I => \N__7673\
        );

    \I__1466\ : Span12Mux_v
    port map (
            O => \N__7678\,
            I => \N__7673\
        );

    \I__1465\ : Odrv12
    port map (
            O => \N__7673\,
            I => \CLK40_PLL_i\
        );

    \I__1464\ : CascadeMux
    port map (
            O => \N__7670\,
            I => \N__7666\
        );

    \I__1463\ : InMux
    port map (
            O => \N__7669\,
            I => \N__7662\
        );

    \I__1462\ : InMux
    port map (
            O => \N__7666\,
            I => \N__7657\
        );

    \I__1461\ : InMux
    port map (
            O => \N__7665\,
            I => \N__7657\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__7662\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__7657\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1458\ : IoInMux
    port map (
            O => \N__7652\,
            I => \N__7648\
        );

    \I__1457\ : IoInMux
    port map (
            O => \N__7651\,
            I => \N__7644\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__7648\,
            I => \N__7641\
        );

    \I__1455\ : IoInMux
    port map (
            O => \N__7647\,
            I => \N__7638\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__7644\,
            I => \N__7635\
        );

    \I__1453\ : IoSpan4Mux
    port map (
            O => \N__7641\,
            I => \N__7632\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__7638\,
            I => \N__7629\
        );

    \I__1451\ : Span4Mux_s3_v
    port map (
            O => \N__7635\,
            I => \N__7626\
        );

    \I__1450\ : Span4Mux_s3_h
    port map (
            O => \N__7632\,
            I => \N__7623\
        );

    \I__1449\ : Span4Mux_s0_v
    port map (
            O => \N__7629\,
            I => \N__7620\
        );

    \I__1448\ : Sp12to4
    port map (
            O => \N__7626\,
            I => \N__7617\
        );

    \I__1447\ : Sp12to4
    port map (
            O => \N__7623\,
            I => \N__7614\
        );

    \I__1446\ : Sp12to4
    port map (
            O => \N__7620\,
            I => \N__7611\
        );

    \I__1445\ : Span12Mux_s9_h
    port map (
            O => \N__7617\,
            I => \N__7608\
        );

    \I__1444\ : Span12Mux_v
    port map (
            O => \N__7614\,
            I => \N__7605\
        );

    \I__1443\ : Span12Mux_h
    port map (
            O => \N__7611\,
            I => \N__7602\
        );

    \I__1442\ : Span12Mux_v
    port map (
            O => \N__7608\,
            I => \N__7598\
        );

    \I__1441\ : Span12Mux_h
    port map (
            O => \N__7605\,
            I => \N__7593\
        );

    \I__1440\ : Span12Mux_v
    port map (
            O => \N__7602\,
            I => \N__7593\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7601\,
            I => \N__7590\
        );

    \I__1438\ : Odrv12
    port map (
            O => \N__7598\,
            I => \TACK_OUTn\
        );

    \I__1437\ : Odrv12
    port map (
            O => \N__7593\,
            I => \TACK_OUTn\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__7590\,
            I => \TACK_OUTn\
        );

    \I__1435\ : InMux
    port map (
            O => \N__7583\,
            I => \N__7580\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__7580\,
            I => \N__7577\
        );

    \I__1433\ : Span12Mux_v
    port map (
            O => \N__7577\,
            I => \N__7574\
        );

    \I__1432\ : Span12Mux_h
    port map (
            O => \N__7574\,
            I => \N__7571\
        );

    \I__1431\ : Odrv12
    port map (
            O => \N__7571\,
            I => \A_c_15\
        );

    \I__1430\ : InMux
    port map (
            O => \N__7568\,
            I => \N__7565\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__7565\,
            I => \N__7562\
        );

    \I__1428\ : Span4Mux_h
    port map (
            O => \N__7562\,
            I => \N__7559\
        );

    \I__1427\ : Span4Mux_h
    port map (
            O => \N__7559\,
            I => \N__7556\
        );

    \I__1426\ : Odrv4
    port map (
            O => \N__7556\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\
        );

    \I__1425\ : SRMux
    port map (
            O => \N__7553\,
            I => \N__7550\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__7550\,
            I => \N__7547\
        );

    \I__1423\ : Span4Mux_h
    port map (
            O => \N__7547\,
            I => \N__7543\
        );

    \I__1422\ : InMux
    port map (
            O => \N__7546\,
            I => \N__7540\
        );

    \I__1421\ : Span4Mux_h
    port map (
            O => \N__7543\,
            I => \N__7537\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__7540\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__1419\ : Odrv4
    port map (
            O => \N__7537\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__1418\ : IoInMux
    port map (
            O => \N__7532\,
            I => \N__7529\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__7529\,
            I => \N__7525\
        );

    \I__1416\ : InMux
    port map (
            O => \N__7528\,
            I => \N__7522\
        );

    \I__1415\ : Span12Mux_s4_v
    port map (
            O => \N__7525\,
            I => \N__7519\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__7522\,
            I => \N__7516\
        );

    \I__1413\ : Span12Mux_v
    port map (
            O => \N__7519\,
            I => \N__7511\
        );

    \I__1412\ : Span12Mux_v
    port map (
            O => \N__7516\,
            I => \N__7511\
        );

    \I__1411\ : Span12Mux_h
    port map (
            O => \N__7511\,
            I => \N__7508\
        );

    \I__1410\ : Odrv12
    port map (
            O => \N__7508\,
            I => \A_c_9\
        );

    \I__1409\ : InMux
    port map (
            O => \N__7505\,
            I => \N__7502\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__7502\,
            I => \N__7499\
        );

    \I__1407\ : Odrv12
    port map (
            O => \N__7499\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\
        );

    \I__1406\ : CascadeMux
    port map (
            O => \N__7496\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\
        );

    \I__1405\ : IoInMux
    port map (
            O => \N__7493\,
            I => \N__7490\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__7490\,
            I => \N__7487\
        );

    \I__1403\ : IoSpan4Mux
    port map (
            O => \N__7487\,
            I => \N__7484\
        );

    \I__1402\ : IoSpan4Mux
    port map (
            O => \N__7484\,
            I => \N__7481\
        );

    \I__1401\ : IoSpan4Mux
    port map (
            O => \N__7481\,
            I => \N__7478\
        );

    \I__1400\ : Span4Mux_s2_v
    port map (
            O => \N__7478\,
            I => \N__7475\
        );

    \I__1399\ : Sp12to4
    port map (
            O => \N__7475\,
            I => \N__7471\
        );

    \I__1398\ : InMux
    port map (
            O => \N__7474\,
            I => \N__7468\
        );

    \I__1397\ : Span12Mux_s8_v
    port map (
            O => \N__7471\,
            I => \N__7465\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__7468\,
            I => \N__7462\
        );

    \I__1395\ : Span12Mux_v
    port map (
            O => \N__7465\,
            I => \N__7457\
        );

    \I__1394\ : Span12Mux_h
    port map (
            O => \N__7462\,
            I => \N__7457\
        );

    \I__1393\ : Odrv12
    port map (
            O => \N__7457\,
            I => \A_c_10\
        );

    \I__1392\ : InMux
    port map (
            O => \N__7454\,
            I => \N__7451\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__7451\,
            I => \N__7448\
        );

    \I__1390\ : Odrv12
    port map (
            O => \N__7448\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__7445\,
            I => \U712_CHIP_RAM.N_305_cascade_\
        );

    \I__1388\ : InMux
    port map (
            O => \N__7442\,
            I => \N__7439\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__7439\,
            I => \N__7436\
        );

    \I__1386\ : Span4Mux_v
    port map (
            O => \N__7436\,
            I => \N__7433\
        );

    \I__1385\ : Span4Mux_v
    port map (
            O => \N__7433\,
            I => \N__7430\
        );

    \I__1384\ : Sp12to4
    port map (
            O => \N__7430\,
            I => \N__7427\
        );

    \I__1383\ : Span12Mux_h
    port map (
            O => \N__7427\,
            I => \N__7424\
        );

    \I__1382\ : Odrv12
    port map (
            O => \N__7424\,
            I => \A_c_14\
        );

    \I__1381\ : InMux
    port map (
            O => \N__7421\,
            I => \N__7418\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__7418\,
            I => \N__7415\
        );

    \I__1379\ : Span12Mux_v
    port map (
            O => \N__7415\,
            I => \N__7412\
        );

    \I__1378\ : Odrv12
    port map (
            O => \N__7412\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\
        );

    \I__1377\ : InMux
    port map (
            O => \N__7409\,
            I => \N__7401\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7408\,
            I => \N__7401\
        );

    \I__1375\ : InMux
    port map (
            O => \N__7407\,
            I => \N__7398\
        );

    \I__1374\ : InMux
    port map (
            O => \N__7406\,
            I => \N__7395\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__7401\,
            I => \U712_CHIP_RAM.N_469\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__7398\,
            I => \U712_CHIP_RAM.N_469\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__7395\,
            I => \U712_CHIP_RAM.N_469\
        );

    \I__1370\ : CascadeMux
    port map (
            O => \N__7388\,
            I => \U712_CHIP_RAM.N_438_cascade_\
        );

    \I__1369\ : InMux
    port map (
            O => \N__7385\,
            I => \N__7382\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__7382\,
            I => \N__7379\
        );

    \I__1367\ : Odrv4
    port map (
            O => \N__7379\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__7376\,
            I => \N__7370\
        );

    \I__1365\ : CascadeMux
    port map (
            O => \N__7375\,
            I => \N__7364\
        );

    \I__1364\ : InMux
    port map (
            O => \N__7374\,
            I => \N__7359\
        );

    \I__1363\ : InMux
    port map (
            O => \N__7373\,
            I => \N__7356\
        );

    \I__1362\ : InMux
    port map (
            O => \N__7370\,
            I => \N__7353\
        );

    \I__1361\ : InMux
    port map (
            O => \N__7369\,
            I => \N__7350\
        );

    \I__1360\ : InMux
    port map (
            O => \N__7368\,
            I => \N__7347\
        );

    \I__1359\ : InMux
    port map (
            O => \N__7367\,
            I => \N__7344\
        );

    \I__1358\ : InMux
    port map (
            O => \N__7364\,
            I => \N__7339\
        );

    \I__1357\ : InMux
    port map (
            O => \N__7363\,
            I => \N__7339\
        );

    \I__1356\ : CascadeMux
    port map (
            O => \N__7362\,
            I => \N__7335\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__7359\,
            I => \N__7331\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__7356\,
            I => \N__7328\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__7353\,
            I => \N__7321\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__7350\,
            I => \N__7321\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__7347\,
            I => \N__7321\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__7344\,
            I => \N__7311\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__7339\,
            I => \N__7311\
        );

    \I__1348\ : InMux
    port map (
            O => \N__7338\,
            I => \N__7308\
        );

    \I__1347\ : InMux
    port map (
            O => \N__7335\,
            I => \N__7305\
        );

    \I__1346\ : InMux
    port map (
            O => \N__7334\,
            I => \N__7302\
        );

    \I__1345\ : Span4Mux_h
    port map (
            O => \N__7331\,
            I => \N__7297\
        );

    \I__1344\ : Span4Mux_h
    port map (
            O => \N__7328\,
            I => \N__7297\
        );

    \I__1343\ : Span4Mux_h
    port map (
            O => \N__7321\,
            I => \N__7291\
        );

    \I__1342\ : InMux
    port map (
            O => \N__7320\,
            I => \N__7288\
        );

    \I__1341\ : InMux
    port map (
            O => \N__7319\,
            I => \N__7281\
        );

    \I__1340\ : InMux
    port map (
            O => \N__7318\,
            I => \N__7281\
        );

    \I__1339\ : InMux
    port map (
            O => \N__7317\,
            I => \N__7281\
        );

    \I__1338\ : InMux
    port map (
            O => \N__7316\,
            I => \N__7278\
        );

    \I__1337\ : Span4Mux_h
    port map (
            O => \N__7311\,
            I => \N__7275\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__7308\,
            I => \N__7268\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__7305\,
            I => \N__7268\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__7302\,
            I => \N__7268\
        );

    \I__1333\ : Sp12to4
    port map (
            O => \N__7297\,
            I => \N__7265\
        );

    \I__1332\ : InMux
    port map (
            O => \N__7296\,
            I => \N__7258\
        );

    \I__1331\ : InMux
    port map (
            O => \N__7295\,
            I => \N__7258\
        );

    \I__1330\ : InMux
    port map (
            O => \N__7294\,
            I => \N__7258\
        );

    \I__1329\ : Odrv4
    port map (
            O => \N__7291\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__7288\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__7281\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__7278\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1325\ : Odrv4
    port map (
            O => \N__7275\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1324\ : Odrv4
    port map (
            O => \N__7268\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1323\ : Odrv12
    port map (
            O => \N__7265\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__7258\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1321\ : CascadeMux
    port map (
            O => \N__7241\,
            I => \N__7237\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__7240\,
            I => \N__7233\
        );

    \I__1319\ : InMux
    port map (
            O => \N__7237\,
            I => \N__7230\
        );

    \I__1318\ : InMux
    port map (
            O => \N__7236\,
            I => \N__7227\
        );

    \I__1317\ : InMux
    port map (
            O => \N__7233\,
            I => \N__7223\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__7230\,
            I => \N__7218\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__7227\,
            I => \N__7215\
        );

    \I__1314\ : InMux
    port map (
            O => \N__7226\,
            I => \N__7208\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__7223\,
            I => \N__7205\
        );

    \I__1312\ : CascadeMux
    port map (
            O => \N__7222\,
            I => \N__7202\
        );

    \I__1311\ : InMux
    port map (
            O => \N__7221\,
            I => \N__7198\
        );

    \I__1310\ : Span4Mux_v
    port map (
            O => \N__7218\,
            I => \N__7195\
        );

    \I__1309\ : Span4Mux_h
    port map (
            O => \N__7215\,
            I => \N__7192\
        );

    \I__1308\ : InMux
    port map (
            O => \N__7214\,
            I => \N__7189\
        );

    \I__1307\ : InMux
    port map (
            O => \N__7213\,
            I => \N__7186\
        );

    \I__1306\ : InMux
    port map (
            O => \N__7212\,
            I => \N__7181\
        );

    \I__1305\ : InMux
    port map (
            O => \N__7211\,
            I => \N__7181\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__7208\,
            I => \N__7178\
        );

    \I__1303\ : Span4Mux_v
    port map (
            O => \N__7205\,
            I => \N__7175\
        );

    \I__1302\ : InMux
    port map (
            O => \N__7202\,
            I => \N__7172\
        );

    \I__1301\ : InMux
    port map (
            O => \N__7201\,
            I => \N__7169\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__7198\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1299\ : Odrv4
    port map (
            O => \N__7195\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1298\ : Odrv4
    port map (
            O => \N__7192\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__7189\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__7186\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__7181\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1294\ : Odrv4
    port map (
            O => \N__7178\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1293\ : Odrv4
    port map (
            O => \N__7175\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__7172\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__7169\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1290\ : InMux
    port map (
            O => \N__7148\,
            I => \N__7141\
        );

    \I__1289\ : CascadeMux
    port map (
            O => \N__7147\,
            I => \N__7136\
        );

    \I__1288\ : InMux
    port map (
            O => \N__7146\,
            I => \N__7133\
        );

    \I__1287\ : CascadeMux
    port map (
            O => \N__7145\,
            I => \N__7128\
        );

    \I__1286\ : InMux
    port map (
            O => \N__7144\,
            I => \N__7125\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__7141\,
            I => \N__7122\
        );

    \I__1284\ : InMux
    port map (
            O => \N__7140\,
            I => \N__7119\
        );

    \I__1283\ : InMux
    port map (
            O => \N__7139\,
            I => \N__7116\
        );

    \I__1282\ : InMux
    port map (
            O => \N__7136\,
            I => \N__7113\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__7133\,
            I => \N__7106\
        );

    \I__1280\ : InMux
    port map (
            O => \N__7132\,
            I => \N__7103\
        );

    \I__1279\ : InMux
    port map (
            O => \N__7131\,
            I => \N__7098\
        );

    \I__1278\ : InMux
    port map (
            O => \N__7128\,
            I => \N__7098\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__7125\,
            I => \N__7087\
        );

    \I__1276\ : Span4Mux_v
    port map (
            O => \N__7122\,
            I => \N__7087\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__7119\,
            I => \N__7087\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__7116\,
            I => \N__7087\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__7113\,
            I => \N__7087\
        );

    \I__1272\ : InMux
    port map (
            O => \N__7112\,
            I => \N__7080\
        );

    \I__1271\ : InMux
    port map (
            O => \N__7111\,
            I => \N__7080\
        );

    \I__1270\ : InMux
    port map (
            O => \N__7110\,
            I => \N__7080\
        );

    \I__1269\ : InMux
    port map (
            O => \N__7109\,
            I => \N__7077\
        );

    \I__1268\ : Odrv4
    port map (
            O => \N__7106\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__7103\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__7098\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1265\ : Odrv4
    port map (
            O => \N__7087\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__7080\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__7077\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1262\ : InMux
    port map (
            O => \N__7064\,
            I => \N__7061\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__7061\,
            I => \N__7058\
        );

    \I__1260\ : Span4Mux_h
    port map (
            O => \N__7058\,
            I => \N__7055\
        );

    \I__1259\ : Odrv4
    port map (
            O => \N__7055\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_a2_1\
        );

    \I__1258\ : CascadeMux
    port map (
            O => \N__7052\,
            I => \N__7048\
        );

    \I__1257\ : InMux
    port map (
            O => \N__7051\,
            I => \N__7043\
        );

    \I__1256\ : InMux
    port map (
            O => \N__7048\,
            I => \N__7043\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__7043\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_a2_2\
        );

    \I__1254\ : IoInMux
    port map (
            O => \N__7040\,
            I => \N__7037\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__7037\,
            I => \N__7034\
        );

    \I__1252\ : Span4Mux_s3_v
    port map (
            O => \N__7034\,
            I => \N__7031\
        );

    \I__1251\ : Sp12to4
    port map (
            O => \N__7031\,
            I => \N__7027\
        );

    \I__1250\ : InMux
    port map (
            O => \N__7030\,
            I => \N__7024\
        );

    \I__1249\ : Span12Mux_h
    port map (
            O => \N__7027\,
            I => \N__7019\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__7024\,
            I => \N__7016\
        );

    \I__1247\ : InMux
    port map (
            O => \N__7023\,
            I => \N__7013\
        );

    \I__1246\ : InMux
    port map (
            O => \N__7022\,
            I => \N__7010\
        );

    \I__1245\ : Odrv12
    port map (
            O => \N__7019\,
            I => \DBENn_c\
        );

    \I__1244\ : Odrv4
    port map (
            O => \N__7016\,
            I => \DBENn_c\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__7013\,
            I => \DBENn_c\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__7010\,
            I => \DBENn_c\
        );

    \I__1241\ : CascadeMux
    port map (
            O => \N__7001\,
            I => \N__6998\
        );

    \I__1240\ : InMux
    port map (
            O => \N__6998\,
            I => \N__6991\
        );

    \I__1239\ : InMux
    port map (
            O => \N__6997\,
            I => \N__6988\
        );

    \I__1238\ : InMux
    port map (
            O => \N__6996\,
            I => \N__6985\
        );

    \I__1237\ : InMux
    port map (
            O => \N__6995\,
            I => \N__6982\
        );

    \I__1236\ : InMux
    port map (
            O => \N__6994\,
            I => \N__6979\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__6991\,
            I => \N__6974\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__6988\,
            I => \N__6971\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__6985\,
            I => \N__6968\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__6982\,
            I => \N__6965\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__6979\,
            I => \N__6962\
        );

    \I__1230\ : InMux
    port map (
            O => \N__6978\,
            I => \N__6959\
        );

    \I__1229\ : InMux
    port map (
            O => \N__6977\,
            I => \N__6956\
        );

    \I__1228\ : Span4Mux_v
    port map (
            O => \N__6974\,
            I => \N__6949\
        );

    \I__1227\ : Span4Mux_h
    port map (
            O => \N__6971\,
            I => \N__6949\
        );

    \I__1226\ : Span4Mux_v
    port map (
            O => \N__6968\,
            I => \N__6949\
        );

    \I__1225\ : Span4Mux_v
    port map (
            O => \N__6965\,
            I => \N__6942\
        );

    \I__1224\ : Span4Mux_v
    port map (
            O => \N__6962\,
            I => \N__6942\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__6959\,
            I => \N__6942\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__6956\,
            I => \DMA_CYCLEm\
        );

    \I__1221\ : Odrv4
    port map (
            O => \N__6949\,
            I => \DMA_CYCLEm\
        );

    \I__1220\ : Odrv4
    port map (
            O => \N__6942\,
            I => \DMA_CYCLEm\
        );

    \I__1219\ : InMux
    port map (
            O => \N__6935\,
            I => \N__6932\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__6932\,
            I => \U712_CYCLE_TERM.N_321\
        );

    \I__1217\ : IoInMux
    port map (
            O => \N__6929\,
            I => \N__6925\
        );

    \I__1216\ : IoInMux
    port map (
            O => \N__6928\,
            I => \N__6922\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__6925\,
            I => \N__6918\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__6922\,
            I => \N__6915\
        );

    \I__1213\ : IoInMux
    port map (
            O => \N__6921\,
            I => \N__6912\
        );

    \I__1212\ : IoSpan4Mux
    port map (
            O => \N__6918\,
            I => \N__6909\
        );

    \I__1211\ : IoSpan4Mux
    port map (
            O => \N__6915\,
            I => \N__6906\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__6912\,
            I => \N__6903\
        );

    \I__1209\ : Span4Mux_s1_h
    port map (
            O => \N__6909\,
            I => \N__6900\
        );

    \I__1208\ : Sp12to4
    port map (
            O => \N__6906\,
            I => \N__6897\
        );

    \I__1207\ : Span4Mux_s3_v
    port map (
            O => \N__6903\,
            I => \N__6894\
        );

    \I__1206\ : Sp12to4
    port map (
            O => \N__6900\,
            I => \N__6891\
        );

    \I__1205\ : Span12Mux_s3_v
    port map (
            O => \N__6897\,
            I => \N__6888\
        );

    \I__1204\ : Sp12to4
    port map (
            O => \N__6894\,
            I => \N__6885\
        );

    \I__1203\ : Span12Mux_h
    port map (
            O => \N__6891\,
            I => \N__6881\
        );

    \I__1202\ : Span12Mux_h
    port map (
            O => \N__6888\,
            I => \N__6876\
        );

    \I__1201\ : Span12Mux_h
    port map (
            O => \N__6885\,
            I => \N__6876\
        );

    \I__1200\ : InMux
    port map (
            O => \N__6884\,
            I => \N__6873\
        );

    \I__1199\ : Odrv12
    port map (
            O => \N__6881\,
            I => \TACK_EN\
        );

    \I__1198\ : Odrv12
    port map (
            O => \N__6876\,
            I => \TACK_EN\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__6873\,
            I => \TACK_EN\
        );

    \I__1196\ : InMux
    port map (
            O => \N__6866\,
            I => \N__6863\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__6863\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__1194\ : IoInMux
    port map (
            O => \N__6860\,
            I => \N__6857\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__6857\,
            I => \N__6854\
        );

    \I__1192\ : IoSpan4Mux
    port map (
            O => \N__6854\,
            I => \N__6851\
        );

    \I__1191\ : Sp12to4
    port map (
            O => \N__6851\,
            I => \N__6848\
        );

    \I__1190\ : Odrv12
    port map (
            O => \N__6848\,
            I => \CMA_c_2\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6845\,
            I => \N__6842\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__6842\,
            I => \N__6839\
        );

    \I__1187\ : Span12Mux_h
    port map (
            O => \N__6839\,
            I => \N__6836\
        );

    \I__1186\ : Odrv12
    port map (
            O => \N__6836\,
            I => \A_c_13\
        );

    \I__1185\ : InMux
    port map (
            O => \N__6833\,
            I => \N__6830\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__6830\,
            I => \N__6827\
        );

    \I__1183\ : Odrv12
    port map (
            O => \N__6827\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\
        );

    \I__1182\ : CascadeMux
    port map (
            O => \N__6824\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\
        );

    \I__1181\ : InMux
    port map (
            O => \N__6821\,
            I => \N__6813\
        );

    \I__1180\ : InMux
    port map (
            O => \N__6820\,
            I => \N__6813\
        );

    \I__1179\ : InMux
    port map (
            O => \N__6819\,
            I => \N__6810\
        );

    \I__1178\ : InMux
    port map (
            O => \N__6818\,
            I => \N__6807\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__6813\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__6810\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6807\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__1174\ : CascadeMux
    port map (
            O => \N__6800\,
            I => \U712_CHIP_RAM.N_442_cascade_\
        );

    \I__1173\ : InMux
    port map (
            O => \N__6797\,
            I => \N__6791\
        );

    \I__1172\ : InMux
    port map (
            O => \N__6796\,
            I => \N__6791\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__6791\,
            I => \U712_CHIP_RAM.N_441\
        );

    \I__1170\ : InMux
    port map (
            O => \N__6788\,
            I => \N__6785\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__6785\,
            I => \N__6782\
        );

    \I__1168\ : Span4Mux_h
    port map (
            O => \N__6782\,
            I => \N__6779\
        );

    \I__1167\ : Odrv4
    port map (
            O => \N__6779\,
            I => \U712_CHIP_RAM.CPU_TACK_8_iv_i_a2_1\
        );

    \I__1166\ : CascadeMux
    port map (
            O => \N__6776\,
            I => \N__6772\
        );

    \I__1165\ : CascadeMux
    port map (
            O => \N__6775\,
            I => \N__6769\
        );

    \I__1164\ : InMux
    port map (
            O => \N__6772\,
            I => \N__6762\
        );

    \I__1163\ : InMux
    port map (
            O => \N__6769\,
            I => \N__6762\
        );

    \I__1162\ : InMux
    port map (
            O => \N__6768\,
            I => \N__6756\
        );

    \I__1161\ : InMux
    port map (
            O => \N__6767\,
            I => \N__6753\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__6762\,
            I => \N__6750\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6761\,
            I => \N__6745\
        );

    \I__1158\ : InMux
    port map (
            O => \N__6760\,
            I => \N__6745\
        );

    \I__1157\ : InMux
    port map (
            O => \N__6759\,
            I => \N__6742\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__6756\,
            I => \U712_CHIP_RAM.N_295\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__6753\,
            I => \U712_CHIP_RAM.N_295\
        );

    \I__1154\ : Odrv4
    port map (
            O => \N__6750\,
            I => \U712_CHIP_RAM.N_295\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__6745\,
            I => \U712_CHIP_RAM.N_295\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__6742\,
            I => \U712_CHIP_RAM.N_295\
        );

    \I__1151\ : InMux
    port map (
            O => \N__6731\,
            I => \N__6728\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__6728\,
            I => \N__6724\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6727\,
            I => \N__6720\
        );

    \I__1148\ : Span4Mux_v
    port map (
            O => \N__6724\,
            I => \N__6717\
        );

    \I__1147\ : InMux
    port map (
            O => \N__6723\,
            I => \N__6714\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__6720\,
            I => \N__6707\
        );

    \I__1145\ : Sp12to4
    port map (
            O => \N__6717\,
            I => \N__6707\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__6714\,
            I => \N__6707\
        );

    \I__1143\ : Span12Mux_h
    port map (
            O => \N__6707\,
            I => \N__6704\
        );

    \I__1142\ : Span12Mux_v
    port map (
            O => \N__6704\,
            I => \N__6701\
        );

    \I__1141\ : Odrv12
    port map (
            O => \N__6701\,
            I => \AWEn_c\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6698\,
            I => \N__6693\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6697\,
            I => \N__6690\
        );

    \I__1138\ : InMux
    port map (
            O => \N__6696\,
            I => \N__6687\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__6693\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__6690\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__6687\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\
        );

    \I__1134\ : InMux
    port map (
            O => \N__6680\,
            I => \N__6677\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__6677\,
            I => \N__6672\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6676\,
            I => \N__6669\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6675\,
            I => \N__6666\
        );

    \I__1130\ : Odrv4
    port map (
            O => \N__6672\,
            I => \U712_CHIP_RAM.N_551\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6669\,
            I => \U712_CHIP_RAM.N_551\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__6666\,
            I => \U712_CHIP_RAM.N_551\
        );

    \I__1127\ : CascadeMux
    port map (
            O => \N__6659\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_cascade_\
        );

    \I__1126\ : CEMux
    port map (
            O => \N__6656\,
            I => \N__6653\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__6653\,
            I => \N__6650\
        );

    \I__1124\ : Span4Mux_v
    port map (
            O => \N__6650\,
            I => \N__6647\
        );

    \I__1123\ : Odrv4
    port map (
            O => \N__6647\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0\
        );

    \I__1122\ : InMux
    port map (
            O => \N__6644\,
            I => \N__6639\
        );

    \I__1121\ : CascadeMux
    port map (
            O => \N__6643\,
            I => \N__6636\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6642\,
            I => \N__6630\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__6639\,
            I => \N__6627\
        );

    \I__1118\ : InMux
    port map (
            O => \N__6636\,
            I => \N__6624\
        );

    \I__1117\ : InMux
    port map (
            O => \N__6635\,
            I => \N__6617\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6634\,
            I => \N__6617\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6633\,
            I => \N__6614\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__6630\,
            I => \N__6607\
        );

    \I__1113\ : Span4Mux_v
    port map (
            O => \N__6627\,
            I => \N__6607\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__6624\,
            I => \N__6607\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6623\,
            I => \N__6602\
        );

    \I__1110\ : InMux
    port map (
            O => \N__6622\,
            I => \N__6602\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__6617\,
            I => \U712_CHIP_RAM.N_458\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__6614\,
            I => \U712_CHIP_RAM.N_458\
        );

    \I__1107\ : Odrv4
    port map (
            O => \N__6607\,
            I => \U712_CHIP_RAM.N_458\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__6602\,
            I => \U712_CHIP_RAM.N_458\
        );

    \I__1105\ : InMux
    port map (
            O => \N__6593\,
            I => \N__6590\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__6590\,
            I => \N__6587\
        );

    \I__1103\ : Span4Mux_h
    port map (
            O => \N__6587\,
            I => \N__6584\
        );

    \I__1102\ : Odrv4
    port map (
            O => \N__6584\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_0_0_0_a2_1\
        );

    \I__1101\ : InMux
    port map (
            O => \N__6581\,
            I => \N__6578\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__6578\,
            I => \N__6575\
        );

    \I__1099\ : Odrv4
    port map (
            O => \N__6575\,
            I => \U712_CHIP_RAM.N_428\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__6572\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_0_cascade_\
        );

    \I__1097\ : CascadeMux
    port map (
            O => \N__6569\,
            I => \N__6566\
        );

    \I__1096\ : InMux
    port map (
            O => \N__6566\,
            I => \N__6563\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__6563\,
            I => \N__6559\
        );

    \I__1094\ : InMux
    port map (
            O => \N__6562\,
            I => \N__6556\
        );

    \I__1093\ : Span4Mux_v
    port map (
            O => \N__6559\,
            I => \N__6551\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__6556\,
            I => \N__6551\
        );

    \I__1091\ : Odrv4
    port map (
            O => \N__6551\,
            I => \U712_CHIP_RAM.N_300\
        );

    \I__1090\ : CascadeMux
    port map (
            O => \N__6548\,
            I => \N__6543\
        );

    \I__1089\ : CascadeMux
    port map (
            O => \N__6547\,
            I => \N__6528\
        );

    \I__1088\ : InMux
    port map (
            O => \N__6546\,
            I => \N__6520\
        );

    \I__1087\ : InMux
    port map (
            O => \N__6543\,
            I => \N__6512\
        );

    \I__1086\ : CascadeMux
    port map (
            O => \N__6542\,
            I => \N__6509\
        );

    \I__1085\ : InMux
    port map (
            O => \N__6541\,
            I => \N__6506\
        );

    \I__1084\ : InMux
    port map (
            O => \N__6540\,
            I => \N__6503\
        );

    \I__1083\ : InMux
    port map (
            O => \N__6539\,
            I => \N__6498\
        );

    \I__1082\ : InMux
    port map (
            O => \N__6538\,
            I => \N__6498\
        );

    \I__1081\ : InMux
    port map (
            O => \N__6537\,
            I => \N__6495\
        );

    \I__1080\ : InMux
    port map (
            O => \N__6536\,
            I => \N__6488\
        );

    \I__1079\ : InMux
    port map (
            O => \N__6535\,
            I => \N__6488\
        );

    \I__1078\ : InMux
    port map (
            O => \N__6534\,
            I => \N__6488\
        );

    \I__1077\ : InMux
    port map (
            O => \N__6533\,
            I => \N__6479\
        );

    \I__1076\ : InMux
    port map (
            O => \N__6532\,
            I => \N__6479\
        );

    \I__1075\ : InMux
    port map (
            O => \N__6531\,
            I => \N__6479\
        );

    \I__1074\ : InMux
    port map (
            O => \N__6528\,
            I => \N__6479\
        );

    \I__1073\ : InMux
    port map (
            O => \N__6527\,
            I => \N__6471\
        );

    \I__1072\ : InMux
    port map (
            O => \N__6526\,
            I => \N__6471\
        );

    \I__1071\ : InMux
    port map (
            O => \N__6525\,
            I => \N__6464\
        );

    \I__1070\ : InMux
    port map (
            O => \N__6524\,
            I => \N__6464\
        );

    \I__1069\ : InMux
    port map (
            O => \N__6523\,
            I => \N__6464\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__6520\,
            I => \N__6461\
        );

    \I__1067\ : InMux
    port map (
            O => \N__6519\,
            I => \N__6450\
        );

    \I__1066\ : InMux
    port map (
            O => \N__6518\,
            I => \N__6450\
        );

    \I__1065\ : InMux
    port map (
            O => \N__6517\,
            I => \N__6450\
        );

    \I__1064\ : InMux
    port map (
            O => \N__6516\,
            I => \N__6450\
        );

    \I__1063\ : InMux
    port map (
            O => \N__6515\,
            I => \N__6450\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__6512\,
            I => \N__6447\
        );

    \I__1061\ : InMux
    port map (
            O => \N__6509\,
            I => \N__6444\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__6506\,
            I => \N__6439\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__6503\,
            I => \N__6439\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__6498\,
            I => \N__6430\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__6495\,
            I => \N__6430\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__6488\,
            I => \N__6430\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__6479\,
            I => \N__6430\
        );

    \I__1054\ : InMux
    port map (
            O => \N__6478\,
            I => \N__6424\
        );

    \I__1053\ : InMux
    port map (
            O => \N__6477\,
            I => \N__6424\
        );

    \I__1052\ : InMux
    port map (
            O => \N__6476\,
            I => \N__6421\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__6471\,
            I => \N__6416\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__6464\,
            I => \N__6416\
        );

    \I__1049\ : Span4Mux_v
    port map (
            O => \N__6461\,
            I => \N__6411\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__6450\,
            I => \N__6411\
        );

    \I__1047\ : Span4Mux_v
    port map (
            O => \N__6447\,
            I => \N__6402\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__6444\,
            I => \N__6402\
        );

    \I__1045\ : Span4Mux_v
    port map (
            O => \N__6439\,
            I => \N__6402\
        );

    \I__1044\ : Span4Mux_v
    port map (
            O => \N__6430\,
            I => \N__6402\
        );

    \I__1043\ : InMux
    port map (
            O => \N__6429\,
            I => \N__6399\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__6424\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__6421\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1040\ : Odrv12
    port map (
            O => \N__6416\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1039\ : Odrv4
    port map (
            O => \N__6411\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1038\ : Odrv4
    port map (
            O => \N__6402\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__6399\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1036\ : CascadeMux
    port map (
            O => \N__6386\,
            I => \N__6383\
        );

    \I__1035\ : InMux
    port map (
            O => \N__6383\,
            I => \N__6380\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__6380\,
            I => \U712_CHIP_RAM.N_438\
        );

    \I__1033\ : IoInMux
    port map (
            O => \N__6377\,
            I => \N__6374\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__6374\,
            I => \N__6371\
        );

    \I__1031\ : Span4Mux_s3_v
    port map (
            O => \N__6371\,
            I => \N__6367\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6370\,
            I => \N__6364\
        );

    \I__1029\ : Span4Mux_v
    port map (
            O => \N__6367\,
            I => \N__6361\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__6364\,
            I => \N__6358\
        );

    \I__1027\ : Span4Mux_h
    port map (
            O => \N__6361\,
            I => \N__6355\
        );

    \I__1026\ : Span4Mux_v
    port map (
            O => \N__6358\,
            I => \N__6352\
        );

    \I__1025\ : Odrv4
    port map (
            O => \N__6355\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1024\ : Odrv4
    port map (
            O => \N__6352\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1023\ : IoInMux
    port map (
            O => \N__6347\,
            I => \N__6344\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__6344\,
            I => \N__6341\
        );

    \I__1021\ : IoSpan4Mux
    port map (
            O => \N__6341\,
            I => \N__6338\
        );

    \I__1020\ : Span4Mux_s2_v
    port map (
            O => \N__6338\,
            I => \N__6334\
        );

    \I__1019\ : InMux
    port map (
            O => \N__6337\,
            I => \N__6331\
        );

    \I__1018\ : Sp12to4
    port map (
            O => \N__6334\,
            I => \N__6328\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__6331\,
            I => \N__6325\
        );

    \I__1016\ : Span12Mux_s8_v
    port map (
            O => \N__6328\,
            I => \N__6322\
        );

    \I__1015\ : Span4Mux_v
    port map (
            O => \N__6325\,
            I => \N__6319\
        );

    \I__1014\ : Span12Mux_v
    port map (
            O => \N__6322\,
            I => \N__6316\
        );

    \I__1013\ : Sp12to4
    port map (
            O => \N__6319\,
            I => \N__6313\
        );

    \I__1012\ : Span12Mux_h
    port map (
            O => \N__6316\,
            I => \N__6310\
        );

    \I__1011\ : Span12Mux_h
    port map (
            O => \N__6313\,
            I => \N__6307\
        );

    \I__1010\ : Odrv12
    port map (
            O => \N__6310\,
            I => \A_c_11\
        );

    \I__1009\ : Odrv12
    port map (
            O => \N__6307\,
            I => \A_c_11\
        );

    \I__1008\ : InMux
    port map (
            O => \N__6302\,
            I => \N__6299\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__6299\,
            I => \N__6296\
        );

    \I__1006\ : Span4Mux_v
    port map (
            O => \N__6296\,
            I => \N__6293\
        );

    \I__1005\ : Odrv4
    port map (
            O => \N__6293\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\
        );

    \I__1004\ : CascadeMux
    port map (
            O => \N__6290\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\
        );

    \I__1003\ : IoInMux
    port map (
            O => \N__6287\,
            I => \N__6284\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__6284\,
            I => \N__6281\
        );

    \I__1001\ : Span4Mux_s3_v
    port map (
            O => \N__6281\,
            I => \N__6278\
        );

    \I__1000\ : Span4Mux_h
    port map (
            O => \N__6278\,
            I => \N__6275\
        );

    \I__999\ : Span4Mux_h
    port map (
            O => \N__6275\,
            I => \N__6272\
        );

    \I__998\ : Sp12to4
    port map (
            O => \N__6272\,
            I => \N__6269\
        );

    \I__997\ : Span12Mux_v
    port map (
            O => \N__6269\,
            I => \N__6265\
        );

    \I__996\ : InMux
    port map (
            O => \N__6268\,
            I => \N__6262\
        );

    \I__995\ : Odrv12
    port map (
            O => \N__6265\,
            I => \LATCH_CLK_c\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__6262\,
            I => \LATCH_CLK_c\
        );

    \I__993\ : InMux
    port map (
            O => \N__6257\,
            I => \N__6254\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__6254\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_a2_0_1\
        );

    \I__991\ : CascadeMux
    port map (
            O => \N__6251\,
            I => \N__6246\
        );

    \I__990\ : InMux
    port map (
            O => \N__6250\,
            I => \N__6243\
        );

    \I__989\ : InMux
    port map (
            O => \N__6249\,
            I => \N__6240\
        );

    \I__988\ : InMux
    port map (
            O => \N__6246\,
            I => \N__6237\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__6243\,
            I => \U712_CHIP_RAM.N_533\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__6240\,
            I => \U712_CHIP_RAM.N_533\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__6237\,
            I => \U712_CHIP_RAM.N_533\
        );

    \I__984\ : CascadeMux
    port map (
            O => \N__6230\,
            I => \U712_CHIP_RAM.N_296_cascade_\
        );

    \I__983\ : CascadeMux
    port map (
            O => \N__6227\,
            I => \N__6224\
        );

    \I__982\ : InMux
    port map (
            O => \N__6224\,
            I => \N__6221\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__6221\,
            I => \N__6217\
        );

    \I__980\ : InMux
    port map (
            O => \N__6220\,
            I => \N__6214\
        );

    \I__979\ : Odrv4
    port map (
            O => \N__6217\,
            I => \U712_CHIP_RAM.N_550\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__6214\,
            I => \U712_CHIP_RAM.N_550\
        );

    \I__977\ : CascadeMux
    port map (
            O => \N__6209\,
            I => \N__6206\
        );

    \I__976\ : InMux
    port map (
            O => \N__6206\,
            I => \N__6202\
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__6205\,
            I => \N__6199\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__6202\,
            I => \N__6196\
        );

    \I__973\ : InMux
    port map (
            O => \N__6199\,
            I => \N__6187\
        );

    \I__972\ : Span4Mux_v
    port map (
            O => \N__6196\,
            I => \N__6184\
        );

    \I__971\ : InMux
    port map (
            O => \N__6195\,
            I => \N__6177\
        );

    \I__970\ : InMux
    port map (
            O => \N__6194\,
            I => \N__6177\
        );

    \I__969\ : InMux
    port map (
            O => \N__6193\,
            I => \N__6177\
        );

    \I__968\ : InMux
    port map (
            O => \N__6192\,
            I => \N__6170\
        );

    \I__967\ : InMux
    port map (
            O => \N__6191\,
            I => \N__6170\
        );

    \I__966\ : InMux
    port map (
            O => \N__6190\,
            I => \N__6170\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__6187\,
            I => \U712_CHIP_RAM.N_463\
        );

    \I__964\ : Odrv4
    port map (
            O => \N__6184\,
            I => \U712_CHIP_RAM.N_463\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__6177\,
            I => \U712_CHIP_RAM.N_463\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__6170\,
            I => \U712_CHIP_RAM.N_463\
        );

    \I__961\ : InMux
    port map (
            O => \N__6161\,
            I => \N__6158\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__6158\,
            I => \N__6154\
        );

    \I__959\ : InMux
    port map (
            O => \N__6157\,
            I => \N__6151\
        );

    \I__958\ : Span4Mux_h
    port map (
            O => \N__6154\,
            I => \N__6148\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__6151\,
            I => \N__6145\
        );

    \I__956\ : Odrv4
    port map (
            O => \N__6148\,
            I => \U712_CHIP_RAM.N_546\
        );

    \I__955\ : Odrv4
    port map (
            O => \N__6145\,
            I => \U712_CHIP_RAM.N_546\
        );

    \I__954\ : InMux
    port map (
            O => \N__6140\,
            I => \N__6137\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__6137\,
            I => \N__6134\
        );

    \I__952\ : Span4Mux_h
    port map (
            O => \N__6134\,
            I => \N__6122\
        );

    \I__951\ : InMux
    port map (
            O => \N__6133\,
            I => \N__6119\
        );

    \I__950\ : InMux
    port map (
            O => \N__6132\,
            I => \N__6116\
        );

    \I__949\ : InMux
    port map (
            O => \N__6131\,
            I => \N__6111\
        );

    \I__948\ : InMux
    port map (
            O => \N__6130\,
            I => \N__6111\
        );

    \I__947\ : InMux
    port map (
            O => \N__6129\,
            I => \N__6106\
        );

    \I__946\ : InMux
    port map (
            O => \N__6128\,
            I => \N__6106\
        );

    \I__945\ : InMux
    port map (
            O => \N__6127\,
            I => \N__6099\
        );

    \I__944\ : InMux
    port map (
            O => \N__6126\,
            I => \N__6099\
        );

    \I__943\ : InMux
    port map (
            O => \N__6125\,
            I => \N__6099\
        );

    \I__942\ : Odrv4
    port map (
            O => \N__6122\,
            I => \U712_CHIP_RAM.N_464\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__6119\,
            I => \U712_CHIP_RAM.N_464\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__6116\,
            I => \U712_CHIP_RAM.N_464\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__6111\,
            I => \U712_CHIP_RAM.N_464\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__6106\,
            I => \U712_CHIP_RAM.N_464\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__6099\,
            I => \U712_CHIP_RAM.N_464\
        );

    \I__936\ : InMux
    port map (
            O => \N__6086\,
            I => \N__6081\
        );

    \I__935\ : InMux
    port map (
            O => \N__6085\,
            I => \N__6078\
        );

    \I__934\ : InMux
    port map (
            O => \N__6084\,
            I => \N__6075\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__6081\,
            I => \U712_CHIP_RAM.N_465\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__6078\,
            I => \U712_CHIP_RAM.N_465\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__6075\,
            I => \U712_CHIP_RAM.N_465\
        );

    \I__930\ : CascadeMux
    port map (
            O => \N__6068\,
            I => \U712_CHIP_RAM.N_465_cascade_\
        );

    \I__929\ : InMux
    port map (
            O => \N__6065\,
            I => \N__6062\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__6062\,
            I => \N__6059\
        );

    \I__927\ : Span12Mux_v
    port map (
            O => \N__6059\,
            I => \N__6056\
        );

    \I__926\ : Span12Mux_h
    port map (
            O => \N__6056\,
            I => \N__6053\
        );

    \I__925\ : Odrv12
    port map (
            O => \N__6053\,
            I => \A_c_20\
        );

    \I__924\ : InMux
    port map (
            O => \N__6050\,
            I => \N__6047\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__6047\,
            I => \N__6043\
        );

    \I__922\ : InMux
    port map (
            O => \N__6046\,
            I => \N__6040\
        );

    \I__921\ : Odrv4
    port map (
            O => \N__6043\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__6040\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\
        );

    \I__919\ : InMux
    port map (
            O => \N__6035\,
            I => \N__6031\
        );

    \I__918\ : InMux
    port map (
            O => \N__6034\,
            I => \N__6028\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__6031\,
            I => \N__6025\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__6028\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\
        );

    \I__915\ : Odrv12
    port map (
            O => \N__6025\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\
        );

    \I__914\ : InMux
    port map (
            O => \N__6020\,
            I => \N__6017\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__6017\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0\
        );

    \I__912\ : CascadeMux
    port map (
            O => \N__6014\,
            I => \N__6011\
        );

    \I__911\ : InMux
    port map (
            O => \N__6011\,
            I => \N__6008\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__6008\,
            I => \N__6005\
        );

    \I__909\ : Odrv4
    port map (
            O => \N__6005\,
            I => \U712_CHIP_RAM.DBENn_8_0_0\
        );

    \I__908\ : IoInMux
    port map (
            O => \N__6002\,
            I => \N__5999\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__5999\,
            I => \N__5996\
        );

    \I__906\ : Span4Mux_s2_v
    port map (
            O => \N__5996\,
            I => \N__5993\
        );

    \I__905\ : Span4Mux_v
    port map (
            O => \N__5993\,
            I => \N__5990\
        );

    \I__904\ : Span4Mux_v
    port map (
            O => \N__5990\,
            I => \N__5987\
        );

    \I__903\ : Span4Mux_v
    port map (
            O => \N__5987\,
            I => \N__5983\
        );

    \I__902\ : InMux
    port map (
            O => \N__5986\,
            I => \N__5980\
        );

    \I__901\ : Odrv4
    port map (
            O => \N__5983\,
            I => \DBDIR_c\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__5980\,
            I => \DBDIR_c\
        );

    \I__899\ : IoInMux
    port map (
            O => \N__5975\,
            I => \N__5971\
        );

    \I__898\ : IoInMux
    port map (
            O => \N__5974\,
            I => \N__5968\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__5971\,
            I => \N__5965\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__5968\,
            I => \N__5962\
        );

    \I__895\ : Span4Mux_s0_v
    port map (
            O => \N__5965\,
            I => \N__5959\
        );

    \I__894\ : Span4Mux_s3_v
    port map (
            O => \N__5962\,
            I => \N__5956\
        );

    \I__893\ : Span4Mux_v
    port map (
            O => \N__5959\,
            I => \N__5953\
        );

    \I__892\ : Span4Mux_h
    port map (
            O => \N__5956\,
            I => \N__5950\
        );

    \I__891\ : Sp12to4
    port map (
            O => \N__5953\,
            I => \N__5946\
        );

    \I__890\ : Span4Mux_h
    port map (
            O => \N__5950\,
            I => \N__5943\
        );

    \I__889\ : IoInMux
    port map (
            O => \N__5949\,
            I => \N__5940\
        );

    \I__888\ : Span12Mux_s11_h
    port map (
            O => \N__5946\,
            I => \N__5935\
        );

    \I__887\ : Sp12to4
    port map (
            O => \N__5943\,
            I => \N__5935\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__5940\,
            I => \N__5932\
        );

    \I__885\ : Span12Mux_v
    port map (
            O => \N__5935\,
            I => \N__5927\
        );

    \I__884\ : Span12Mux_s8_h
    port map (
            O => \N__5932\,
            I => \N__5927\
        );

    \I__883\ : Odrv12
    port map (
            O => \N__5927\,
            I => \CLK40_PLL_i_i\
        );

    \I__882\ : IoInMux
    port map (
            O => \N__5924\,
            I => \N__5921\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__5921\,
            I => \N__5918\
        );

    \I__880\ : IoSpan4Mux
    port map (
            O => \N__5918\,
            I => \N__5915\
        );

    \I__879\ : Span4Mux_s3_v
    port map (
            O => \N__5915\,
            I => \N__5912\
        );

    \I__878\ : Span4Mux_v
    port map (
            O => \N__5912\,
            I => \N__5909\
        );

    \I__877\ : Odrv4
    port map (
            O => \N__5909\,
            I => \N_167_i\
        );

    \I__876\ : CascadeMux
    port map (
            O => \N__5906\,
            I => \U712_CHIP_RAM.N_533_cascade_\
        );

    \I__875\ : InMux
    port map (
            O => \N__5903\,
            I => \N__5900\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__5900\,
            I => \U712_CHIP_RAM.N_370\
        );

    \I__873\ : CascadeMux
    port map (
            O => \N__5897\,
            I => \U712_CHIP_RAM.N_391_cascade_\
        );

    \I__872\ : CascadeMux
    port map (
            O => \N__5894\,
            I => \N__5891\
        );

    \I__871\ : InMux
    port map (
            O => \N__5891\,
            I => \N__5888\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__5888\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0\
        );

    \I__869\ : IoInMux
    port map (
            O => \N__5885\,
            I => \N__5882\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__5882\,
            I => \N__5879\
        );

    \I__867\ : Span12Mux_s6_h
    port map (
            O => \N__5879\,
            I => \N__5876\
        );

    \I__866\ : Span12Mux_h
    port map (
            O => \N__5876\,
            I => \N__5873\
        );

    \I__865\ : Odrv12
    port map (
            O => \N__5873\,
            I => \CLK_EN_c\
        );

    \I__864\ : InMux
    port map (
            O => \N__5870\,
            I => \N__5866\
        );

    \I__863\ : InMux
    port map (
            O => \N__5869\,
            I => \N__5863\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__5866\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__5863\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__860\ : InMux
    port map (
            O => \N__5858\,
            I => \N__5854\
        );

    \I__859\ : InMux
    port map (
            O => \N__5857\,
            I => \N__5851\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5854\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__5851\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__856\ : CascadeMux
    port map (
            O => \N__5846\,
            I => \N__5842\
        );

    \I__855\ : InMux
    port map (
            O => \N__5845\,
            I => \N__5839\
        );

    \I__854\ : InMux
    port map (
            O => \N__5842\,
            I => \N__5836\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__5839\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__5836\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__851\ : InMux
    port map (
            O => \N__5831\,
            I => \N__5827\
        );

    \I__850\ : InMux
    port map (
            O => \N__5830\,
            I => \N__5824\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__5827\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__5824\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__847\ : CascadeMux
    port map (
            O => \N__5819\,
            I => \U712_CHIP_RAM.N_295_cascade_\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__5816\,
            I => \N__5812\
        );

    \I__845\ : InMux
    port map (
            O => \N__5815\,
            I => \N__5807\
        );

    \I__844\ : InMux
    port map (
            O => \N__5812\,
            I => \N__5807\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__5807\,
            I => \N__5802\
        );

    \I__842\ : InMux
    port map (
            O => \N__5806\,
            I => \N__5794\
        );

    \I__841\ : InMux
    port map (
            O => \N__5805\,
            I => \N__5791\
        );

    \I__840\ : Span4Mux_h
    port map (
            O => \N__5802\,
            I => \N__5788\
        );

    \I__839\ : InMux
    port map (
            O => \N__5801\,
            I => \N__5785\
        );

    \I__838\ : InMux
    port map (
            O => \N__5800\,
            I => \N__5782\
        );

    \I__837\ : InMux
    port map (
            O => \N__5799\,
            I => \N__5777\
        );

    \I__836\ : InMux
    port map (
            O => \N__5798\,
            I => \N__5777\
        );

    \I__835\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5774\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__5794\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__5791\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__832\ : Odrv4
    port map (
            O => \N__5788\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__5785\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__5782\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__5777\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__5774\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__827\ : CascadeMux
    port map (
            O => \N__5759\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_cascade_\
        );

    \I__826\ : InMux
    port map (
            O => \N__5756\,
            I => \N__5753\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__5753\,
            I => \N__5749\
        );

    \I__824\ : InMux
    port map (
            O => \N__5752\,
            I => \N__5746\
        );

    \I__823\ : Span4Mux_v
    port map (
            O => \N__5749\,
            I => \N__5738\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__5746\,
            I => \N__5738\
        );

    \I__821\ : InMux
    port map (
            O => \N__5745\,
            I => \N__5733\
        );

    \I__820\ : InMux
    port map (
            O => \N__5744\,
            I => \N__5733\
        );

    \I__819\ : InMux
    port map (
            O => \N__5743\,
            I => \N__5730\
        );

    \I__818\ : Odrv4
    port map (
            O => \N__5738\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__5733\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__5730\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__815\ : CascadeMux
    port map (
            O => \N__5723\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_cascade_\
        );

    \I__814\ : CEMux
    port map (
            O => \N__5720\,
            I => \N__5717\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__5717\,
            I => \N__5714\
        );

    \I__812\ : Span4Mux_h
    port map (
            O => \N__5714\,
            I => \N__5711\
        );

    \I__811\ : Odrv4
    port map (
            O => \N__5711\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_1\
        );

    \I__810\ : InMux
    port map (
            O => \N__5708\,
            I => \N__5704\
        );

    \I__809\ : InMux
    port map (
            O => \N__5707\,
            I => \N__5700\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__5704\,
            I => \N__5693\
        );

    \I__807\ : InMux
    port map (
            O => \N__5703\,
            I => \N__5690\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__5700\,
            I => \N__5687\
        );

    \I__805\ : InMux
    port map (
            O => \N__5699\,
            I => \N__5684\
        );

    \I__804\ : InMux
    port map (
            O => \N__5698\,
            I => \N__5679\
        );

    \I__803\ : InMux
    port map (
            O => \N__5697\,
            I => \N__5679\
        );

    \I__802\ : CascadeMux
    port map (
            O => \N__5696\,
            I => \N__5674\
        );

    \I__801\ : Span4Mux_h
    port map (
            O => \N__5693\,
            I => \N__5671\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__5690\,
            I => \N__5666\
        );

    \I__799\ : Span4Mux_h
    port map (
            O => \N__5687\,
            I => \N__5666\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__5684\,
            I => \N__5661\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5679\,
            I => \N__5661\
        );

    \I__796\ : InMux
    port map (
            O => \N__5678\,
            I => \N__5658\
        );

    \I__795\ : InMux
    port map (
            O => \N__5677\,
            I => \N__5653\
        );

    \I__794\ : InMux
    port map (
            O => \N__5674\,
            I => \N__5653\
        );

    \I__793\ : Odrv4
    port map (
            O => \N__5671\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__792\ : Odrv4
    port map (
            O => \N__5666\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__791\ : Odrv4
    port map (
            O => \N__5661\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__5658\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__5653\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__788\ : CascadeMux
    port map (
            O => \N__5642\,
            I => \U712_CHIP_RAM.N_463_cascade_\
        );

    \I__787\ : CascadeMux
    port map (
            O => \N__5639\,
            I => \N__5636\
        );

    \I__786\ : InMux
    port map (
            O => \N__5636\,
            I => \N__5632\
        );

    \I__785\ : InMux
    port map (
            O => \N__5635\,
            I => \N__5629\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__5632\,
            I => \N__5625\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__5629\,
            I => \N__5622\
        );

    \I__782\ : CascadeMux
    port map (
            O => \N__5628\,
            I => \N__5619\
        );

    \I__781\ : Span4Mux_h
    port map (
            O => \N__5625\,
            I => \N__5615\
        );

    \I__780\ : Span4Mux_h
    port map (
            O => \N__5622\,
            I => \N__5612\
        );

    \I__779\ : InMux
    port map (
            O => \N__5619\,
            I => \N__5607\
        );

    \I__778\ : InMux
    port map (
            O => \N__5618\,
            I => \N__5607\
        );

    \I__777\ : Odrv4
    port map (
            O => \N__5615\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__776\ : Odrv4
    port map (
            O => \N__5612\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__5607\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__774\ : CascadeMux
    port map (
            O => \N__5600\,
            I => \U712_CHIP_RAM.N_385_cascade_\
        );

    \I__773\ : InMux
    port map (
            O => \N__5597\,
            I => \N__5594\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__5594\,
            I => \U712_CHIP_RAM.N_384\
        );

    \I__771\ : CascadeMux
    port map (
            O => \N__5591\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0_cascade_\
        );

    \I__770\ : InMux
    port map (
            O => \N__5588\,
            I => \N__5585\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__5585\,
            I => \U712_CHIP_RAM.N_461\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__5582\,
            I => \N__5579\
        );

    \I__767\ : InMux
    port map (
            O => \N__5579\,
            I => \N__5576\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__5576\,
            I => \N__5573\
        );

    \I__765\ : Span4Mux_v
    port map (
            O => \N__5573\,
            I => \N__5568\
        );

    \I__764\ : InMux
    port map (
            O => \N__5572\,
            I => \N__5563\
        );

    \I__763\ : InMux
    port map (
            O => \N__5571\,
            I => \N__5563\
        );

    \I__762\ : Odrv4
    port map (
            O => \N__5568\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__5563\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\
        );

    \I__760\ : CascadeMux
    port map (
            O => \N__5558\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERlde_0_a3_0_0_a2_0_cascade_\
        );

    \I__759\ : CEMux
    port map (
            O => \N__5555\,
            I => \N__5550\
        );

    \I__758\ : CEMux
    port map (
            O => \N__5554\,
            I => \N__5547\
        );

    \I__757\ : CEMux
    port map (
            O => \N__5553\,
            I => \N__5544\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__5550\,
            I => \N__5541\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__5547\,
            I => \N__5538\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__5544\,
            I => \N__5535\
        );

    \I__753\ : Span4Mux_h
    port map (
            O => \N__5541\,
            I => \N__5530\
        );

    \I__752\ : Span4Mux_h
    port map (
            O => \N__5538\,
            I => \N__5530\
        );

    \I__751\ : Span4Mux_v
    port map (
            O => \N__5535\,
            I => \N__5527\
        );

    \I__750\ : Odrv4
    port map (
            O => \N__5530\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__749\ : Odrv4
    port map (
            O => \N__5527\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__748\ : InMux
    port map (
            O => \N__5522\,
            I => \N__5519\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__5519\,
            I => \N__5516\
        );

    \I__746\ : Span4Mux_h
    port map (
            O => \N__5516\,
            I => \N__5513\
        );

    \I__745\ : Odrv4
    port map (
            O => \N__5513\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERlde_0_a3_0_0_a2_0\
        );

    \I__744\ : CascadeMux
    port map (
            O => \N__5510\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_1_cascade_\
        );

    \I__743\ : InMux
    port map (
            O => \N__5507\,
            I => \N__5504\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__5504\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__741\ : CascadeMux
    port map (
            O => \N__5501\,
            I => \N__5495\
        );

    \I__740\ : CascadeMux
    port map (
            O => \N__5500\,
            I => \N__5492\
        );

    \I__739\ : InMux
    port map (
            O => \N__5499\,
            I => \N__5482\
        );

    \I__738\ : InMux
    port map (
            O => \N__5498\,
            I => \N__5482\
        );

    \I__737\ : InMux
    port map (
            O => \N__5495\,
            I => \N__5482\
        );

    \I__736\ : InMux
    port map (
            O => \N__5492\,
            I => \N__5482\
        );

    \I__735\ : InMux
    port map (
            O => \N__5491\,
            I => \N__5477\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__5482\,
            I => \N__5474\
        );

    \I__733\ : InMux
    port map (
            O => \N__5481\,
            I => \N__5471\
        );

    \I__732\ : InMux
    port map (
            O => \N__5480\,
            I => \N__5468\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__5477\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__730\ : Odrv4
    port map (
            O => \N__5474\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__5471\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__5468\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__727\ : InMux
    port map (
            O => \N__5459\,
            I => \N__5456\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__5456\,
            I => \U712_CHIP_RAM.N_419\
        );

    \I__725\ : InMux
    port map (
            O => \N__5453\,
            I => \N__5450\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__5450\,
            I => \N__5447\
        );

    \I__723\ : Odrv12
    port map (
            O => \N__5447\,
            I => \U712_BYTE_ENABLE.N_326\
        );

    \I__722\ : InMux
    port map (
            O => \N__5444\,
            I => \N__5441\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__5441\,
            I => \N__5438\
        );

    \I__720\ : Odrv4
    port map (
            O => \N__5438\,
            I => \U712_BYTE_ENABLE.N_323\
        );

    \I__719\ : InMux
    port map (
            O => \N__5435\,
            I => \N__5432\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__5432\,
            I => \N__5429\
        );

    \I__717\ : Odrv12
    port map (
            O => \N__5429\,
            I => \U712_BYTE_ENABLE.N_324\
        );

    \I__716\ : InMux
    port map (
            O => \N__5426\,
            I => \N__5423\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__5423\,
            I => \N__5420\
        );

    \I__714\ : Span4Mux_h
    port map (
            O => \N__5420\,
            I => \N__5417\
        );

    \I__713\ : Sp12to4
    port map (
            O => \N__5417\,
            I => \N__5414\
        );

    \I__712\ : Span12Mux_v
    port map (
            O => \N__5414\,
            I => \N__5411\
        );

    \I__711\ : Odrv12
    port map (
            O => \N__5411\,
            I => \A_c_17\
        );

    \I__710\ : InMux
    port map (
            O => \N__5408\,
            I => \N__5399\
        );

    \I__709\ : InMux
    port map (
            O => \N__5407\,
            I => \N__5392\
        );

    \I__708\ : InMux
    port map (
            O => \N__5406\,
            I => \N__5392\
        );

    \I__707\ : InMux
    port map (
            O => \N__5405\,
            I => \N__5392\
        );

    \I__706\ : InMux
    port map (
            O => \N__5404\,
            I => \N__5385\
        );

    \I__705\ : InMux
    port map (
            O => \N__5403\,
            I => \N__5385\
        );

    \I__704\ : InMux
    port map (
            O => \N__5402\,
            I => \N__5385\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__5399\,
            I => \N__5382\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__5392\,
            I => \U712_CHIP_RAM.N_90_i\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__5385\,
            I => \U712_CHIP_RAM.N_90_i\
        );

    \I__700\ : Odrv4
    port map (
            O => \N__5382\,
            I => \U712_CHIP_RAM.N_90_i\
        );

    \I__699\ : InMux
    port map (
            O => \N__5375\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__698\ : IoInMux
    port map (
            O => \N__5372\,
            I => \N__5369\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__5369\,
            I => \N__5366\
        );

    \I__696\ : IoSpan4Mux
    port map (
            O => \N__5366\,
            I => \N__5363\
        );

    \I__695\ : Span4Mux_s2_v
    port map (
            O => \N__5363\,
            I => \N__5360\
        );

    \I__694\ : Sp12to4
    port map (
            O => \N__5360\,
            I => \N__5357\
        );

    \I__693\ : Odrv12
    port map (
            O => \N__5357\,
            I => \N_188_i\
        );

    \I__692\ : InMux
    port map (
            O => \N__5354\,
            I => \N__5350\
        );

    \I__691\ : InMux
    port map (
            O => \N__5353\,
            I => \N__5347\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__5350\,
            I => \N__5342\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__5347\,
            I => \N__5342\
        );

    \I__688\ : Odrv4
    port map (
            O => \N__5342\,
            I => \U712_CHIP_RAM.N_302\
        );

    \I__687\ : CascadeMux
    port map (
            O => \N__5339\,
            I => \N__5336\
        );

    \I__686\ : InMux
    port map (
            O => \N__5336\,
            I => \N__5332\
        );

    \I__685\ : InMux
    port map (
            O => \N__5335\,
            I => \N__5329\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__5332\,
            I => \N__5324\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__5329\,
            I => \N__5324\
        );

    \I__682\ : Span4Mux_v
    port map (
            O => \N__5324\,
            I => \N__5321\
        );

    \I__681\ : Odrv4
    port map (
            O => \N__5321\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3\
        );

    \I__680\ : InMux
    port map (
            O => \N__5318\,
            I => \N__5315\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__5315\,
            I => \U712_CHIP_RAM.N_455\
        );

    \I__678\ : CascadeMux
    port map (
            O => \N__5312\,
            I => \U712_CHIP_RAM.N_417_cascade_\
        );

    \I__677\ : InMux
    port map (
            O => \N__5309\,
            I => \N__5306\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__5306\,
            I => \N__5303\
        );

    \I__675\ : Span12Mux_h
    port map (
            O => \N__5303\,
            I => \N__5300\
        );

    \I__674\ : Span12Mux_v
    port map (
            O => \N__5300\,
            I => \N__5297\
        );

    \I__673\ : Odrv12
    port map (
            O => \N__5297\,
            I => \RAMSPACEn_c\
        );

    \I__672\ : InMux
    port map (
            O => \N__5294\,
            I => \N__5291\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__5291\,
            I => \N__5285\
        );

    \I__670\ : InMux
    port map (
            O => \N__5290\,
            I => \N__5278\
        );

    \I__669\ : InMux
    port map (
            O => \N__5289\,
            I => \N__5278\
        );

    \I__668\ : InMux
    port map (
            O => \N__5288\,
            I => \N__5278\
        );

    \I__667\ : Odrv4
    port map (
            O => \N__5285\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__5278\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__665\ : InMux
    port map (
            O => \N__5273\,
            I => \N__5270\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__5270\,
            I => \N__5266\
        );

    \I__663\ : InMux
    port map (
            O => \N__5269\,
            I => \N__5263\
        );

    \I__662\ : Span4Mux_h
    port map (
            O => \N__5266\,
            I => \N__5260\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__5263\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__660\ : Odrv4
    port map (
            O => \N__5260\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__659\ : InMux
    port map (
            O => \N__5255\,
            I => \N__5252\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__5252\,
            I => \N__5249\
        );

    \I__657\ : Span4Mux_h
    port map (
            O => \N__5249\,
            I => \N__5246\
        );

    \I__656\ : Odrv4
    port map (
            O => \N__5246\,
            I => \U712_CHIP_RAM.REFRESH5lto7_0\
        );

    \I__655\ : InMux
    port map (
            O => \N__5243\,
            I => \N__5240\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__5240\,
            I => \N__5237\
        );

    \I__653\ : Span4Mux_h
    port map (
            O => \N__5237\,
            I => \N__5234\
        );

    \I__652\ : Odrv4
    port map (
            O => \N__5234\,
            I => \U712_CHIP_RAM.REFRESH5lt7\
        );

    \I__651\ : InMux
    port map (
            O => \N__5231\,
            I => \N__5228\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__5228\,
            I => \N__5224\
        );

    \I__649\ : InMux
    port map (
            O => \N__5227\,
            I => \N__5221\
        );

    \I__648\ : Odrv4
    port map (
            O => \N__5224\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_o2_0_0\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__5221\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_o2_0_0\
        );

    \I__646\ : InMux
    port map (
            O => \N__5216\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__645\ : InMux
    port map (
            O => \N__5213\,
            I => \N__5210\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__5210\,
            I => \N__5207\
        );

    \I__643\ : Odrv4
    port map (
            O => \N__5207\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__642\ : InMux
    port map (
            O => \N__5204\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__641\ : InMux
    port map (
            O => \N__5201\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__640\ : InMux
    port map (
            O => \N__5198\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__639\ : InMux
    port map (
            O => \N__5195\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__638\ : InMux
    port map (
            O => \N__5192\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__637\ : InMux
    port map (
            O => \N__5189\,
            I => \N__5183\
        );

    \I__636\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5183\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__5183\,
            I => \N__5180\
        );

    \I__634\ : Odrv4
    port map (
            O => \N__5180\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0\
        );

    \I__633\ : IoInMux
    port map (
            O => \N__5177\,
            I => \N__5174\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__5174\,
            I => \N__5171\
        );

    \I__631\ : IoSpan4Mux
    port map (
            O => \N__5171\,
            I => \N__5168\
        );

    \I__630\ : Sp12to4
    port map (
            O => \N__5168\,
            I => \N__5165\
        );

    \I__629\ : Span12Mux_s7_h
    port map (
            O => \N__5165\,
            I => \N__5162\
        );

    \I__628\ : Odrv12
    port map (
            O => \N__5162\,
            I => \N_176_i\
        );

    \I__627\ : InMux
    port map (
            O => \N__5159\,
            I => \N__5156\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__5156\,
            I => \N__5153\
        );

    \I__625\ : Odrv12
    port map (
            O => \N__5153\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\
        );

    \I__624\ : InMux
    port map (
            O => \N__5150\,
            I => \N__5147\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__5147\,
            I => \N__5144\
        );

    \I__622\ : Span4Mux_v
    port map (
            O => \N__5144\,
            I => \N__5141\
        );

    \I__621\ : Span4Mux_h
    port map (
            O => \N__5141\,
            I => \N__5138\
        );

    \I__620\ : Sp12to4
    port map (
            O => \N__5138\,
            I => \N__5135\
        );

    \I__619\ : Odrv12
    port map (
            O => \N__5135\,
            I => \A_c_12\
        );

    \I__618\ : InMux
    port map (
            O => \N__5132\,
            I => \N__5129\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__5129\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER19\
        );

    \I__616\ : CascadeMux
    port map (
            O => \N__5126\,
            I => \U712_CHIP_RAM.N_464_cascade_\
        );

    \I__615\ : CascadeMux
    port map (
            O => \N__5123\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_\
        );

    \I__614\ : InMux
    port map (
            O => \N__5120\,
            I => \N__5117\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__5117\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0\
        );

    \I__612\ : InMux
    port map (
            O => \N__5114\,
            I => \N__5111\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__5111\,
            I => \U712_CHIP_RAM.N_390\
        );

    \I__610\ : InMux
    port map (
            O => \N__5108\,
            I => \N__5105\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__5105\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0\
        );

    \I__608\ : InMux
    port map (
            O => \N__5102\,
            I => \N__5098\
        );

    \I__607\ : InMux
    port map (
            O => \N__5101\,
            I => \N__5095\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__5098\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__5095\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\
        );

    \I__604\ : CascadeMux
    port map (
            O => \N__5090\,
            I => \N__5087\
        );

    \I__603\ : InMux
    port map (
            O => \N__5087\,
            I => \N__5084\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__5084\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3\
        );

    \I__601\ : InMux
    port map (
            O => \N__5081\,
            I => \N__5077\
        );

    \I__600\ : InMux
    port map (
            O => \N__5080\,
            I => \N__5074\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__5077\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__5074\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\
        );

    \I__597\ : InMux
    port map (
            O => \N__5069\,
            I => \N__5065\
        );

    \I__596\ : CascadeMux
    port map (
            O => \N__5068\,
            I => \N__5062\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__5065\,
            I => \N__5059\
        );

    \I__594\ : InMux
    port map (
            O => \N__5062\,
            I => \N__5056\
        );

    \I__593\ : Odrv4
    port map (
            O => \N__5059\,
            I => \DBR_SYNC_i_1\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__5056\,
            I => \DBR_SYNC_i_1\
        );

    \I__591\ : InMux
    port map (
            O => \N__5051\,
            I => \N__5048\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__5048\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__589\ : InMux
    port map (
            O => \N__5045\,
            I => \N__5042\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__5042\,
            I => \N__5039\
        );

    \I__587\ : Span4Mux_h
    port map (
            O => \N__5039\,
            I => \N__5036\
        );

    \I__586\ : Sp12to4
    port map (
            O => \N__5036\,
            I => \N__5033\
        );

    \I__585\ : Span12Mux_v
    port map (
            O => \N__5033\,
            I => \N__5030\
        );

    \I__584\ : Odrv12
    port map (
            O => \N__5030\,
            I => \A_c_5\
        );

    \I__583\ : CEMux
    port map (
            O => \N__5027\,
            I => \N__5023\
        );

    \I__582\ : CEMux
    port map (
            O => \N__5026\,
            I => \N__5018\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__5023\,
            I => \N__5015\
        );

    \I__580\ : CEMux
    port map (
            O => \N__5022\,
            I => \N__5012\
        );

    \I__579\ : CEMux
    port map (
            O => \N__5021\,
            I => \N__5009\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__5018\,
            I => \N__5006\
        );

    \I__577\ : Span4Mux_v
    port map (
            O => \N__5015\,
            I => \N__5001\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__5012\,
            I => \N__5001\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__5009\,
            I => \N__4998\
        );

    \I__574\ : Span4Mux_h
    port map (
            O => \N__5006\,
            I => \N__4995\
        );

    \I__573\ : Span4Mux_h
    port map (
            O => \N__5001\,
            I => \N__4992\
        );

    \I__572\ : Span4Mux_v
    port map (
            O => \N__4998\,
            I => \N__4989\
        );

    \I__571\ : Odrv4
    port map (
            O => \N__4995\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\
        );

    \I__570\ : Odrv4
    port map (
            O => \N__4992\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\
        );

    \I__569\ : Odrv4
    port map (
            O => \N__4989\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\
        );

    \I__568\ : InMux
    port map (
            O => \N__4982\,
            I => \N__4979\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__4979\,
            I => \N__4976\
        );

    \I__566\ : Sp12to4
    port map (
            O => \N__4976\,
            I => \N__4973\
        );

    \I__565\ : Span12Mux_v
    port map (
            O => \N__4973\,
            I => \N__4970\
        );

    \I__564\ : Span12Mux_h
    port map (
            O => \N__4970\,
            I => \N__4967\
        );

    \I__563\ : Odrv12
    port map (
            O => \N__4967\,
            I => \A_c_16\
        );

    \I__562\ : InMux
    port map (
            O => \N__4964\,
            I => \N__4961\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__4961\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\
        );

    \I__560\ : InMux
    port map (
            O => \N__4958\,
            I => \N__4955\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__4955\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a3_0_a2_0\
        );

    \I__558\ : IoInMux
    port map (
            O => \N__4952\,
            I => \N__4949\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__4949\,
            I => \N__4946\
        );

    \I__556\ : IoSpan4Mux
    port map (
            O => \N__4946\,
            I => \N__4943\
        );

    \I__555\ : Sp12to4
    port map (
            O => \N__4943\,
            I => \N__4940\
        );

    \I__554\ : Span12Mux_s7_h
    port map (
            O => \N__4940\,
            I => \N__4937\
        );

    \I__553\ : Span12Mux_h
    port map (
            O => \N__4937\,
            I => \N__4934\
        );

    \I__552\ : Odrv12
    port map (
            O => \N__4934\,
            I => \N_178_i\
        );

    \I__551\ : InMux
    port map (
            O => \N__4931\,
            I => \N__4925\
        );

    \I__550\ : InMux
    port map (
            O => \N__4930\,
            I => \N__4925\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__4925\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\
        );

    \I__548\ : CascadeMux
    port map (
            O => \N__4922\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3_cascade_\
        );

    \I__547\ : InMux
    port map (
            O => \N__4919\,
            I => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\
        );

    \I__546\ : InMux
    port map (
            O => \N__4916\,
            I => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\
        );

    \I__545\ : InMux
    port map (
            O => \N__4913\,
            I => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2\
        );

    \I__544\ : InMux
    port map (
            O => \N__4910\,
            I => \N__4907\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__4907\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2\
        );

    \I__542\ : CascadeMux
    port map (
            O => \N__4904\,
            I => \N__4900\
        );

    \I__541\ : InMux
    port map (
            O => \N__4903\,
            I => \N__4897\
        );

    \I__540\ : InMux
    port map (
            O => \N__4900\,
            I => \N__4894\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__4897\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__4894\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\
        );

    \I__537\ : CascadeMux
    port map (
            O => \N__4889\,
            I => \N__4886\
        );

    \I__536\ : InMux
    port map (
            O => \N__4886\,
            I => \N__4883\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__4883\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1\
        );

    \I__534\ : InMux
    port map (
            O => \N__4880\,
            I => \N__4876\
        );

    \I__533\ : InMux
    port map (
            O => \N__4879\,
            I => \N__4873\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__4876\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ0Z_1\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__4873\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ0Z_1\
        );

    \I__530\ : CascadeMux
    port map (
            O => \N__4868\,
            I => \U712_CHIP_RAM.N_298_cascade_\
        );

    \I__529\ : CascadeMux
    port map (
            O => \N__4865\,
            I => \U712_CHIP_RAM.N_300_cascade_\
        );

    \I__528\ : InMux
    port map (
            O => \N__4862\,
            I => \N__4859\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__4859\,
            I => \N__4856\
        );

    \I__526\ : Odrv4
    port map (
            O => \N__4856\,
            I => \U712_CHIP_RAM.N_310\
        );

    \I__525\ : CascadeMux
    port map (
            O => \N__4853\,
            I => \U712_CHIP_RAM.N_310_cascade_\
        );

    \I__524\ : InMux
    port map (
            O => \N__4850\,
            I => \N__4846\
        );

    \I__523\ : InMux
    port map (
            O => \N__4849\,
            I => \N__4843\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__4846\,
            I => \U712_CHIP_RAM.N_313\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__4843\,
            I => \U712_CHIP_RAM.N_313\
        );

    \I__520\ : InMux
    port map (
            O => \N__4838\,
            I => \N__4835\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__4835\,
            I => \U712_CHIP_RAM.N_389\
        );

    \I__518\ : InMux
    port map (
            O => \N__4832\,
            I => \N__4829\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__4829\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_5\
        );

    \I__516\ : InMux
    port map (
            O => \N__4826\,
            I => \N__4823\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__4823\,
            I => \N__4820\
        );

    \I__514\ : Span4Mux_h
    port map (
            O => \N__4820\,
            I => \N__4817\
        );

    \I__513\ : Sp12to4
    port map (
            O => \N__4817\,
            I => \N__4814\
        );

    \I__512\ : Span12Mux_v
    port map (
            O => \N__4814\,
            I => \N__4811\
        );

    \I__511\ : Odrv12
    port map (
            O => \N__4811\,
            I => \A_c_18\
        );

    \I__510\ : CEMux
    port map (
            O => \N__4808\,
            I => \N__4805\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__4805\,
            I => \N__4802\
        );

    \I__508\ : Odrv4
    port map (
            O => \N__4802\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0\
        );

    \I__507\ : InMux
    port map (
            O => \N__4799\,
            I => \N__4796\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__4796\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__505\ : CascadeMux
    port map (
            O => \N__4793\,
            I => \N__4790\
        );

    \I__504\ : InMux
    port map (
            O => \N__4790\,
            I => \N__4787\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4787\,
            I => \N__4784\
        );

    \I__502\ : Odrv4
    port map (
            O => \N__4784\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_a2_1_0\
        );

    \I__501\ : CascadeMux
    port map (
            O => \N__4781\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_165_i_i_0_cascade_\
        );

    \I__500\ : InMux
    port map (
            O => \N__4778\,
            I => \N__4775\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__4775\,
            I => \N__4772\
        );

    \I__498\ : Odrv4
    port map (
            O => \N__4772\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__497\ : CascadeMux
    port map (
            O => \N__4769\,
            I => \U712_CHIP_RAM.N_90_i_cascade_\
        );

    \I__496\ : InMux
    port map (
            O => \N__4766\,
            I => \N__4763\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__4763\,
            I => \N__4760\
        );

    \I__494\ : Span4Mux_v
    port map (
            O => \N__4760\,
            I => \N__4757\
        );

    \I__493\ : Span4Mux_v
    port map (
            O => \N__4757\,
            I => \N__4754\
        );

    \I__492\ : Sp12to4
    port map (
            O => \N__4754\,
            I => \N__4751\
        );

    \I__491\ : Odrv12
    port map (
            O => \N__4751\,
            I => \A_c_7\
        );

    \I__490\ : InMux
    port map (
            O => \N__4748\,
            I => \N__4745\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__4745\,
            I => \N__4742\
        );

    \I__488\ : Span4Mux_v
    port map (
            O => \N__4742\,
            I => \N__4739\
        );

    \I__487\ : Span4Mux_v
    port map (
            O => \N__4739\,
            I => \N__4736\
        );

    \I__486\ : Sp12to4
    port map (
            O => \N__4736\,
            I => \N__4733\
        );

    \I__485\ : Odrv12
    port map (
            O => \N__4733\,
            I => \A_c_8\
        );

    \I__484\ : CEMux
    port map (
            O => \N__4730\,
            I => \N__4727\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__4727\,
            I => \N__4724\
        );

    \I__482\ : Span4Mux_v
    port map (
            O => \N__4724\,
            I => \N__4721\
        );

    \I__481\ : Odrv4
    port map (
            O => \N__4721\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0\
        );

    \I__480\ : InMux
    port map (
            O => \N__4718\,
            I => \N__4715\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4715\,
            I => \N__4711\
        );

    \I__478\ : InMux
    port map (
            O => \N__4714\,
            I => \N__4708\
        );

    \I__477\ : Span4Mux_v
    port map (
            O => \N__4711\,
            I => \N__4703\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__4708\,
            I => \N__4703\
        );

    \I__475\ : Span4Mux_v
    port map (
            O => \N__4703\,
            I => \N__4700\
        );

    \I__474\ : Sp12to4
    port map (
            O => \N__4700\,
            I => \N__4697\
        );

    \I__473\ : Span12Mux_h
    port map (
            O => \N__4697\,
            I => \N__4694\
        );

    \I__472\ : Odrv12
    port map (
            O => \N__4694\,
            I => \DBRn_c\
        );

    \I__471\ : IoInMux
    port map (
            O => \N__4691\,
            I => \N__4688\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__4688\,
            I => \N__4685\
        );

    \I__469\ : Span12Mux_s9_v
    port map (
            O => \N__4685\,
            I => \N__4682\
        );

    \I__468\ : Odrv12
    port map (
            O => \N__4682\,
            I => \VBENn_c\
        );

    \I__467\ : InMux
    port map (
            O => \N__4679\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__466\ : InMux
    port map (
            O => \N__4676\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__465\ : ClkMux
    port map (
            O => \N__4673\,
            I => \N__4649\
        );

    \I__464\ : ClkMux
    port map (
            O => \N__4672\,
            I => \N__4649\
        );

    \I__463\ : ClkMux
    port map (
            O => \N__4671\,
            I => \N__4649\
        );

    \I__462\ : ClkMux
    port map (
            O => \N__4670\,
            I => \N__4649\
        );

    \I__461\ : ClkMux
    port map (
            O => \N__4669\,
            I => \N__4649\
        );

    \I__460\ : ClkMux
    port map (
            O => \N__4668\,
            I => \N__4649\
        );

    \I__459\ : ClkMux
    port map (
            O => \N__4667\,
            I => \N__4649\
        );

    \I__458\ : ClkMux
    port map (
            O => \N__4666\,
            I => \N__4649\
        );

    \I__457\ : GlobalMux
    port map (
            O => \N__4649\,
            I => \N__4646\
        );

    \I__456\ : gio2CtrlBuf
    port map (
            O => \N__4646\,
            I => \C1_c_g\
        );

    \I__455\ : InMux
    port map (
            O => \N__4643\,
            I => \N__4639\
        );

    \I__454\ : InMux
    port map (
            O => \N__4642\,
            I => \N__4636\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__4639\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__4636\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__451\ : InMux
    port map (
            O => \N__4631\,
            I => \N__4627\
        );

    \I__450\ : InMux
    port map (
            O => \N__4630\,
            I => \N__4624\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__4627\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__4624\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__447\ : CascadeMux
    port map (
            O => \N__4619\,
            I => \N__4615\
        );

    \I__446\ : InMux
    port map (
            O => \N__4618\,
            I => \N__4612\
        );

    \I__445\ : InMux
    port map (
            O => \N__4615\,
            I => \N__4609\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__4612\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__4609\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__442\ : InMux
    port map (
            O => \N__4604\,
            I => \N__4600\
        );

    \I__441\ : InMux
    port map (
            O => \N__4603\,
            I => \N__4597\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__4600\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__4597\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__438\ : InMux
    port map (
            O => \N__4592\,
            I => \N__4588\
        );

    \I__437\ : InMux
    port map (
            O => \N__4591\,
            I => \N__4585\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__4588\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__4585\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__434\ : InMux
    port map (
            O => \N__4580\,
            I => \N__4576\
        );

    \I__433\ : InMux
    port map (
            O => \N__4579\,
            I => \N__4573\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__4576\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__4573\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__430\ : InMux
    port map (
            O => \N__4568\,
            I => \N__4565\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__4565\,
            I => \N__4562\
        );

    \I__428\ : Span4Mux_v
    port map (
            O => \N__4562\,
            I => \N__4559\
        );

    \I__427\ : Span4Mux_v
    port map (
            O => \N__4559\,
            I => \N__4556\
        );

    \I__426\ : Sp12to4
    port map (
            O => \N__4556\,
            I => \N__4553\
        );

    \I__425\ : Odrv12
    port map (
            O => \N__4553\,
            I => \A_c_6\
        );

    \I__424\ : InMux
    port map (
            O => \N__4550\,
            I => \N__4547\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__4547\,
            I => \N__4544\
        );

    \I__422\ : Span4Mux_v
    port map (
            O => \N__4544\,
            I => \N__4541\
        );

    \I__421\ : Sp12to4
    port map (
            O => \N__4541\,
            I => \N__4538\
        );

    \I__420\ : Span12Mux_v
    port map (
            O => \N__4538\,
            I => \N__4535\
        );

    \I__419\ : Odrv12
    port map (
            O => \N__4535\,
            I => \A_c_2\
        );

    \I__418\ : InMux
    port map (
            O => \N__4532\,
            I => \N__4529\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__4529\,
            I => \N__4526\
        );

    \I__416\ : Span4Mux_v
    port map (
            O => \N__4526\,
            I => \N__4523\
        );

    \I__415\ : Sp12to4
    port map (
            O => \N__4523\,
            I => \N__4520\
        );

    \I__414\ : Span12Mux_h
    port map (
            O => \N__4520\,
            I => \N__4517\
        );

    \I__413\ : Span12Mux_v
    port map (
            O => \N__4517\,
            I => \N__4514\
        );

    \I__412\ : Odrv12
    port map (
            O => \N__4514\,
            I => \A_c_3\
        );

    \I__411\ : InMux
    port map (
            O => \N__4511\,
            I => \N__4508\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__4508\,
            I => \N__4505\
        );

    \I__409\ : Span4Mux_h
    port map (
            O => \N__4505\,
            I => \N__4502\
        );

    \I__408\ : Sp12to4
    port map (
            O => \N__4502\,
            I => \N__4499\
        );

    \I__407\ : Span12Mux_v
    port map (
            O => \N__4499\,
            I => \N__4496\
        );

    \I__406\ : Odrv12
    port map (
            O => \N__4496\,
            I => \A_c_4\
        );

    \I__405\ : IoInMux
    port map (
            O => \N__4493\,
            I => \N__4490\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__4490\,
            I => \N__4487\
        );

    \I__403\ : Odrv12
    port map (
            O => \N__4487\,
            I => \DBRn_c_i_0\
        );

    \I__402\ : IoInMux
    port map (
            O => \N__4484\,
            I => \N__4481\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__4481\,
            I => \N__4478\
        );

    \I__400\ : IoSpan4Mux
    port map (
            O => \N__4478\,
            I => \N__4475\
        );

    \I__399\ : Span4Mux_s3_v
    port map (
            O => \N__4475\,
            I => \N__4472\
        );

    \I__398\ : Odrv4
    port map (
            O => \N__4472\,
            I => \CLK80_PLL_i_i\
        );

    \I__397\ : InMux
    port map (
            O => \N__4469\,
            I => \N__4466\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__4466\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__395\ : InMux
    port map (
            O => \N__4463\,
            I => \bfn_6_7_0_\
        );

    \I__394\ : InMux
    port map (
            O => \N__4460\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__393\ : InMux
    port map (
            O => \N__4457\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__392\ : InMux
    port map (
            O => \N__4454\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__391\ : InMux
    port map (
            O => \N__4451\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__390\ : InMux
    port map (
            O => \N__4448\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__389\ : IoInMux
    port map (
            O => \N__4445\,
            I => \N__4442\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__4442\,
            I => \N__4439\
        );

    \I__387\ : Span4Mux_s0_v
    port map (
            O => \N__4439\,
            I => \N__4436\
        );

    \I__386\ : Span4Mux_v
    port map (
            O => \N__4436\,
            I => \N__4433\
        );

    \I__385\ : Sp12to4
    port map (
            O => \N__4433\,
            I => \N__4430\
        );

    \I__384\ : Span12Mux_h
    port map (
            O => \N__4430\,
            I => \N__4427\
        );

    \I__383\ : Span12Mux_v
    port map (
            O => \N__4427\,
            I => \N__4424\
        );

    \I__382\ : Odrv12
    port map (
            O => \N__4424\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__4670\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            I => \N__4671\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            I => \N__4672\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            I => \N__4669\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            I => \N__4667\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__4668\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\,
            I => \N__4666\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_6_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_7_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_12_0_\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8602\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7997\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4493\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8237\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__8155\,
            in1 => \N__11576\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_2_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11060\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4469\,
            in2 => \_gnd_net_\,
            in3 => \N__4463\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_6_7_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__4673\,
            ce => 'H',
            sr => \N__7553\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4631\,
            in2 => \_gnd_net_\,
            in3 => \N__4460\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__4673\,
            ce => 'H',
            sr => \N__7553\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4604\,
            in2 => \_gnd_net_\,
            in3 => \N__4457\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__4673\,
            ce => 'H',
            sr => \N__7553\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4643\,
            in2 => \_gnd_net_\,
            in3 => \N__4454\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__4673\,
            ce => 'H',
            sr => \N__7553\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4618\,
            in2 => \_gnd_net_\,
            in3 => \N__4451\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__4673\,
            ce => 'H',
            sr => \N__7553\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4580\,
            in2 => \_gnd_net_\,
            in3 => \N__4448\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__4673\,
            ce => 'H',
            sr => \N__7553\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4592\,
            in2 => \_gnd_net_\,
            in3 => \N__4679\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__4673\,
            ce => 'H',
            sr => \N__7553\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5269\,
            in2 => \_gnd_net_\,
            in3 => \N__4676\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4673\,
            ce => 'H',
            sr => \N__7553\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__4642\,
            in1 => \N__4630\,
            in2 => \N__4619\,
            in3 => \N__4603\,
            lcout => \U712_CHIP_RAM.REFRESH5lt7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4591\,
            in2 => \_gnd_net_\,
            in3 => \N__4579\,
            lcout => \U712_CHIP_RAM.REFRESH5lto7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBRn_ibuf_RNIBAB_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4718\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBRn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4568\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11023\,
            ce => \N__5026\,
            sr => \N__11538\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4550\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11029\,
            ce => \N__5022\,
            sr => \N__11535\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4532\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11029\,
            ce => \N__5022\,
            sr => \N__11535\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4511\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11029\,
            ce => \N__5022\,
            sr => \N__11535\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4766\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11029\,
            ce => \N__5022\,
            sr => \N__11535\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4748\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11029\,
            ce => \N__5022\,
            sr => \N__11535\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__6723\,
            in1 => \N__10880\,
            in2 => \_gnd_net_\,
            in3 => \N__5708\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11035\,
            ce => \N__4730\,
            sr => \N__11529\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6140\,
            in1 => \N__5707\,
            in2 => \N__6548\,
            in3 => \N__6644\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11040\,
            ce => \N__5720\,
            sr => \N__11518\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11575\,
            in2 => \_gnd_net_\,
            in3 => \N__4799\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBR_SYNC_0_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4714\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11055\,
            ce => 'H',
            sr => \N__11488\
        );

    \U712_BUFFERS.un1_VBENn_0_a2_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8393\,
            in2 => \_gnd_net_\,
            in3 => \N__9075\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__4958\,
            in1 => \N__5408\,
            in2 => \N__6209\,
            in3 => \N__5213\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11017\,
            ce => \N__5553\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQ8AQ_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6476\,
            in2 => \_gnd_net_\,
            in3 => \N__5801\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_a2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6370\,
            in2 => \_gnd_net_\,
            in3 => \N__7369\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4826\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11024\,
            ce => \N__5027\,
            sr => \N__11530\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI09RS_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__5743\,
            in1 => \N__6429\,
            in2 => \_gnd_net_\,
            in3 => \N__8997\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11573\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5120\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_2_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11574\,
            in2 => \_gnd_net_\,
            in3 => \N__6046\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__6129\,
            in1 => \N__6527\,
            in2 => \N__5339\,
            in3 => \N__6642\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11030\,
            ce => \N__4808\,
            sr => \N__11519\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_1_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6128\,
            in1 => \N__5353\,
            in2 => \N__6643\,
            in3 => \N__6526\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI722C3_1_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__7139\,
            in1 => \N__11334\,
            in2 => \N__4793\,
            in3 => \N__4849\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_165_i_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI30J08_1_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100001101"
        )
    port map (
            in0 => \N__11333\,
            in1 => \N__4862\,
            in2 => \N__4781\,
            in3 => \N__5227\,
            lcout => \U712_CHIP_RAM.N_90_i\,
            ltout => \U712_CHIP_RAM.N_90_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011001010"
        )
    port map (
            in0 => \N__4778\,
            in1 => \N__5114\,
            in2 => \N__4769\,
            in3 => \N__4838\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11036\,
            ce => \N__5555\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000110000"
        )
    port map (
            in0 => \N__7211\,
            in1 => \N__6523\,
            in2 => \N__7145\,
            in3 => \N__7318\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_298_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4868\,
            in3 => \N__5815\,
            lcout => \U712_CHIP_RAM.N_546\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIVFJO_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__5745\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7317\,
            lcout => \U712_CHIP_RAM.N_300\,
            ltout => \U712_CHIP_RAM.N_300_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6525\,
            in1 => \N__7131\,
            in2 => \N__4865\,
            in3 => \N__7212\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_0_0_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIPOTI1_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100011111"
        )
    port map (
            in0 => \N__5744\,
            in1 => \N__6524\,
            in2 => \N__5816\,
            in3 => \N__7319\,
            lcout => \U712_CHIP_RAM.N_313\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7030\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6977\,
            lcout => \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000010001"
        )
    port map (
            in0 => \N__7320\,
            in1 => \N__7213\,
            in2 => \_gnd_net_\,
            in3 => \N__7132\,
            lcout => \U712_CHIP_RAM.N_310\,
            ltout => \U712_CHIP_RAM.N_310_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001010"
        )
    port map (
            in0 => \N__11332\,
            in1 => \N__5231\,
            in2 => \N__4853\,
            in3 => \N__4850\,
            lcout => \U712_CHIP_RAM.N_389\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_5_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11291\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4931\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__4832\,
            in1 => \N__4930\,
            in2 => \_gnd_net_\,
            in3 => \N__5481\,
            lcout => \U712_CHIP_RAM.N_455\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_4_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11290\,
            in2 => \_gnd_net_\,
            in3 => \N__8024\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5080\,
            in1 => \N__5480\,
            in2 => \N__4904\,
            in3 => \N__5102\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4880\,
            in2 => \N__4922\,
            in3 => \N__8329\,
            lcout => \U712_CHIP_RAM.N_419\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5101\,
            in2 => \N__5068\,
            in3 => \N__5069\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4879\,
            in2 => \_gnd_net_\,
            in3 => \N__4919\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4903\,
            in2 => \_gnd_net_\,
            in3 => \N__4916\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5081\,
            in2 => \_gnd_net_\,
            in3 => \N__4913\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_2_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__11251\,
            in1 => \N__4910\,
            in2 => \N__5501\,
            in3 => \N__8333\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11050\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_1_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__8330\,
            in1 => \N__5498\,
            in2 => \N__4889\,
            in3 => \N__11250\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11050\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_0_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__11249\,
            in1 => \N__5108\,
            in2 => \N__5500\,
            in3 => \N__8332\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11050\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_3_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__8331\,
            in1 => \N__5499\,
            in2 => \N__5090\,
            in3 => \N__11252\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11050\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBR_SYNC_RNITKK4_1_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8299\,
            lcout => \DBR_SYNC_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBR_SYNC_1_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5051\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11053\,
            ce => 'H',
            sr => \N__11484\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5045\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11005\,
            ce => \N__5021\,
            sr => \N__11536\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4982\,
            in1 => \N__4964\,
            in2 => \_gnd_net_\,
            in3 => \N__10541\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__5132\,
            in1 => \N__11359\,
            in2 => \_gnd_net_\,
            in3 => \N__5806\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11018\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__5354\,
            in1 => \N__6133\,
            in2 => \_gnd_net_\,
            in3 => \N__6478\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a3_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_178_i_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000111110011"
        )
    port map (
            in0 => \N__9002\,
            in1 => \N__5189\,
            in2 => \N__10775\,
            in3 => \N__5435\,
            lcout => \N_178_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_176_i_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__10689\,
            in1 => \N__5188\,
            in2 => \N__9035\,
            in3 => \N__5453\,
            lcout => \N_176_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5159\,
            in1 => \N__5150\,
            in2 => \_gnd_net_\,
            in3 => \N__10554\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__7373\,
            in1 => \N__8998\,
            in2 => \N__7240\,
            in3 => \N__6477\,
            lcout => \U712_CHIP_RAM.CPU_TACK_8_iv_i_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6085\,
            in1 => \N__7296\,
            in2 => \N__6776\,
            in3 => \N__6518\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOV791_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6515\,
            in1 => \N__5798\,
            in2 => \_gnd_net_\,
            in3 => \N__7111\,
            lcout => \U712_CHIP_RAM.N_370\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_3_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__7110\,
            in1 => \_gnd_net_\,
            in2 => \N__7222\,
            in3 => \N__7294\,
            lcout => \U712_CHIP_RAM.N_464\,
            ltout => \U712_CHIP_RAM.N_464_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIU7TF5_2_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6516\,
            in1 => \N__5335\,
            in2 => \N__5126\,
            in3 => \N__6633\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__5752\,
            in1 => \N__6517\,
            in2 => \N__5123\,
            in3 => \N__6675\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6519\,
            in1 => \N__11358\,
            in2 => \_gnd_net_\,
            in3 => \N__7112\,
            lcout => \U712_CHIP_RAM.N_390\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNIBERN2_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__5799\,
            in1 => \N__6996\,
            in2 => \N__6775\,
            in3 => \N__7295\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_o2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIHSKQ_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5635\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5294\,
            lcout => \U712_CHIP_RAM.N_461\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7316\,
            in2 => \_gnd_net_\,
            in3 => \N__7406\,
            lcout => \U712_CHIP_RAM.N_551\,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5405\,
            in1 => \N__7140\,
            in2 => \_gnd_net_\,
            in3 => \N__5216\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__11031\,
            ce => \N__5554\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6546\,
            in2 => \_gnd_net_\,
            in3 => \N__5204\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5406\,
            in1 => \N__7221\,
            in2 => \_gnd_net_\,
            in3 => \N__5201\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__11031\,
            ce => \N__5554\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5402\,
            in1 => \N__5845\,
            in2 => \_gnd_net_\,
            in3 => \N__5198\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__11031\,
            ce => \N__5554\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5407\,
            in1 => \N__5858\,
            in2 => \_gnd_net_\,
            in3 => \N__5195\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__11031\,
            ce => \N__5554\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5403\,
            in1 => \N__5870\,
            in2 => \_gnd_net_\,
            in3 => \N__5192\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__11031\,
            ce => \N__5554\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__5831\,
            in1 => \N__5404\,
            in2 => \_gnd_net_\,
            in3 => \N__5375\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11031\,
            ce => \N__5554\,
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_188_i_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000111110011"
        )
    port map (
            in0 => \N__5444\,
            in1 => \N__7799\,
            in2 => \N__10771\,
            in3 => \N__9074\,
            lcout => \N_188_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001110"
        )
    port map (
            in0 => \N__5289\,
            in1 => \N__5677\,
            in2 => \N__5628\,
            in3 => \N__5572\,
            lcout => \U712_CHIP_RAM.N_302\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_0_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__5571\,
            in1 => \N__5288\,
            in2 => \N__5696\,
            in3 => \N__5618\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000001000"
        )
    port map (
            in0 => \N__5703\,
            in1 => \N__11352\,
            in2 => \N__7001\,
            in3 => \N__5318\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11037\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5290\,
            in2 => \_gnd_net_\,
            in3 => \N__9073\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_417_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011000100"
        )
    port map (
            in0 => \N__8053\,
            in1 => \N__11351\,
            in2 => \N__5312\,
            in3 => \N__5309\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11037\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010110000"
        )
    port map (
            in0 => \N__5273\,
            in1 => \N__5255\,
            in2 => \N__11360\,
            in3 => \N__5243\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11037\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11349\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5507\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11041\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__10679\,
            in1 => \N__11348\,
            in2 => \_gnd_net_\,
            in3 => \N__10764\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11041\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100000000"
        )
    port map (
            in0 => \N__5491\,
            in1 => \N__5459\,
            in2 => \N__8344\,
            in3 => \N__11350\,
            lcout => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11041\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UUBE_i_o2_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100011111"
        )
    port map (
            in0 => \N__9612\,
            in1 => \N__9766\,
            in2 => \N__9528\,
            in3 => \N__9702\,
            lcout => \U712_BYTE_ENABLE.N_326\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LLBE_i_o2_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010101111"
        )
    port map (
            in0 => \N__9765\,
            in1 => \N__9611\,
            in2 => \N__9706\,
            in3 => \N__9515\,
            lcout => \U712_BYTE_ENABLE.N_323\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UMBE_i_o2_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101101110101"
        )
    port map (
            in0 => \N__9475\,
            in1 => \N__9756\,
            in2 => \N__9623\,
            in3 => \N__9684\,
            lcout => \U712_BYTE_ENABLE.N_324\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5426\,
            in1 => \N__6035\,
            in2 => \_gnd_net_\,
            in3 => \N__10542\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7236\,
            in1 => \N__5805\,
            in2 => \N__6542\,
            in3 => \N__7368\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__6194\,
            in1 => \N__6536\,
            in2 => \N__7241\,
            in3 => \N__7374\,
            lcout => \U712_CHIP_RAM.N_384\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIR80N2_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__11357\,
            in1 => \N__5800\,
            in2 => \_gnd_net_\,
            in3 => \N__6759\,
            lcout => \U712_CHIP_RAM.N_463\,
            ltout => \U712_CHIP_RAM.N_463_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIONRK3_1_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6535\,
            in2 => \N__5642\,
            in3 => \N__7146\,
            lcout => \U712_CHIP_RAM.N_550\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__6131\,
            in1 => \N__5698\,
            in2 => \N__5639\,
            in3 => \N__6195\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_385_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__6161\,
            in1 => \_gnd_net_\,
            in2 => \N__5600\,
            in3 => \N__6250\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110100000001"
        )
    port map (
            in0 => \N__5597\,
            in1 => \N__6818\,
            in2 => \N__5591\,
            in3 => \N__10548\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11010\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNICG3P2_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__5588\,
            in1 => \N__6130\,
            in2 => \N__5582\,
            in3 => \N__6534\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERlde_0_a3_0_0_a2_0\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTERlde_0_a3_0_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5697\,
            in2 => \N__5558\,
            in3 => \N__6193\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI36AQC_2_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__6538\,
            in1 => \N__6191\,
            in2 => \N__5894\,
            in3 => \N__6132\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNINN3QI_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__6192\,
            in1 => \N__5522\,
            in2 => \N__5510\,
            in3 => \N__5699\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11338\,
            in2 => \_gnd_net_\,
            in3 => \N__6760\,
            lcout => \U712_CHIP_RAM.N_533\,
            ltout => \U712_CHIP_RAM.N_533_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_3_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7363\,
            in1 => \N__7214\,
            in2 => \N__5906\,
            in3 => \N__5903\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_391_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIEVI78_3_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6190\,
            in2 => \N__5897\,
            in3 => \N__6084\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__6761\,
            in1 => \N__6539\,
            in2 => \N__7375\,
            in3 => \N__6086\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11019\,
            ce => \N__6656\,
            sr => \N__11505\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5869\,
            in1 => \N__5857\,
            in2 => \N__5846\,
            in3 => \N__5830\,
            lcout => \U712_CHIP_RAM.N_295\,
            ltout => \U712_CHIP_RAM.N_295_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5819\,
            in3 => \N__5797\,
            lcout => \U712_CHIP_RAM.N_458\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNILJ788_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__6978\,
            in1 => \N__6696\,
            in2 => \N__7362\,
            in3 => \N__7407\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIMAOKC_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__6531\,
            in1 => \N__6676\,
            in2 => \N__5759\,
            in3 => \N__5756\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5723\,
            in3 => \N__11571\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5678\,
            in1 => \N__6125\,
            in2 => \N__6547\,
            in3 => \N__6623\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIF4EE6_2_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100000"
        )
    port map (
            in0 => \N__6126\,
            in1 => \N__6533\,
            in2 => \N__6251\,
            in3 => \N__6157\,
            lcout => \U712_CHIP_RAM.N_441\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6532\,
            in1 => \N__6127\,
            in2 => \_gnd_net_\,
            in3 => \N__6768\,
            lcout => \U712_CHIP_RAM.DBENn_8_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__7201\,
            in1 => \N__7109\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_465\,
            ltout => \U712_CHIP_RAM.N_465_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_3_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6068\,
            in3 => \N__6622\,
            lcout => \U712_CHIP_RAM.N_469\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__6065\,
            in1 => \N__6034\,
            in2 => \N__11837\,
            in3 => \N__6050\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11032\,
            ce => 'H',
            sr => \N__11492\
        );

    \U712_CHIP_RAM.DBENn_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100111011101110"
        )
    port map (
            in0 => \N__6020\,
            in1 => \N__7022\,
            in2 => \N__6014\,
            in3 => \N__10178\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11032\,
            ce => 'H',
            sr => \N__11492\
        );

    \U712_CHIP_RAM.DBDIR_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__6731\,
            in1 => \N__5986\,
            in2 => \_gnd_net_\,
            in3 => \N__6697\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11032\,
            ce => 'H',
            sr => \N__11492\
        );

    \pll_RNI8MQ3_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__7718\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.N_167_i_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__10807\,
            in1 => \N__10667\,
            in2 => \_gnd_net_\,
            in3 => \N__10762\,
            lcout => \N_167_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6337\,
            in1 => \N__6302\,
            in2 => \_gnd_net_\,
            in3 => \N__10586\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__10587\,
            in1 => \N__9084\,
            in2 => \N__6290\,
            in3 => \N__10139\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__6994\,
            in1 => \N__6268\,
            in2 => \N__7376\,
            in3 => \N__7385\,
            lcout => \LATCH_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11002\,
            ce => 'H',
            sr => \N__11511\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__10502\,
            in1 => \N__9163\,
            in2 => \N__12174\,
            in3 => \N__10411\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__6257\,
            in1 => \N__6249\,
            in2 => \N__6569\,
            in3 => \N__6220\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_296_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6819\,
            in2 => \N__6230\,
            in3 => \N__9164\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11006\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000011"
        )
    port map (
            in0 => \N__12173\,
            in1 => \N__6797\,
            in2 => \N__6227\,
            in3 => \N__6821\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11011\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6541\,
            in1 => \N__7148\,
            in2 => \N__6205\,
            in3 => \N__7367\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_442_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001011"
        )
    port map (
            in0 => \N__10421\,
            in1 => \N__6820\,
            in2 => \N__6800\,
            in3 => \N__6796\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11011\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6788\,
            in2 => \_gnd_net_\,
            in3 => \N__6767\,
            lcout => \U712_CHIP_RAM.N_428\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011000000"
        )
    port map (
            in0 => \N__6727\,
            in1 => \N__10788\,
            in2 => \N__11356\,
            in3 => \N__6698\,
            lcout => \DMA_WRITE_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11011\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__6540\,
            in1 => \N__6634\,
            in2 => \N__7052\,
            in3 => \N__6680\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6659\,
            in3 => \N__11570\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__7051\,
            in1 => \N__6635\,
            in2 => \N__6386\,
            in3 => \N__6593\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011111010"
        )
    port map (
            in0 => \N__7754\,
            in1 => \N__6581\,
            in2 => \N__6572\,
            in3 => \N__7144\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11020\,
            ce => 'H',
            sr => \N__11493\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI1NGC4_2_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__6562\,
            in1 => \N__6537\,
            in2 => \_gnd_net_\,
            in3 => \N__7408\,
            lcout => \U712_CHIP_RAM.N_438\,
            ltout => \U712_CHIP_RAM.N_438_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__7409\,
            in1 => \N__6997\,
            in2 => \N__7388\,
            in3 => \N__7338\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIREK92_3_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__7334\,
            in1 => \N__7226\,
            in2 => \N__7147\,
            in3 => \N__7064\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__7844\,
            in1 => \N__7860\,
            in2 => \_gnd_net_\,
            in3 => \N__7753\,
            lcout => \U712_CYCLE_TERM.N_321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7023\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6995\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011111111"
        )
    port map (
            in0 => \N__7877\,
            in1 => \N__6884\,
            in2 => \_gnd_net_\,
            in3 => \N__6935\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11033\,
            ce => 'H',
            sr => \N__11489\
        );

    \U712_BYTE_ENABLE.LMBE_i_o2_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000101111"
        )
    port map (
            in0 => \N__9767\,
            in1 => \N__9624\,
            in2 => \N__9707\,
            in3 => \N__9519\,
            lcout => \U712_BYTE_ENABLE.N_325\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__9368\,
            in1 => \N__11921\,
            in2 => \N__9329\,
            in3 => \N__6866\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11001\,
            ce => \N__9244\,
            sr => \N__11510\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10599\,
            in1 => \N__6845\,
            in2 => \_gnd_net_\,
            in3 => \N__6833\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9083\,
            in1 => \N__10600\,
            in2 => \N__6824\,
            in3 => \N__8618\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7583\,
            in1 => \N__7568\,
            in2 => \_gnd_net_\,
            in3 => \N__10598\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__10549\,
            in1 => \N__12166\,
            in2 => \N__10422\,
            in3 => \N__7546\,
            lcout => \U712_CHIP_RAM.un1_CMA25_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7528\,
            in1 => \N__7505\,
            in2 => \_gnd_net_\,
            in3 => \N__10550\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__10551\,
            in1 => \N__9081\,
            in2 => \N__7496\,
            in3 => \N__8702\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7474\,
            in1 => \N__7454\,
            in2 => \_gnd_net_\,
            in3 => \N__10552\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10415\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9165\,
            lcout => \U712_CHIP_RAM.N_305\,
            ltout => \U712_CHIP_RAM.N_305_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000001111"
        )
    port map (
            in0 => \N__9082\,
            in1 => \N__10267\,
            in2 => \N__7445\,
            in3 => \N__10553\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9079\,
            in1 => \N__7442\,
            in2 => \_gnd_net_\,
            in3 => \N__8720\,
            lcout => \U712_CHIP_RAM.N_346\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7421\,
            in1 => \N__9080\,
            in2 => \_gnd_net_\,
            in3 => \N__8681\,
            lcout => \U712_CHIP_RAM.N_352\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_186_i_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__10691\,
            in1 => \N__7798\,
            in2 => \N__7784\,
            in3 => \N__9085\,
            lcout => \N_186_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7845\,
            in2 => \_gnd_net_\,
            in3 => \N__7751\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__7709\,
            in1 => \N__11245\,
            in2 => \_gnd_net_\,
            in3 => \N__7908\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100010101"
        )
    port map (
            in0 => \N__7907\,
            in1 => \N__7846\,
            in2 => \N__7865\,
            in3 => \N__7752\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_450_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__7710\,
            in1 => \N__7864\,
            in2 => \N__7733\,
            in3 => \N__11244\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__11246\,
            in1 => \_gnd_net_\,
            in2 => \N__7730\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7665\,
            in2 => \_gnd_net_\,
            in3 => \N__7726\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__11247\,
            in1 => \_gnd_net_\,
            in2 => \N__7670\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111000100"
        )
    port map (
            in0 => \N__7910\,
            in1 => \N__7601\,
            in2 => \N__7714\,
            in3 => \N__7669\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11022\,
            ce => 'H',
            sr => \N__11483\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010101000000"
        )
    port map (
            in0 => \N__7909\,
            in1 => \N__7892\,
            in2 => \N__7886\,
            in3 => \N__7876\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11022\,
            ce => 'H',
            sr => \N__11483\
        );

    \U712_REG_SM.REG_TACK_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__8015\,
            in1 => \N__7847\,
            in2 => \N__8354\,
            in3 => \N__7826\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11022\,
            ce => 'H',
            sr => \N__11483\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__9983\,
            in1 => \N__8360\,
            in2 => \_gnd_net_\,
            in3 => \N__8915\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11022\,
            ce => 'H',
            sr => \N__11483\
        );

    \U712_REG_SM.STATE_COUNT_5_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11194\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7805\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11025\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111110"
        )
    port map (
            in0 => \N__8889\,
            in1 => \N__7819\,
            in2 => \N__9979\,
            in3 => \N__8913\,
            lcout => \U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_7_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11196\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7811\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11025\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_6_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11195\,
            in2 => \_gnd_net_\,
            in3 => \N__7820\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11025\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11193\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8014\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11025\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIH4AH_1_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__10030\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8334\,
            lcout => \U712_REG_SM.N_320\,
            ltout => \U712_REG_SM.N_320_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_0_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__8250\,
            in1 => \N__9978\,
            in2 => \N__8000\,
            in3 => \N__12304\,
            lcout => \U712_REG_SM.N_409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11248\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__9119\,
            in1 => \N__7985\,
            in2 => \N__10370\,
            in3 => \N__10605\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__10601\,
            in1 => \N__9120\,
            in2 => \N__7979\,
            in3 => \N__10127\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11572\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7964\,
            lcout => \U712_CHIP_RAM.un1_CMA25_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__7958\,
            in1 => \N__9121\,
            in2 => \N__10612\,
            in3 => \N__8126\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9115\,
            in1 => \N__7949\,
            in2 => \N__10597\,
            in3 => \N__8690\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7916\,
            in2 => \N__7943\,
            in3 => \N__7940\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11007\,
            ce => \N__9250\,
            sr => \N__11506\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111010101"
        )
    port map (
            in0 => \N__10562\,
            in1 => \N__9355\,
            in2 => \N__9123\,
            in3 => \N__10268\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__8189\,
            in1 => \N__9359\,
            in2 => \N__10616\,
            in3 => \N__8183\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11012\,
            ce => \N__9240\,
            sr => \N__11499\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__11831\,
            in1 => \N__8156\,
            in2 => \N__11906\,
            in3 => \N__8125\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\,
            ce => 'H',
            sr => \N__11494\
        );

    \U712_BUFFERS.N_169_i_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101010"
        )
    port map (
            in0 => \N__9122\,
            in1 => \N__10690\,
            in2 => \N__10763\,
            in3 => \N__8386\,
            lcout => \N_169_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8935\,
            in2 => \_gnd_net_\,
            in3 => \N__8858\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_397_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100010"
        )
    port map (
            in0 => \N__11301\,
            in1 => \N__8087\,
            in2 => \N__8063\,
            in3 => \N__8060\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_3_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11300\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10166\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIJUGT_3_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000001000"
        )
    port map (
            in0 => \N__10038\,
            in1 => \N__8275\,
            in2 => \N__12324\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.N_548\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12297\,
            in2 => \_gnd_net_\,
            in3 => \N__10037\,
            lcout => \U712_REG_SM.N_319\,
            ltout => \U712_REG_SM.N_319_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_1_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__9883\,
            in1 => \N__8378\,
            in2 => \N__8003\,
            in3 => \N__9963\,
            lcout => OPEN,
            ltout => \U712_REG_SM.REG_CYCLE_5_iv_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011100010"
        )
    port map (
            in0 => \N__8379\,
            in1 => \N__11192\,
            in2 => \N__8402\,
            in3 => \N__8399\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11038\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100000000"
        )
    port map (
            in0 => \N__8861\,
            in1 => \N__10039\,
            in2 => \N__12325\,
            in3 => \N__8888\,
            lcout => \U712_REG_SM.STATE_COUNTsr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9882\,
            in1 => \N__8274\,
            in2 => \_gnd_net_\,
            in3 => \N__9962\,
            lcout => \U712_REG_SM.N_328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__10031\,
            in1 => \N__8276\,
            in2 => \N__8345\,
            in3 => \N__8251\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_412_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001010"
        )
    port map (
            in0 => \N__11317\,
            in1 => \N__12307\,
            in2 => \N__8279\,
            in3 => \N__10033\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11042\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111000101"
        )
    port map (
            in0 => \N__8252\,
            in1 => \N__12305\,
            in2 => \N__10082\,
            in3 => \N__10032\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_360_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000000100"
        )
    port map (
            in0 => \N__12306\,
            in1 => \N__11316\,
            in2 => \N__8261\,
            in3 => \N__8258\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11042\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_0_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8224\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11045\,
            ce => 'H',
            sr => \N__11479\
        );

    \U712_REG_SM.C3_SYNC_1_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8195\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11045\,
            ce => 'H',
            sr => \N__11479\
        );

    \U712_REG_SM.C1_SYNC_1_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8567\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11049\,
            ce => 'H',
            sr => \N__11478\
        );

    \U712_REG_SM.C1_SYNC_0_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8603\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11051\,
            ce => 'H',
            sr => \N__11477\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__9390\,
            in1 => \N__9311\,
            in2 => \N__10115\,
            in3 => \N__8561\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11003\,
            ce => \N__9249\,
            sr => \N__11531\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_14_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__12184\,
            in1 => \N__9391\,
            in2 => \_gnd_net_\,
            in3 => \N__10610\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11003\,
            ce => \N__9249\,
            sr => \N__11531\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__8711\,
            in1 => \N__9392\,
            in2 => \N__9326\,
            in3 => \N__8513\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11003\,
            ce => \N__9249\,
            sr => \N__11531\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__10151\,
            in1 => \N__9388\,
            in2 => \N__9328\,
            in3 => \N__8486\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11008\,
            ce => \N__9245\,
            sr => \N__11520\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__9386\,
            in1 => \N__8729\,
            in2 => \N__9325\,
            in3 => \N__8456\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11008\,
            ce => \N__9245\,
            sr => \N__11520\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__12026\,
            in1 => \N__9387\,
            in2 => \N__9327\,
            in3 => \N__8426\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11008\,
            ce => \N__9245\,
            sr => \N__11520\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__9140\,
            in1 => \N__8771\,
            in2 => \N__9125\,
            in3 => \N__11660\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11013\,
            ce => \N__9251\,
            sr => \N__11512\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10313\,
            in1 => \N__11757\,
            in2 => \_gnd_net_\,
            in3 => \N__10353\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11648\,
            ce => \N__11612\,
            sr => \N__11507\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10354\,
            in1 => \N__11759\,
            in2 => \_gnd_net_\,
            in3 => \N__8668\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11648\,
            ce => \N__11612\,
            sr => \N__11507\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8669\,
            in1 => \N__11758\,
            in2 => \_gnd_net_\,
            in3 => \N__12122\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11648\,
            ce => \N__11612\,
            sr => \N__11507\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11760\,
            in1 => \N__12005\,
            in2 => \_gnd_net_\,
            in3 => \N__10249\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__11610\,
            sr => \N__11500\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12006\,
            in1 => \N__11761\,
            in2 => \_gnd_net_\,
            in3 => \N__11965\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__11610\,
            sr => \N__11500\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8666\,
            in1 => \N__11827\,
            in2 => \_gnd_net_\,
            in3 => \N__12121\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__11610\,
            sr => \N__11500\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11812\,
            in1 => \N__8667\,
            in2 => \_gnd_net_\,
            in3 => \N__10352\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__11609\,
            sr => \N__11495\
        );

    \U712_REG_SM.REGENn_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100011011000100"
        )
    port map (
            in0 => \N__8792\,
            in1 => \N__8811\,
            in2 => \N__12332\,
            in3 => \N__8896\,
            lcout => \BLSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11039\,
            ce => 'H',
            sr => \N__11490\
        );

    \U712_REG_SM.START_RST_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__10078\,
            in1 => \N__8936\,
            in2 => \_gnd_net_\,
            in3 => \N__10099\,
            lcout => \U712_REG_SM.START_RSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11039\,
            ce => 'H',
            sr => \N__11490\
        );

    \U712_REG_SM.STATE_COUNT_8_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__8924\,
            in1 => \N__11265\,
            in2 => \N__9977\,
            in3 => \N__8914\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11043\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8859\,
            in1 => \N__10041\,
            in2 => \N__12329\,
            in3 => \N__8897\,
            lcout => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10042\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12314\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_318_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__11264\,
            in1 => \N__10100\,
            in2 => \N__8864\,
            in3 => \N__10079\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11043\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_RNO_0_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001000100"
        )
    port map (
            in0 => \N__8860\,
            in1 => \N__10040\,
            in2 => \N__10081\,
            in3 => \N__8810\,
            lcout => \U712_REG_SM.REGENn_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDSn_RNO_0_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001000"
        )
    port map (
            in0 => \N__9614\,
            in1 => \N__9532\,
            in2 => \N__10888\,
            in3 => \N__9683\,
            lcout => \U712_REG_SM.N_400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_RNO_0_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__10870\,
            in1 => \N__9613\,
            in2 => \N__9533\,
            in3 => \N__9682\,
            lcout => \U712_REG_SM.N_398\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_326_i_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001001000"
        )
    port map (
            in0 => \N__9681\,
            in1 => \N__9755\,
            in2 => \N__9521\,
            in3 => \N__9622\,
            lcout => \N_326_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_325_i_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101000010010"
        )
    port map (
            in0 => \N__9680\,
            in1 => \N__9754\,
            in2 => \N__9520\,
            in3 => \N__9621\,
            lcout => \N_325_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_323_i_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101000100"
        )
    port map (
            in0 => \N__9752\,
            in1 => \N__9678\,
            in2 => \N__9625\,
            in3 => \N__9502\,
            lcout => \N_323_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_324_i_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001110001000"
        )
    port map (
            in0 => \N__9753\,
            in1 => \N__9679\,
            in2 => \N__9626\,
            in3 => \N__9503\,
            lcout => \N_324_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WEn_LC_15_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9179\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11004\,
            ce => 'H',
            sr => \N__11539\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_15_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9108\,
            in2 => \_gnd_net_\,
            in3 => \N__10609\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__9389\,
            in1 => \N__8945\,
            in2 => \N__9324\,
            in3 => \N__8951\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11014\,
            ce => \N__9233\,
            sr => \N__11532\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__10429\,
            in1 => \N__10560\,
            in2 => \_gnd_net_\,
            in3 => \N__9178\,
            lcout => \U712_CHIP_RAM.CMA_5_i_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__9134\,
            in1 => \N__10561\,
            in2 => \N__9124\,
            in3 => \N__10274\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11799\,
            in1 => \N__10312\,
            in2 => \_gnd_net_\,
            in3 => \N__11969\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11647\,
            ce => \N__11615\,
            sr => \N__11513\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12071\,
            in1 => \N__11800\,
            in2 => \_gnd_net_\,
            in3 => \N__11902\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11647\,
            ce => \N__11615\,
            sr => \N__11513\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11823\,
            in1 => \N__10305\,
            in2 => \_gnd_net_\,
            in3 => \N__11964\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__11613\,
            sr => \N__11508\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__11895\,
            in1 => \_gnd_net_\,
            in2 => \N__11836\,
            in3 => \N__12070\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__11613\,
            sr => \N__11508\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10202\,
            in1 => \N__11811\,
            in2 => \_gnd_net_\,
            in3 => \N__10239\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11643\,
            ce => \N__11611\,
            sr => \N__11501\
        );

    \U712_REG_SM.WRITE_CYCLE_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__10889\,
            in1 => \N__9878\,
            in2 => \_gnd_net_\,
            in3 => \N__10098\,
            lcout => \U712_REG_SM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11046\,
            ce => 'H',
            sr => \N__11491\
        );

    \U712_REG_SM.STATE_COUNT_RNI3HF31_1_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__10080\,
            in1 => \N__12320\,
            in2 => \N__10043\,
            in3 => \N__9967\,
            lcout => \U712_REG_SM.N_152\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDSn_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__12318\,
            in1 => \N__9920\,
            in2 => \N__9901\,
            in3 => \N__12357\,
            lcout => \UDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11052\,
            ce => 'H',
            sr => \N__11481\
        );

    \U712_REG_SM.PRnW_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101111111010000"
        )
    port map (
            in0 => \N__9884\,
            in1 => \N__12319\,
            in2 => \N__12359\,
            in3 => \N__9844\,
            lcout => \PRnW_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11052\,
            ce => 'H',
            sr => \N__11481\
        );

    \U712_REG_SM.LDSn_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__9833\,
            in1 => \N__12358\,
            in2 => \N__9817\,
            in3 => \N__12330\,
            lcout => \LDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11054\,
            ce => 'H',
            sr => \N__11480\
        );

    \U712_CHIP_RAM.CASn_LC_16_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10611\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11009\,
            ce => 'H',
            sr => \N__11544\
        );

    \U712_CHIP_RAM.RASn_LC_16_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10433\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11015\,
            ce => 'H',
            sr => \N__11540\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12069\,
            in1 => \N__11835\,
            in2 => \_gnd_net_\,
            in3 => \N__12119\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__11619\,
            sr => \N__11533\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11798\,
            in1 => \N__10355\,
            in2 => \_gnd_net_\,
            in3 => \N__10304\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            ce => \N__11617\,
            sr => \N__11521\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12013\,
            in1 => \N__11819\,
            in2 => \_gnd_net_\,
            in3 => \N__10250\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11644\,
            ce => \N__11616\,
            sr => \N__11514\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10238\,
            in1 => \N__11801\,
            in2 => \_gnd_net_\,
            in3 => \N__10201\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__11614\,
            sr => \N__11509\
        );

    \U712_CHIP_RAM.RAS_SYNC_2_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11243\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10157\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11047\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_1_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11242\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11066\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11047\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_ess_RNO_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11569\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12350\,
            lcout => \U712_REG_SM.N_152_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_ess_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12331\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11056\,
            ce => \N__12197\,
            sr => \N__11482\
        );

    \U712_CHIP_RAM.CRCSn_LC_17_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12185\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11021\,
            ce => 'H',
            sr => \N__11545\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12120\,
            in1 => \N__11830\,
            in2 => \_gnd_net_\,
            in3 => \N__12068\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11646\,
            ce => \N__11621\,
            sr => \N__11537\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12014\,
            in1 => \N__11829\,
            in2 => \_gnd_net_\,
            in3 => \N__11947\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11645\,
            ce => \N__11620\,
            sr => \N__11534\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11885\,
            in1 => \N__11828\,
            in2 => \_gnd_net_\,
            in3 => \N__11089\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11642\,
            ce => \N__11618\,
            sr => \N__11522\
        );

    \U712_CHIP_RAM.RAS_SYNC_0_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__11263\,
            in1 => \N__11105\,
            in2 => \_gnd_net_\,
            in3 => \N__11093\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11048\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_i_m2_LC_24_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001100110011"
        )
    port map (
            in0 => \N__10887\,
            in1 => \N__10808\,
            in2 => \N__10727\,
            in3 => \N__10666\,
            lcout => \N_362\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

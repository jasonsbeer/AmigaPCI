-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     May 31 2025 15:09:50

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U111_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U111_TOP
entity U111_TOP is
port (
    D_UU_AMIGA : inout std_logic_vector(7 downto 0);
    D_LL_AMIGA : inout std_logic_vector(7 downto 0);
    D_UM_AMIGA : inout std_logic_vector(7 downto 0);
    D_LM_AMIGA : inout std_logic_vector(7 downto 0);
    D_UU_040 : inout std_logic_vector(7 downto 0);
    D_LM_040 : inout std_logic_vector(7 downto 0);
    D_UM_040 : inout std_logic_vector(7 downto 0);
    D_LL_040 : inout std_logic_vector(7 downto 0);
    A_AMIGA : out std_logic_vector(1 downto 0);
    A_040 : in std_logic_vector(1 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    TEAn : in std_logic;
    TSn : out std_logic;
    RESETn : in std_logic;
    CLKRAMA : out std_logic;
    PORTSIZE : in std_logic;
    TEA_CPUn : out std_logic;
    LBENn : in std_logic;
    CLK40B : out std_logic;
    TBI_CPUn : out std_logic;
    TAn : inout std_logic;
    CPUBGn : out std_logic;
    BUFENn : out std_logic;
    RnW : in std_logic;
    CLK80_CPU : out std_logic;
    BUFDIR : out std_logic;
    TCI_CPUn : out std_logic;
    TS_CPUn : in std_logic;
    CLKRAMB : out std_logic;
    CLK40A : out std_logic;
    TCIn : in std_logic;
    TBIn : in std_logic;
    DMAn : out std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    TACKn : inout std_logic;
    BGn : in std_logic);
end U111_TOP;

-- Architecture of U111_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U111_TOP is

signal \N__8833\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7827\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7260\ : std_logic;
signal \N__7257\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3959\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3853\ : std_logic;
signal \N__3850\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3809\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3622\ : std_logic;
signal \N__3619\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3587\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3548\ : std_logic;
signal \N__3545\ : std_logic;
signal \N__3542\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3520\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3482\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3476\ : std_logic;
signal \N__3473\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3457\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3442\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3404\ : std_logic;
signal \N__3401\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3392\ : std_logic;
signal \N__3389\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3383\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3353\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3339\ : std_logic;
signal \N__3336\ : std_logic;
signal \N__3333\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3265\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3253\ : std_logic;
signal \N__3250\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3209\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3176\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3140\ : std_logic;
signal \N__3137\ : std_logic;
signal \N__3134\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3121\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3115\ : std_logic;
signal \N__3112\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3067\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3056\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2987\ : std_logic;
signal \N__2984\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2875\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2863\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2768\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2747\ : std_logic;
signal \N__2744\ : std_logic;
signal \N__2741\ : std_logic;
signal \N__2738\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2705\ : std_logic;
signal \N__2702\ : std_logic;
signal \N__2699\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2672\ : std_logic;
signal \N__2669\ : std_logic;
signal \N__2666\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2650\ : std_logic;
signal \N__2647\ : std_logic;
signal \N__2644\ : std_logic;
signal \N__2641\ : std_logic;
signal \N__2638\ : std_logic;
signal \N__2635\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2612\ : std_logic;
signal \N__2609\ : std_logic;
signal \N__2606\ : std_logic;
signal \N__2603\ : std_logic;
signal \N__2600\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2579\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2546\ : std_logic;
signal \N__2543\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2507\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2501\ : std_logic;
signal \N__2498\ : std_logic;
signal \N__2495\ : std_logic;
signal \TCIn_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \TAn_in\ : std_logic;
signal \A_040_c_0\ : std_logic;
signal \A_AMIGA_c_0\ : std_logic;
signal \U111_CYCLE_SM_A_AMIGA_0_i_1\ : std_logic;
signal \D_LL_AMIGA_in_0\ : std_logic;
signal \un1_D_LL_AMIGA_0\ : std_logic;
signal \D_LL_AMIGA_in_1\ : std_logic;
signal \un1_D_LL_AMIGA_1\ : std_logic;
signal \D_LL_AMIGA_in_3\ : std_logic;
signal \un1_D_LL_AMIGA_3\ : std_logic;
signal \D_UM_040_in_6\ : std_logic;
signal \D_LL_040_in_6\ : std_logic;
signal \un1_D_UM_040_6\ : std_logic;
signal \LBENn_c_i\ : std_logic;
signal \D_LM_AMIGA_in_4\ : std_logic;
signal \un1_D_LM_AMIGA_4\ : std_logic;
signal \D_LM_AMIGA_in_5\ : std_logic;
signal \un1_D_LM_AMIGA_5\ : std_logic;
signal \D_LM_AMIGA_in_7\ : std_logic;
signal \un1_D_LM_AMIGA_7\ : std_logic;
signal \D_LM_AMIGA_in_6\ : std_logic;
signal \un1_D_LM_AMIGA_6\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \D_LM_040_in_7\ : std_logic;
signal \D_UU_040_in_7\ : std_logic;
signal \un1_D_UU_040_7\ : std_logic;
signal \D_LM_AMIGA_in_3\ : std_logic;
signal \un1_D_LM_AMIGA_3\ : std_logic;
signal \D_UM_040_in_0\ : std_logic;
signal \D_LL_040_in_0\ : std_logic;
signal \un1_D_UM_040_0\ : std_logic;
signal \D_UU_040_in_1\ : std_logic;
signal \D_LM_040_in_1\ : std_logic;
signal \un1_D_UU_040_1\ : std_logic;
signal \D_UU_040_in_4\ : std_logic;
signal \D_LM_040_in_4\ : std_logic;
signal \un1_D_UU_040_4\ : std_logic;
signal \D_UU_040_in_0\ : std_logic;
signal \D_LM_040_in_0\ : std_logic;
signal \un1_D_UU_040_0\ : std_logic;
signal \un1_D_UM_AMIGA_0\ : std_logic;
signal \D_LM_AMIGA_in_1\ : std_logic;
signal \un1_D_LM_AMIGA_1\ : std_logic;
signal \D_UM_AMIGA_in_0\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\ : std_logic;
signal \un1_D_UM_AMIGA_1\ : std_logic;
signal \D_UM_AMIGA_in_1\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\ : std_logic;
signal \un1_D_UU_AMIGA_1\ : std_logic;
signal \D_UU_AMIGA_in_1\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\ : std_logic;
signal \D_UU_040_in_2\ : std_logic;
signal \D_LM_040_in_2\ : std_logic;
signal \un1_D_UU_040_2\ : std_logic;
signal \D_LL_040_in_5\ : std_logic;
signal \D_UM_040_in_5\ : std_logic;
signal \un1_D_UM_040_5\ : std_logic;
signal \LBENn_c_i_0\ : std_logic;
signal \D_LL_AMIGA_in_6\ : std_logic;
signal \un1_D_LL_AMIGA_6\ : std_logic;
signal \D_LL_AMIGA_in_5\ : std_logic;
signal \un1_D_LL_AMIGA_5\ : std_logic;
signal \A_040_c_1\ : std_logic;
signal \D_LL_AMIGA_in_7\ : std_logic;
signal \un1_D_LL_AMIGA_7\ : std_logic;
signal \D_LM_AMIGA_in_0\ : std_logic;
signal \un1_D_LM_AMIGA_0\ : std_logic;
signal \TSn_c\ : std_logic;
signal \INVU111_CYCLE_SM.TSnC_net\ : std_logic;
signal \D_UU_AMIGA_1_i\ : std_logic;
signal \U111_CYCLE_SM.TS_ENZ0\ : std_logic;
signal \U111_CYCLE_SM.FLIP_WORD_2\ : std_logic;
signal \D_UM_040_in_2\ : std_logic;
signal \D_LL_040_in_2\ : std_logic;
signal \un1_D_UM_040_2\ : std_logic;
signal \GB_BUFFER_CLK40_THRU_CO\ : std_logic;
signal \U111_CYCLE_SM.PORT_MISMATCH_2\ : std_logic;
signal \U111_CYCLE_SM.N_123_0_cascade_\ : std_logic;
signal \U111_CYCLE_SM.N_121_0\ : std_logic;
signal \U111_CYCLE_SM.un1_CYCLE_STATE_0\ : std_logic;
signal \D_UU_040_1_i\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81_cascade_\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\ : std_logic;
signal \D_UU_AMIGA_in_6\ : std_logic;
signal \un1_D_UU_AMIGA_6\ : std_logic;
signal \D_UU_AMIGA_in_0\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\ : std_logic;
signal \un1_D_UU_AMIGA_0\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\ : std_logic;
signal \un1_D_UU_AMIGA_2\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\ : std_logic;
signal \D_UM_AMIGA_in_5\ : std_logic;
signal \un1_D_UM_AMIGA_5\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\ : std_logic;
signal \D_UU_AMIGA_in_7\ : std_logic;
signal \un1_D_UU_AMIGA_7\ : std_logic;
signal \D_LL_AMIGA_in_2\ : std_logic;
signal \un1_D_LL_AMIGA_2\ : std_logic;
signal \D_LL_AMIGA_in_4\ : std_logic;
signal \un1_D_LL_AMIGA_4\ : std_logic;
signal \U111_CYCLE_SM.A2_ENZ0\ : std_logic;
signal \U111_CYCLE_SM.N_148\ : std_logic;
signal \U111_CYCLE_SM.N_148_cascade_\ : std_logic;
signal \U111_CYCLE_SM.TS_EN_6\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_srsts_i_o2_0_5_cascade_\ : std_logic;
signal \LBENn_c\ : std_logic;
signal \U111_CYCLE_SM.TA_DISZ0\ : std_logic;
signal \TAn_1_i\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\ : std_logic;
signal \U111_CYCLE_SM.N_135_cascade_\ : std_logic;
signal \U111_CYCLE_SM.N_128_0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_srsts_0_1_0_cascade_\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\ : std_logic;
signal \TEAn_c\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_srsts_i_1_2_cascade_\ : std_logic;
signal \CLK80\ : std_logic;
signal \GB_BUFFER_CLK80_THRU_CO\ : std_logic;
signal \D_LM_AMIGA_in_2\ : std_logic;
signal \D_UU_AMIGA_in_2\ : std_logic;
signal \un1_D_LM_AMIGA_2\ : std_logic;
signal \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81\ : std_logic;
signal \D_UM_AMIGA_in_4\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\ : std_logic;
signal \un1_D_UM_AMIGA_4\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\ : std_logic;
signal \D_UU_AMIGA_in_3\ : std_logic;
signal \un1_D_UU_AMIGA_3\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\ : std_logic;
signal \D_UM_AMIGA_in_3\ : std_logic;
signal \un1_D_UM_AMIGA_3\ : std_logic;
signal \D_UM_040_in_3\ : std_logic;
signal \D_LL_040_in_3\ : std_logic;
signal \un1_D_UM_040_3\ : std_logic;
signal \D_UM_AMIGA_in_7\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\ : std_logic;
signal \un1_D_UM_AMIGA_7\ : std_logic;
signal \D_UM_040_in_4\ : std_logic;
signal \D_LL_040_in_4\ : std_logic;
signal \un1_D_UM_040_4\ : std_logic;
signal \D_UM_040_in_7\ : std_logic;
signal \D_LL_040_in_7\ : std_logic;
signal \un1_D_UM_040_7\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\ : std_logic;
signal \D_UU_AMIGA_in_5\ : std_logic;
signal \un1_D_UU_AMIGA_5\ : std_logic;
signal \D_LM_040_in_3\ : std_logic;
signal \D_UU_040_in_3\ : std_logic;
signal \un1_D_UU_040_3\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\ : std_logic;
signal \D_UU_AMIGA_in_4\ : std_logic;
signal \un1_D_UU_AMIGA_4\ : std_logic;
signal \U111_CYCLE_SM.LW_TRANSZ0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\ : std_logic;
signal \PORTSIZE_c\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\ : std_logic;
signal \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa\ : std_logic;
signal \TS_CPUn_c\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\ : std_logic;
signal \U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0\ : std_logic;
signal \CLK40\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U111_CYCLE_SM.BURST_COUNTZ0Z_1\ : std_logic;
signal \U111_CYCLE_SM.BURST_COUNTZ0Z_0\ : std_logic;
signal \TBIn_c\ : std_logic;
signal \U111_CYCLE_SM.BURSTZ0\ : std_logic;
signal \U111_CYCLE_SM.un7_CYCLE_STATE_0\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \U111_CYCLE_SM.PORT_MISMATCHZ0\ : std_logic;
signal \U111_CYCLE_SM.un7_CYCLE_STATE_0_cascade_\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\ : std_logic;
signal \U111_CYCLE_SM.N_136\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\ : std_logic;
signal \D_UM_AMIGA_in_2\ : std_logic;
signal \un1_D_UM_AMIGA_2\ : std_logic;
signal \D_UM_040_in_1\ : std_logic;
signal \D_LL_040_in_1\ : std_logic;
signal \un1_D_UM_040_1\ : std_logic;
signal \D_UM_AMIGA_in_6\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\ : std_logic;
signal \U111_CYCLE_SM.LATCH_ENZ0\ : std_logic;
signal \un1_D_UM_AMIGA_6\ : std_logic;
signal \D_UU_040_in_6\ : std_logic;
signal \D_LM_040_in_6\ : std_logic;
signal \un1_D_UU_040_6\ : std_logic;
signal \D_LM_040_in_5\ : std_logic;
signal \U111_CYCLE_SM.FLIP_WORDZ0\ : std_logic;
signal \D_UU_040_in_5\ : std_logic;
signal \un1_D_UU_040_5\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK40_IN_wire\ : std_logic;
signal \LBENn_wire\ : std_logic;
signal \CPUBGn_wire\ : std_logic;
signal \TEA_CPUn_wire\ : std_logic;
signal \A_040_wire\ : std_logic_vector(1 downto 0);
signal \A_AMIGA_wire\ : std_logic_vector(1 downto 0);
signal \CLK40B_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \BUFDIR_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \TS_CPUn_wire\ : std_logic;
signal \CLKRAMA_wire\ : std_logic;
signal \TCI_CPUn_wire\ : std_logic;
signal \CLKRAMB_wire\ : std_logic;
signal \TEAn_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \DMAn_wire\ : std_logic;
signal \CLK80_CPU_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \TBI_CPUn_wire\ : std_logic;
signal \CLK40A_wire\ : std_logic;
signal \pll_pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK40_IN_wire\ <= CLK40_IN;
    \LBENn_wire\ <= LBENn;
    CPUBGn <= \CPUBGn_wire\;
    TEA_CPUn <= \TEA_CPUn_wire\;
    \A_040_wire\ <= A_040;
    A_AMIGA <= \A_AMIGA_wire\;
    CLK40B <= \CLK40B_wire\;
    \TBIn_wire\ <= TBIn;
    BUFDIR <= \BUFDIR_wire\;
    \SIZ_wire\ <= SIZ;
    \TS_CPUn_wire\ <= TS_CPUn;
    CLKRAMA <= \CLKRAMA_wire\;
    TCI_CPUn <= \TCI_CPUn_wire\;
    CLKRAMB <= \CLKRAMB_wire\;
    \TEAn_wire\ <= TEAn;
    BUFENn <= \BUFENn_wire\;
    \RnW_wire\ <= RnW;
    DMAn <= \DMAn_wire\;
    CLK80_CPU <= \CLK80_CPU_wire\;
    TSn <= \TSn_wire\;
    \PORTSIZE_wire\ <= PORTSIZE;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    \TCIn_wire\ <= TCIn;
    TBI_CPUn <= \TBI_CPUn_wire\;
    CLK40A <= \CLK40A_wire\;
    \pll_pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll_pll\ : PLL40_2F
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            SCLK => '0',
            PLLOUTGLOBALA => \CLK80\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALB => \CLK40\,
            SDI => '0',
            PLLOUTCOREA => OPEN,
            BYPASS => '0',
            RESETB => \N__3121\,
            PLLOUTCOREB => OPEN,
            LOCK => OPEN,
            SDO => OPEN,
            EXTFEEDBACK => '0',
            DYNAMICDELAY => \pll_pll_DYNAMICDELAY_wire\,
            PLLIN => \N__8833\
        );

    \pll_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \VCCG0\,
            DIN => '0',
            DOUT => \N__8833\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \LBENn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8817\,
            DIN => \N__8816\,
            DOUT => \N__8815\,
            PACKAGEPIN => \LBENn_wire\
        );

    \LBENn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8817\,
            PADOUT => \N__8816\,
            PADIN => \N__8815\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \LBENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8808\,
            DIN => \N__8807\,
            DOUT => \N__8806\,
            PACKAGEPIN => D_UM_040(3)
        );

    \D_UM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8808\,
            PADOUT => \N__8807\,
            PADIN => \N__8806\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4585\,
            DIN0 => \D_UM_040_in_3\,
            DOUT0 => \N__6005\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TAn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8799\,
            DIN => \N__8798\,
            DOUT => \N__8797\,
            PACKAGEPIN => TAn
        );

    \TAn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8799\,
            PADOUT => \N__8798\,
            PADIN => \N__8797\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5372\,
            DIN0 => \TAn_in\,
            DOUT0 => \N__7553\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8790\,
            DIN => \N__8789\,
            DOUT => \N__8788\,
            PACKAGEPIN => D_LL_AMIGA(1)
        );

    \D_LL_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8790\,
            PADOUT => \N__8789\,
            PADIN => \N__8788\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4373\,
            DIN0 => \D_LL_AMIGA_in_1\,
            DOUT0 => \N__7334\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8781\,
            DIN => \N__8780\,
            DOUT => \N__8779\,
            PACKAGEPIN => D_UU_AMIGA(5)
        );

    \D_UU_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8781\,
            PADOUT => \N__8780\,
            PADIN => \N__8779\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4337\,
            DIN0 => \D_UU_AMIGA_in_5\,
            DOUT0 => \N__7943\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8772\,
            DIN => \N__8771\,
            DOUT => \N__8770\,
            PACKAGEPIN => D_UU_040(6)
        );

    \D_UU_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8772\,
            PADOUT => \N__8771\,
            PADIN => \N__8770\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4660\,
            DIN0 => \D_UU_040_in_6\,
            DOUT0 => \N__4964\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CPUBGn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8763\,
            DIN => \N__8762\,
            DOUT => \N__8761\,
            PACKAGEPIN => \CPUBGn_wire\
        );

    \CPUBGn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8763\,
            PADOUT => \N__8762\,
            PADIN => \N__8761\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8754\,
            DIN => \N__8753\,
            DOUT => \N__8752\,
            PACKAGEPIN => D_LL_040(7)
        );

    \D_LL_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8754\,
            PADOUT => \N__8753\,
            PADIN => \N__8752\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4726\,
            DIN0 => \D_LL_040_in_7\,
            DOUT0 => \N__3590\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8745\,
            DIN => \N__8744\,
            DOUT => \N__8743\,
            PACKAGEPIN => D_LL_AMIGA(4)
        );

    \D_LL_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8745\,
            PADOUT => \N__8744\,
            PADIN => \N__8743\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4372\,
            DIN0 => \D_LL_AMIGA_in_4\,
            DOUT0 => \N__5797\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8736\,
            DIN => \N__8735\,
            DOUT => \N__8734\,
            PACKAGEPIN => D_UM_AMIGA(3)
        );

    \D_UM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8736\,
            PADOUT => \N__8735\,
            PADIN => \N__8734\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4246\,
            DIN0 => \D_UM_AMIGA_in_3\,
            DOUT0 => \N__5924\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8727\,
            DIN => \N__8726\,
            DOUT => \N__8725\,
            PACKAGEPIN => D_UU_040(3)
        );

    \D_UU_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8727\,
            PADOUT => \N__8726\,
            PADIN => \N__8725\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4701\,
            DIN0 => \D_UU_040_in_3\,
            DOUT0 => \N__6077\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TEA_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8718\,
            DIN => \N__8717\,
            DOUT => \N__8716\,
            PACKAGEPIN => \TEA_CPUn_wire\
        );

    \TEA_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8718\,
            PADOUT => \N__8717\,
            PADIN => \N__8716\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5276\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8709\,
            DIN => \N__8708\,
            DOUT => \N__8707\,
            PACKAGEPIN => \A_040_wire\(1)
        );

    \A_040_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8709\,
            PADOUT => \N__8708\,
            PADIN => \N__8707\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8700\,
            DIN => \N__8699\,
            DOUT => \N__8698\,
            PACKAGEPIN => D_LM_AMIGA(3)
        );

    \D_LM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8700\,
            PADOUT => \N__8699\,
            PADIN => \N__8698\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4304\,
            DIN0 => \D_LM_AMIGA_in_3\,
            DOUT0 => \N__6662\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8691\,
            DIN => \N__8690\,
            DOUT => \N__8689\,
            PACKAGEPIN => D_LM_040(0)
        );

    \D_LM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8691\,
            PADOUT => \N__8690\,
            PADIN => \N__8689\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4727\,
            DIN0 => \D_LM_040_in_0\,
            DOUT0 => \N__4418\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8682\,
            DIN => \N__8681\,
            DOUT => \N__8680\,
            PACKAGEPIN => D_UM_AMIGA(6)
        );

    \D_UM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8682\,
            PADOUT => \N__8681\,
            PADIN => \N__8680\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4336\,
            DIN0 => \D_UM_AMIGA_in_6\,
            DOUT0 => \N__2612\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8673\,
            DIN => \N__8672\,
            DOUT => \N__8671\,
            PACKAGEPIN => D_LM_AMIGA(4)
        );

    \D_LM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8673\,
            PADOUT => \N__8672\,
            PADIN => \N__8671\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4257\,
            DIN0 => \D_LM_AMIGA_in_4\,
            DOUT0 => \N__3551\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8664\,
            DIN => \N__8663\,
            DOUT => \N__8662\,
            PACKAGEPIN => \A_AMIGA_wire\(1)
        );

    \A_AMIGA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8664\,
            PADOUT => \N__8663\,
            PADIN => \N__8662\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2795\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8655\,
            DIN => \N__8654\,
            DOUT => \N__8653\,
            PACKAGEPIN => D_LM_040(7)
        );

    \D_LM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8655\,
            PADOUT => \N__8654\,
            PADIN => \N__8653\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4663\,
            DIN0 => \D_LM_040_in_7\,
            DOUT0 => \N__3167\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8646\,
            DIN => \N__8645\,
            DOUT => \N__8644\,
            PACKAGEPIN => D_UM_040(4)
        );

    \D_UM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8646\,
            PADOUT => \N__8645\,
            PADIN => \N__8644\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4702\,
            DIN0 => \D_UM_040_in_4\,
            DOUT0 => \N__6149\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8637\,
            DIN => \N__8636\,
            DOUT => \N__8635\,
            PACKAGEPIN => \CLK40B_wire\
        );

    \CLK40B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8637\,
            PADOUT => \N__8636\,
            PADIN => \N__8635\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3984\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8628\,
            DIN => \N__8627\,
            DOUT => \N__8626\,
            PACKAGEPIN => D_UU_AMIGA(0)
        );

    \D_UU_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8628\,
            PADOUT => \N__8627\,
            PADIN => \N__8626\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4355\,
            DIN0 => \D_UU_AMIGA_in_0\,
            DOUT0 => \N__3431\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8619\,
            DIN => \N__8618\,
            DOUT => \N__8617\,
            PACKAGEPIN => D_UM_040(1)
        );

    \D_UM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8619\,
            PADOUT => \N__8618\,
            PADIN => \N__8617\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4678\,
            DIN0 => \D_UM_040_in_1\,
            DOUT0 => \N__3308\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8610\,
            DIN => \N__8609\,
            DOUT => \N__8608\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8610\,
            PADOUT => \N__8609\,
            PADIN => \N__8608\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TBIn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8601\,
            DIN => \N__8600\,
            DOUT => \N__8599\,
            PACKAGEPIN => D_LL_040(4)
        );

    \D_LL_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8601\,
            PADOUT => \N__8600\,
            PADIN => \N__8599\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4743\,
            DIN0 => \D_LL_040_in_4\,
            DOUT0 => \N__5072\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8592\,
            DIN => \N__8591\,
            DOUT => \N__8590\,
            PACKAGEPIN => D_LL_AMIGA(7)
        );

    \D_LL_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8592\,
            PADOUT => \N__8591\,
            PADIN => \N__8590\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4338\,
            DIN0 => \D_LL_AMIGA_in_7\,
            DOUT0 => \N__5711\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8583\,
            DIN => \N__8582\,
            DOUT => \N__8581\,
            PACKAGEPIN => D_UU_AMIGA(7)
        );

    \D_UU_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8583\,
            PADOUT => \N__8582\,
            PADIN => \N__8581\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4253\,
            DIN0 => \D_UU_AMIGA_in_7\,
            DOUT0 => \N__3032\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8574\,
            DIN => \N__8573\,
            DOUT => \N__8572\,
            PACKAGEPIN => \BUFDIR_wire\
        );

    \BUFDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8574\,
            PADOUT => \N__8573\,
            PADIN => \N__8572\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7877\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8565\,
            DIN => \N__8564\,
            DOUT => \N__8563\,
            PACKAGEPIN => D_UU_040(4)
        );

    \D_UU_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8565\,
            PADOUT => \N__8564\,
            PADIN => \N__8563\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4657\,
            DIN0 => \D_UU_040_in_4\,
            DOUT0 => \N__6518\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8556\,
            DIN => \N__8555\,
            DOUT => \N__8554\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8556\,
            PADOUT => \N__8555\,
            PADIN => \N__8554\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TS_CPUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8547\,
            DIN => \N__8546\,
            DOUT => \N__8545\,
            PACKAGEPIN => \TS_CPUn_wire\
        );

    \TS_CPUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8547\,
            PADOUT => \N__8546\,
            PADIN => \N__8545\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TS_CPUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8538\,
            DIN => \N__8537\,
            DOUT => \N__8536\,
            PACKAGEPIN => D_LL_040(1)
        );

    \D_LL_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8538\,
            PADOUT => \N__8537\,
            PADIN => \N__8536\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4742\,
            DIN0 => \D_LL_040_in_1\,
            DOUT0 => \N__2723\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8529\,
            DIN => \N__8528\,
            DOUT => \N__8527\,
            PACKAGEPIN => D_UM_AMIGA(5)
        );

    \D_UM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8529\,
            PADOUT => \N__8528\,
            PADIN => \N__8527\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4356\,
            DIN0 => \D_UM_AMIGA_in_5\,
            DOUT0 => \N__3737\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8520\,
            DIN => \N__8519\,
            DOUT => \N__8518\,
            PACKAGEPIN => D_UU_040(1)
        );

    \D_UU_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8520\,
            PADOUT => \N__8519\,
            PADIN => \N__8518\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4703\,
            DIN0 => \D_UU_040_in_1\,
            DOUT0 => \N__3239\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8511\,
            DIN => \N__8510\,
            DOUT => \N__8509\,
            PACKAGEPIN => D_LM_AMIGA(1)
        );

    \D_LM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8511\,
            PADOUT => \N__8510\,
            PADIN => \N__8509\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4256\,
            DIN0 => \D_LM_AMIGA_in_1\,
            DOUT0 => \N__2885\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8502\,
            DIN => \N__8501\,
            DOUT => \N__8500\,
            PACKAGEPIN => D_LM_040(2)
        );

    \D_LM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8502\,
            PADOUT => \N__8501\,
            PADIN => \N__8500\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4637\,
            DIN0 => \D_LM_040_in_2\,
            DOUT0 => \N__5477\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8493\,
            DIN => \N__8492\,
            DOUT => \N__8491\,
            PACKAGEPIN => D_LL_040(5)
        );

    \D_LL_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8493\,
            PADOUT => \N__8492\,
            PADIN => \N__8491\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4728\,
            DIN0 => \D_LL_040_in_5\,
            DOUT0 => \N__3653\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8484\,
            DIN => \N__8483\,
            DOUT => \N__8482\,
            PACKAGEPIN => D_LL_AMIGA(6)
        );

    \D_LL_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8484\,
            PADOUT => \N__8483\,
            PADIN => \N__8482\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4340\,
            DIN0 => \D_LL_AMIGA_in_6\,
            DOUT0 => \N__2657\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8475\,
            DIN => \N__8474\,
            DOUT => \N__8473\,
            PACKAGEPIN => D_UU_AMIGA(6)
        );

    \D_UU_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8475\,
            PADOUT => \N__8474\,
            PADIN => \N__8473\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4254\,
            DIN0 => \D_UU_AMIGA_in_6\,
            DOUT0 => \N__7025\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8466\,
            DIN => \N__8465\,
            DOUT => \N__8464\,
            PACKAGEPIN => D_UM_AMIGA(1)
        );

    \D_UM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8466\,
            PADOUT => \N__8465\,
            PADIN => \N__8464\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4286\,
            DIN0 => \D_UM_AMIGA_in_1\,
            DOUT0 => \N__7286\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8457\,
            DIN => \N__8456\,
            DOUT => \N__8455\,
            PACKAGEPIN => D_UU_040(5)
        );

    \D_UU_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8457\,
            PADOUT => \N__8456\,
            PADIN => \N__8455\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4662\,
            DIN0 => \D_UU_040_in_5\,
            DOUT0 => \N__6683\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8448\,
            DIN => \N__8447\,
            DOUT => \N__8446\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8448\,
            PADOUT => \N__8447\,
            PADIN => \N__8446\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3719\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__2546\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8439\,
            DIN => \N__8438\,
            DOUT => \N__8437\,
            PACKAGEPIN => \CLKRAMA_wire\
        );

    \CLKRAMA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8439\,
            PADOUT => \N__8438\,
            PADIN => \N__8437\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3992\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8430\,
            DIN => \N__8429\,
            DOUT => \N__8428\,
            PACKAGEPIN => D_UM_040(2)
        );

    \D_UM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8430\,
            PADOUT => \N__8429\,
            PADIN => \N__8428\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4648\,
            DIN0 => \D_UM_040_in_2\,
            DOUT0 => \N__7370\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8421\,
            DIN => \N__8420\,
            DOUT => \N__8419\,
            PACKAGEPIN => D_LL_040(2)
        );

    \D_LL_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8421\,
            PADOUT => \N__8420\,
            PADIN => \N__8419\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4730\,
            DIN0 => \D_LL_040_in_2\,
            DOUT0 => \N__5111\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8412\,
            DIN => \N__8411\,
            DOUT => \N__8410\,
            PACKAGEPIN => \TCI_CPUn_wire\
        );

    \TCI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8412\,
            PADOUT => \N__8411\,
            PADIN => \N__8410\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2522\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMB_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8403\,
            DIN => \N__8402\,
            DOUT => \N__8401\,
            PACKAGEPIN => \CLKRAMB_wire\
        );

    \CLKRAMB_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8403\,
            PADOUT => \N__8402\,
            PADIN => \N__8401\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5576\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8394\,
            DIN => \N__8393\,
            DOUT => \N__8392\,
            PACKAGEPIN => D_LL_AMIGA(2)
        );

    \D_LL_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8394\,
            PADOUT => \N__8393\,
            PADIN => \N__8392\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4375\,
            DIN0 => \D_LL_AMIGA_in_2\,
            DOUT0 => \N__4055\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8385\,
            DIN => \N__8384\,
            DOUT => \N__8383\,
            PACKAGEPIN => D_UM_AMIGA(4)
        );

    \D_UM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8385\,
            PADOUT => \N__8384\,
            PADIN => \N__8383\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4303\,
            DIN0 => \D_UM_AMIGA_in_4\,
            DOUT0 => \N__5753\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8376\,
            DIN => \N__8375\,
            DOUT => \N__8374\,
            PACKAGEPIN => D_UU_AMIGA(2)
        );

    \D_UU_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8376\,
            PADOUT => \N__8375\,
            PADIN => \N__8374\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4354\,
            DIN0 => \D_UU_AMIGA_in_2\,
            DOUT0 => \N__3821\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TEAn_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8367\,
            DIN => \N__8366\,
            DOUT => \N__8365\,
            PACKAGEPIN => \TEAn_wire\
        );

    \TEAn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8367\,
            PADOUT => \N__8366\,
            PADIN => \N__8365\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TEAn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8358\,
            DIN => \N__8357\,
            DOUT => \N__8356\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8358\,
            PADOUT => \N__8357\,
            PADIN => \N__8356\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2597\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8349\,
            DIN => \N__8348\,
            DOUT => \N__8347\,
            PACKAGEPIN => D_LM_AMIGA(6)
        );

    \D_LM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8349\,
            PADOUT => \N__8348\,
            PADIN => \N__8347\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4323\,
            DIN0 => \D_LM_AMIGA_in_6\,
            DOUT0 => \N__7067\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8340\,
            DIN => \N__8339\,
            DOUT => \N__8338\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8340\,
            PADOUT => \N__8339\,
            PADIN => \N__8338\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8331\,
            DIN => \N__8330\,
            DOUT => \N__8329\,
            PACKAGEPIN => D_LM_040(5)
        );

    \D_LM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8331\,
            PADOUT => \N__8330\,
            PADIN => \N__8329\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4650\,
            DIN0 => \D_LM_040_in_5\,
            DOUT0 => \N__3203\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8322\,
            DIN => \N__8321\,
            DOUT => \N__8320\,
            PACKAGEPIN => D_UM_040(6)
        );

    \D_UM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8322\,
            PADOUT => \N__8321\,
            PADIN => \N__8320\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4638\,
            DIN0 => \D_UM_040_in_6\,
            DOUT0 => \N__7103\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMAn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8313\,
            DIN => \N__8312\,
            DOUT => \N__8311\,
            PACKAGEPIN => \DMAn_wire\
        );

    \DMAn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8313\,
            PADOUT => \N__8312\,
            PADIN => \N__8311\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3122\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8304\,
            DIN => \N__8303\,
            DOUT => \N__8302\,
            PACKAGEPIN => D_LL_040(6)
        );

    \D_LL_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8304\,
            PADOUT => \N__8303\,
            PADIN => \N__8302\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4729\,
            DIN0 => \D_LL_040_in_6\,
            DOUT0 => \N__3692\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8295\,
            DIN => \N__8294\,
            DOUT => \N__8293\,
            PACKAGEPIN => D_LL_AMIGA(5)
        );

    \D_LL_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8295\,
            PADOUT => \N__8294\,
            PADIN => \N__8293\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4341\,
            DIN0 => \D_LL_AMIGA_in_5\,
            DOUT0 => \N__3803\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8286\,
            DIN => \N__8285\,
            DOUT => \N__8284\,
            PACKAGEPIN => D_UM_AMIGA(0)
        );

    \D_UM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8286\,
            PADOUT => \N__8285\,
            PADIN => \N__8284\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4321\,
            DIN0 => \D_UM_AMIGA_in_0\,
            DOUT0 => \N__2924\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8277\,
            DIN => \N__8276\,
            DOUT => \N__8275\,
            PACKAGEPIN => D_UU_040(2)
        );

    \D_UU_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8277\,
            PADOUT => \N__8276\,
            PADIN => \N__8275\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4574\,
            DIN0 => \D_UU_040_in_2\,
            DOUT0 => \N__4868\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8268\,
            DIN => \N__8267\,
            DOUT => \N__8266\,
            PACKAGEPIN => D_LM_AMIGA(2)
        );

    \D_LM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8268\,
            PADOUT => \N__8267\,
            PADIN => \N__8266\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4320\,
            DIN0 => \D_LM_AMIGA_in_2\,
            DOUT0 => \N__3857\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK80_CPU_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8259\,
            DIN => \N__8258\,
            DOUT => \N__8257\,
            PACKAGEPIN => \CLK80_CPU_wire\
        );

    \CLK80_CPU_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8259\,
            PADOUT => \N__8258\,
            PADIN => \N__8257\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5572\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8250\,
            DIN => \N__8249\,
            DOUT => \N__8248\,
            PACKAGEPIN => D_LL_040(3)
        );

    \D_LL_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8250\,
            PADOUT => \N__8249\,
            PADIN => \N__8248\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4750\,
            DIN0 => \D_LL_040_in_3\,
            DOUT0 => \N__2690\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8241\,
            DIN => \N__8240\,
            DOUT => \N__8239\,
            PACKAGEPIN => D_LM_040(1)
        );

    \D_LM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8241\,
            PADOUT => \N__8240\,
            PADIN => \N__8239\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4636\,
            DIN0 => \D_LM_040_in_1\,
            DOUT0 => \N__3383\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8232\,
            DIN => \N__8231\,
            DOUT => \N__8230\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8232\,
            PADOUT => \N__8231\,
            PADIN => \N__8230\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4394\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8223\,
            DIN => \N__8222\,
            DOUT => \N__8221\,
            PACKAGEPIN => D_UM_AMIGA(7)
        );

    \D_UM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8223\,
            PADOUT => \N__8222\,
            PADIN => \N__8221\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4302\,
            DIN0 => \D_UM_AMIGA_in_7\,
            DOUT0 => \N__5672\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8214\,
            DIN => \N__8213\,
            DOUT => \N__8212\,
            PACKAGEPIN => D_LM_AMIGA(7)
        );

    \D_LM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8214\,
            PADOUT => \N__8213\,
            PADIN => \N__8212\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4322\,
            DIN0 => \D_LM_AMIGA_in_7\,
            DOUT0 => \N__3089\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8205\,
            DIN => \N__8204\,
            DOUT => \N__8203\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8205\,
            PADOUT => \N__8204\,
            PADIN => \N__8203\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \PORTSIZE_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8196\,
            DIN => \N__8195\,
            DOUT => \N__8194\,
            PACKAGEPIN => \A_AMIGA_wire\(0)
        );

    \A_AMIGA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8196\,
            PADOUT => \N__8195\,
            PADIN => \N__8194\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2810\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8187\,
            DIN => \N__8186\,
            DOUT => \N__8185\,
            PACKAGEPIN => D_LM_040(4)
        );

    \D_LM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8187\,
            PADOUT => \N__8186\,
            PADIN => \N__8185\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4674\,
            DIN0 => \D_LM_040_in_4\,
            DOUT0 => \N__2567\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8178\,
            DIN => \N__8177\,
            DOUT => \N__8176\,
            PACKAGEPIN => D_UM_040(7)
        );

    \D_UM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8178\,
            PADOUT => \N__8177\,
            PADIN => \N__8176\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4584\,
            DIN0 => \D_UM_040_in_7\,
            DOUT0 => \N__5843\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8169\,
            DIN => \N__8168\,
            DOUT => \N__8167\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8169\,
            PADOUT => \N__8168\,
            PADIN => \N__8167\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8160\,
            DIN => \N__8159\,
            DOUT => \N__8158\,
            PACKAGEPIN => D_UU_AMIGA(1)
        );

    \D_UU_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8160\,
            PADOUT => \N__8159\,
            PADIN => \N__8158\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4245\,
            DIN0 => \D_UU_AMIGA_in_1\,
            DOUT0 => \N__2843\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8151\,
            DIN => \N__8150\,
            DOUT => \N__8149\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8151\,
            PADOUT => \N__8150\,
            PADIN => \N__8149\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3983\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8142\,
            DIN => \N__8141\,
            DOUT => \N__8140\,
            PACKAGEPIN => D_UM_040(0)
        );

    \D_UM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8142\,
            PADOUT => \N__8141\,
            PADIN => \N__8140\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4649\,
            DIN0 => \D_UM_040_in_0\,
            DOUT0 => \N__3413\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8133\,
            DIN => \N__8132\,
            DOUT => \N__8131\,
            PACKAGEPIN => D_LL_AMIGA(0)
        );

    \D_LL_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8133\,
            PADOUT => \N__8132\,
            PADIN => \N__8131\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4376\,
            DIN0 => \D_LL_AMIGA_in_0\,
            DOUT0 => \N__2963\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8124\,
            DIN => \N__8123\,
            DOUT => \N__8122\,
            PACKAGEPIN => D_UU_AMIGA(4)
        );

    \D_UU_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8124\,
            PADOUT => \N__8123\,
            PADIN => \N__8122\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4353\,
            DIN0 => \D_UU_AMIGA_in_4\,
            DOUT0 => \N__3512\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8115\,
            DIN => \N__8114\,
            DOUT => \N__8113\,
            PACKAGEPIN => D_UU_040(7)
        );

    \D_UU_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8115\,
            PADOUT => \N__8114\,
            PADIN => \N__8113\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4659\,
            DIN0 => \D_UU_040_in_7\,
            DOUT0 => \N__5150\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8106\,
            DIN => \N__8105\,
            DOUT => \N__8104\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8106\,
            PADOUT => \N__8105\,
            PADIN => \N__8104\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8097\,
            DIN => \N__8096\,
            DOUT => \N__8095\,
            PACKAGEPIN => D_LL_040(0)
        );

    \D_LL_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8097\,
            PADOUT => \N__8096\,
            PADIN => \N__8095\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4751\,
            DIN0 => \D_LL_040_in_0\,
            DOUT0 => \N__2762\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8088\,
            DIN => \N__8087\,
            DOUT => \N__8086\,
            PACKAGEPIN => D_UM_AMIGA(2)
        );

    \D_UM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8088\,
            PADOUT => \N__8087\,
            PADIN => \N__8086\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4258\,
            DIN0 => \D_UM_AMIGA_in_2\,
            DOUT0 => \N__4013\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8079\,
            DIN => \N__8078\,
            DOUT => \N__8077\,
            PACKAGEPIN => D_UU_040(0)
        );

    \D_UU_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8079\,
            PADOUT => \N__8078\,
            PADIN => \N__8077\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4658\,
            DIN0 => \D_UU_040_in_0\,
            DOUT0 => \N__4898\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8070\,
            DIN => \N__8069\,
            DOUT => \N__8068\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8070\,
            PADOUT => \N__8069\,
            PADIN => \N__8068\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TCIn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8061\,
            DIN => \N__8060\,
            DOUT => \N__8059\,
            PACKAGEPIN => \A_040_wire\(0)
        );

    \A_040_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8061\,
            PADOUT => \N__8060\,
            PADIN => \N__8059\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8052\,
            DIN => \N__8051\,
            DOUT => \N__8050\,
            PACKAGEPIN => D_LM_AMIGA(0)
        );

    \D_LM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8052\,
            PADOUT => \N__8051\,
            PADIN => \N__8050\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4339\,
            DIN0 => \D_LM_AMIGA_in_0\,
            DOUT0 => \N__3473\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8043\,
            DIN => \N__8042\,
            DOUT => \N__8041\,
            PACKAGEPIN => \TBI_CPUn_wire\
        );

    \TBI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8043\,
            PADOUT => \N__8042\,
            PADIN => \N__8041\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7609\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8034\,
            DIN => \N__8033\,
            DOUT => \N__8032\,
            PACKAGEPIN => \CLK40A_wire\
        );

    \CLK40A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8034\,
            PADOUT => \N__8033\,
            PADIN => \N__8032\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3988\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8025\,
            DIN => \N__8024\,
            DOUT => \N__8023\,
            PACKAGEPIN => D_LM_040(3)
        );

    \D_LM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8025\,
            PADOUT => \N__8024\,
            PADIN => \N__8023\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4592\,
            DIN0 => \D_LM_040_in_3\,
            DOUT0 => \N__3002\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8016\,
            DIN => \N__8015\,
            DOUT => \N__8014\,
            PACKAGEPIN => D_LM_AMIGA(5)
        );

    \D_LM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8016\,
            PADOUT => \N__8015\,
            PADIN => \N__8014\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4279\,
            DIN0 => \D_LM_AMIGA_in_5\,
            DOUT0 => \N__7001\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8007\,
            DIN => \N__8006\,
            DOUT => \N__8005\,
            PACKAGEPIN => D_LM_040(6)
        );

    \D_LM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8007\,
            PADOUT => \N__8006\,
            PADIN => \N__8005\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4639\,
            DIN0 => \D_LM_040_in_6\,
            DOUT0 => \N__3134\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7998\,
            DIN => \N__7997\,
            DOUT => \N__7996\,
            PACKAGEPIN => D_UM_040(5)
        );

    \D_UM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7998\,
            PADOUT => \N__7997\,
            PADIN => \N__7996\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4661\,
            DIN0 => \D_UM_040_in_5\,
            DOUT0 => \N__4796\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7989\,
            DIN => \N__7988\,
            DOUT => \N__7987\,
            PACKAGEPIN => D_LL_AMIGA(3)
        );

    \D_LL_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7989\,
            PADOUT => \N__7988\,
            PADIN => \N__7987\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4374\,
            DIN0 => \D_LL_AMIGA_in_3\,
            DOUT0 => \N__5960\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7980\,
            DIN => \N__7979\,
            DOUT => \N__7978\,
            PACKAGEPIN => D_UU_AMIGA(3)
        );

    \D_UU_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7980\,
            PADOUT => \N__7979\,
            PADIN => \N__7978\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4255\,
            DIN0 => \D_UU_AMIGA_in_3\,
            DOUT0 => \N__6593\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2033\ : InMux
    port map (
            O => \N__7961\,
            I => \N__7958\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__7958\,
            I => \N__7955\
        );

    \I__2031\ : Sp12to4
    port map (
            O => \N__7955\,
            I => \N__7952\
        );

    \I__2030\ : Span12Mux_v
    port map (
            O => \N__7952\,
            I => \N__7949\
        );

    \I__2029\ : Span12Mux_h
    port map (
            O => \N__7949\,
            I => \N__7946\
        );

    \I__2028\ : Odrv12
    port map (
            O => \N__7946\,
            I => \D_UU_040_in_5\
        );

    \I__2027\ : IoInMux
    port map (
            O => \N__7943\,
            I => \N__7940\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__7940\,
            I => \N__7937\
        );

    \I__2025\ : Span4Mux_s3_h
    port map (
            O => \N__7937\,
            I => \N__7934\
        );

    \I__2024\ : Span4Mux_v
    port map (
            O => \N__7934\,
            I => \N__7931\
        );

    \I__2023\ : Sp12to4
    port map (
            O => \N__7931\,
            I => \N__7928\
        );

    \I__2022\ : Span12Mux_s9_h
    port map (
            O => \N__7928\,
            I => \N__7925\
        );

    \I__2021\ : Odrv12
    port map (
            O => \N__7925\,
            I => \un1_D_UU_040_5\
        );

    \I__2020\ : InMux
    port map (
            O => \N__7922\,
            I => \N__7918\
        );

    \I__2019\ : InMux
    port map (
            O => \N__7921\,
            I => \N__7912\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__7918\,
            I => \N__7909\
        );

    \I__2017\ : InMux
    port map (
            O => \N__7917\,
            I => \N__7904\
        );

    \I__2016\ : InMux
    port map (
            O => \N__7916\,
            I => \N__7904\
        );

    \I__2015\ : InMux
    port map (
            O => \N__7915\,
            I => \N__7901\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__7912\,
            I => \N__7898\
        );

    \I__2013\ : Span4Mux_v
    port map (
            O => \N__7909\,
            I => \N__7891\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__7904\,
            I => \N__7891\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__7901\,
            I => \N__7891\
        );

    \I__2010\ : Span4Mux_h
    port map (
            O => \N__7898\,
            I => \N__7886\
        );

    \I__2009\ : Span4Mux_h
    port map (
            O => \N__7891\,
            I => \N__7886\
        );

    \I__2008\ : Sp12to4
    port map (
            O => \N__7886\,
            I => \N__7883\
        );

    \I__2007\ : Span12Mux_v
    port map (
            O => \N__7883\,
            I => \N__7880\
        );

    \I__2006\ : Odrv12
    port map (
            O => \N__7880\,
            I => \TS_CPUn_c\
        );

    \I__2005\ : IoInMux
    port map (
            O => \N__7877\,
            I => \N__7874\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__7874\,
            I => \N__7869\
        );

    \I__2003\ : CascadeMux
    port map (
            O => \N__7873\,
            I => \N__7866\
        );

    \I__2002\ : CascadeMux
    port map (
            O => \N__7872\,
            I => \N__7863\
        );

    \I__2001\ : Span4Mux_s3_v
    port map (
            O => \N__7869\,
            I => \N__7860\
        );

    \I__2000\ : InMux
    port map (
            O => \N__7866\,
            I => \N__7857\
        );

    \I__1999\ : InMux
    port map (
            O => \N__7863\,
            I => \N__7854\
        );

    \I__1998\ : Span4Mux_v
    port map (
            O => \N__7860\,
            I => \N__7851\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__7857\,
            I => \N__7848\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__7854\,
            I => \N__7845\
        );

    \I__1995\ : Span4Mux_v
    port map (
            O => \N__7851\,
            I => \N__7842\
        );

    \I__1994\ : Span4Mux_h
    port map (
            O => \N__7848\,
            I => \N__7839\
        );

    \I__1993\ : Span4Mux_v
    port map (
            O => \N__7845\,
            I => \N__7836\
        );

    \I__1992\ : Sp12to4
    port map (
            O => \N__7842\,
            I => \N__7833\
        );

    \I__1991\ : Span4Mux_v
    port map (
            O => \N__7839\,
            I => \N__7830\
        );

    \I__1990\ : Sp12to4
    port map (
            O => \N__7836\,
            I => \N__7827\
        );

    \I__1989\ : Span12Mux_h
    port map (
            O => \N__7833\,
            I => \N__7822\
        );

    \I__1988\ : Sp12to4
    port map (
            O => \N__7830\,
            I => \N__7822\
        );

    \I__1987\ : Span12Mux_h
    port map (
            O => \N__7827\,
            I => \N__7819\
        );

    \I__1986\ : Span12Mux_h
    port map (
            O => \N__7822\,
            I => \N__7816\
        );

    \I__1985\ : Odrv12
    port map (
            O => \N__7819\,
            I => \RnW_c\
        );

    \I__1984\ : Odrv12
    port map (
            O => \N__7816\,
            I => \RnW_c\
        );

    \I__1983\ : InMux
    port map (
            O => \N__7811\,
            I => \N__7802\
        );

    \I__1982\ : InMux
    port map (
            O => \N__7810\,
            I => \N__7799\
        );

    \I__1981\ : InMux
    port map (
            O => \N__7809\,
            I => \N__7796\
        );

    \I__1980\ : InMux
    port map (
            O => \N__7808\,
            I => \N__7791\
        );

    \I__1979\ : InMux
    port map (
            O => \N__7807\,
            I => \N__7791\
        );

    \I__1978\ : InMux
    port map (
            O => \N__7806\,
            I => \N__7786\
        );

    \I__1977\ : InMux
    port map (
            O => \N__7805\,
            I => \N__7786\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__7802\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__7799\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__7796\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__7791\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__7786\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1971\ : InMux
    port map (
            O => \N__7775\,
            I => \N__7772\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__7772\,
            I => \N__7769\
        );

    \I__1969\ : Span4Mux_v
    port map (
            O => \N__7769\,
            I => \N__7765\
        );

    \I__1968\ : InMux
    port map (
            O => \N__7768\,
            I => \N__7762\
        );

    \I__1967\ : Odrv4
    port map (
            O => \N__7765\,
            I => \U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__7762\,
            I => \U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0\
        );

    \I__1965\ : InMux
    port map (
            O => \N__7757\,
            I => \N__7754\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__7754\,
            I => \N__7745\
        );

    \I__1963\ : ClkMux
    port map (
            O => \N__7753\,
            I => \N__7703\
        );

    \I__1962\ : ClkMux
    port map (
            O => \N__7752\,
            I => \N__7703\
        );

    \I__1961\ : ClkMux
    port map (
            O => \N__7751\,
            I => \N__7703\
        );

    \I__1960\ : ClkMux
    port map (
            O => \N__7750\,
            I => \N__7703\
        );

    \I__1959\ : ClkMux
    port map (
            O => \N__7749\,
            I => \N__7703\
        );

    \I__1958\ : ClkMux
    port map (
            O => \N__7748\,
            I => \N__7703\
        );

    \I__1957\ : Glb2LocalMux
    port map (
            O => \N__7745\,
            I => \N__7703\
        );

    \I__1956\ : ClkMux
    port map (
            O => \N__7744\,
            I => \N__7703\
        );

    \I__1955\ : ClkMux
    port map (
            O => \N__7743\,
            I => \N__7703\
        );

    \I__1954\ : ClkMux
    port map (
            O => \N__7742\,
            I => \N__7703\
        );

    \I__1953\ : ClkMux
    port map (
            O => \N__7741\,
            I => \N__7703\
        );

    \I__1952\ : ClkMux
    port map (
            O => \N__7740\,
            I => \N__7703\
        );

    \I__1951\ : ClkMux
    port map (
            O => \N__7739\,
            I => \N__7703\
        );

    \I__1950\ : ClkMux
    port map (
            O => \N__7738\,
            I => \N__7703\
        );

    \I__1949\ : ClkMux
    port map (
            O => \N__7737\,
            I => \N__7703\
        );

    \I__1948\ : ClkMux
    port map (
            O => \N__7736\,
            I => \N__7703\
        );

    \I__1947\ : GlobalMux
    port map (
            O => \N__7703\,
            I => \CLK40\
        );

    \I__1946\ : SRMux
    port map (
            O => \N__7700\,
            I => \N__7696\
        );

    \I__1945\ : SRMux
    port map (
            O => \N__7699\,
            I => \N__7692\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__7696\,
            I => \N__7688\
        );

    \I__1943\ : SRMux
    port map (
            O => \N__7695\,
            I => \N__7685\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__7692\,
            I => \N__7681\
        );

    \I__1941\ : SRMux
    port map (
            O => \N__7691\,
            I => \N__7678\
        );

    \I__1940\ : Span4Mux_h
    port map (
            O => \N__7688\,
            I => \N__7673\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__7685\,
            I => \N__7673\
        );

    \I__1938\ : SRMux
    port map (
            O => \N__7684\,
            I => \N__7670\
        );

    \I__1937\ : Span4Mux_h
    port map (
            O => \N__7681\,
            I => \N__7665\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__7678\,
            I => \N__7665\
        );

    \I__1935\ : Span4Mux_h
    port map (
            O => \N__7673\,
            I => \N__7662\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__7670\,
            I => \N__7659\
        );

    \I__1933\ : Span4Mux_v
    port map (
            O => \N__7665\,
            I => \N__7656\
        );

    \I__1932\ : Odrv4
    port map (
            O => \N__7662\,
            I => \RESETn_c_i\
        );

    \I__1931\ : Odrv12
    port map (
            O => \N__7659\,
            I => \RESETn_c_i\
        );

    \I__1930\ : Odrv4
    port map (
            O => \N__7656\,
            I => \RESETn_c_i\
        );

    \I__1929\ : InMux
    port map (
            O => \N__7649\,
            I => \N__7645\
        );

    \I__1928\ : InMux
    port map (
            O => \N__7648\,
            I => \N__7642\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__7645\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_1\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__7642\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_1\
        );

    \I__1925\ : InMux
    port map (
            O => \N__7637\,
            I => \N__7630\
        );

    \I__1924\ : InMux
    port map (
            O => \N__7636\,
            I => \N__7630\
        );

    \I__1923\ : InMux
    port map (
            O => \N__7635\,
            I => \N__7627\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__7630\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_0\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__7627\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_0\
        );

    \I__1920\ : CascadeMux
    port map (
            O => \N__7622\,
            I => \N__7619\
        );

    \I__1919\ : InMux
    port map (
            O => \N__7619\,
            I => \N__7616\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__7616\,
            I => \N__7613\
        );

    \I__1917\ : Span4Mux_v
    port map (
            O => \N__7613\,
            I => \N__7610\
        );

    \I__1916\ : Span4Mux_h
    port map (
            O => \N__7610\,
            I => \N__7606\
        );

    \I__1915\ : IoInMux
    port map (
            O => \N__7609\,
            I => \N__7603\
        );

    \I__1914\ : Sp12to4
    port map (
            O => \N__7606\,
            I => \N__7600\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__7603\,
            I => \N__7597\
        );

    \I__1912\ : Span12Mux_v
    port map (
            O => \N__7600\,
            I => \N__7594\
        );

    \I__1911\ : IoSpan4Mux
    port map (
            O => \N__7597\,
            I => \N__7591\
        );

    \I__1910\ : Odrv12
    port map (
            O => \N__7594\,
            I => \TBIn_c\
        );

    \I__1909\ : Odrv4
    port map (
            O => \N__7591\,
            I => \TBIn_c\
        );

    \I__1908\ : InMux
    port map (
            O => \N__7586\,
            I => \N__7579\
        );

    \I__1907\ : InMux
    port map (
            O => \N__7585\,
            I => \N__7574\
        );

    \I__1906\ : InMux
    port map (
            O => \N__7584\,
            I => \N__7574\
        );

    \I__1905\ : InMux
    port map (
            O => \N__7583\,
            I => \N__7571\
        );

    \I__1904\ : InMux
    port map (
            O => \N__7582\,
            I => \N__7568\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__7579\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__7574\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__7571\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__7568\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__1899\ : InMux
    port map (
            O => \N__7559\,
            I => \N__7556\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__7556\,
            I => \U111_CYCLE_SM.un7_CYCLE_STATE_0\
        );

    \I__1897\ : IoInMux
    port map (
            O => \N__7553\,
            I => \N__7549\
        );

    \I__1896\ : CascadeMux
    port map (
            O => \N__7552\,
            I => \N__7545\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__7549\,
            I => \N__7538\
        );

    \I__1894\ : InMux
    port map (
            O => \N__7548\,
            I => \N__7535\
        );

    \I__1893\ : InMux
    port map (
            O => \N__7545\,
            I => \N__7532\
        );

    \I__1892\ : InMux
    port map (
            O => \N__7544\,
            I => \N__7529\
        );

    \I__1891\ : InMux
    port map (
            O => \N__7543\,
            I => \N__7526\
        );

    \I__1890\ : InMux
    port map (
            O => \N__7542\,
            I => \N__7521\
        );

    \I__1889\ : InMux
    port map (
            O => \N__7541\,
            I => \N__7521\
        );

    \I__1888\ : Span4Mux_s1_v
    port map (
            O => \N__7538\,
            I => \N__7518\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__7535\,
            I => \N__7515\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__7532\,
            I => \N__7506\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__7529\,
            I => \N__7506\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__7526\,
            I => \N__7506\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__7521\,
            I => \N__7506\
        );

    \I__1882\ : Sp12to4
    port map (
            O => \N__7518\,
            I => \N__7503\
        );

    \I__1881\ : Span4Mux_v
    port map (
            O => \N__7515\,
            I => \N__7500\
        );

    \I__1880\ : Span4Mux_v
    port map (
            O => \N__7506\,
            I => \N__7497\
        );

    \I__1879\ : Span12Mux_h
    port map (
            O => \N__7503\,
            I => \N__7493\
        );

    \I__1878\ : Sp12to4
    port map (
            O => \N__7500\,
            I => \N__7488\
        );

    \I__1877\ : Sp12to4
    port map (
            O => \N__7497\,
            I => \N__7488\
        );

    \I__1876\ : InMux
    port map (
            O => \N__7496\,
            I => \N__7485\
        );

    \I__1875\ : Span12Mux_v
    port map (
            O => \N__7493\,
            I => \N__7478\
        );

    \I__1874\ : Span12Mux_h
    port map (
            O => \N__7488\,
            I => \N__7478\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__7485\,
            I => \N__7478\
        );

    \I__1872\ : Span12Mux_v
    port map (
            O => \N__7478\,
            I => \N__7475\
        );

    \I__1871\ : Odrv12
    port map (
            O => \N__7475\,
            I => \TACKn_in\
        );

    \I__1870\ : InMux
    port map (
            O => \N__7472\,
            I => \N__7466\
        );

    \I__1869\ : InMux
    port map (
            O => \N__7471\,
            I => \N__7463\
        );

    \I__1868\ : InMux
    port map (
            O => \N__7470\,
            I => \N__7460\
        );

    \I__1867\ : InMux
    port map (
            O => \N__7469\,
            I => \N__7457\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__7466\,
            I => \U111_CYCLE_SM.PORT_MISMATCHZ0\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__7463\,
            I => \U111_CYCLE_SM.PORT_MISMATCHZ0\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__7460\,
            I => \U111_CYCLE_SM.PORT_MISMATCHZ0\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__7457\,
            I => \U111_CYCLE_SM.PORT_MISMATCHZ0\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__7448\,
            I => \U111_CYCLE_SM.un7_CYCLE_STATE_0_cascade_\
        );

    \I__1861\ : InMux
    port map (
            O => \N__7445\,
            I => \N__7438\
        );

    \I__1860\ : InMux
    port map (
            O => \N__7444\,
            I => \N__7435\
        );

    \I__1859\ : InMux
    port map (
            O => \N__7443\,
            I => \N__7432\
        );

    \I__1858\ : InMux
    port map (
            O => \N__7442\,
            I => \N__7427\
        );

    \I__1857\ : InMux
    port map (
            O => \N__7441\,
            I => \N__7427\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__7438\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__7435\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__7432\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__7427\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\
        );

    \I__1852\ : InMux
    port map (
            O => \N__7418\,
            I => \N__7415\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__7415\,
            I => \U111_CYCLE_SM.N_136\
        );

    \I__1850\ : InMux
    port map (
            O => \N__7412\,
            I => \N__7409\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__7409\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\
        );

    \I__1848\ : InMux
    port map (
            O => \N__7406\,
            I => \N__7403\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__7403\,
            I => \N__7400\
        );

    \I__1846\ : Span4Mux_v
    port map (
            O => \N__7400\,
            I => \N__7395\
        );

    \I__1845\ : InMux
    port map (
            O => \N__7399\,
            I => \N__7392\
        );

    \I__1844\ : InMux
    port map (
            O => \N__7398\,
            I => \N__7389\
        );

    \I__1843\ : Span4Mux_v
    port map (
            O => \N__7395\,
            I => \N__7382\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__7392\,
            I => \N__7382\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__7389\,
            I => \N__7382\
        );

    \I__1840\ : Span4Mux_v
    port map (
            O => \N__7382\,
            I => \N__7379\
        );

    \I__1839\ : Sp12to4
    port map (
            O => \N__7379\,
            I => \N__7376\
        );

    \I__1838\ : Span12Mux_h
    port map (
            O => \N__7376\,
            I => \N__7373\
        );

    \I__1837\ : Odrv12
    port map (
            O => \N__7373\,
            I => \D_UM_AMIGA_in_2\
        );

    \I__1836\ : IoInMux
    port map (
            O => \N__7370\,
            I => \N__7367\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__7367\,
            I => \N__7364\
        );

    \I__1834\ : IoSpan4Mux
    port map (
            O => \N__7364\,
            I => \N__7361\
        );

    \I__1833\ : Span4Mux_s2_h
    port map (
            O => \N__7361\,
            I => \N__7358\
        );

    \I__1832\ : Sp12to4
    port map (
            O => \N__7358\,
            I => \N__7355\
        );

    \I__1831\ : Odrv12
    port map (
            O => \N__7355\,
            I => \un1_D_UM_AMIGA_2\
        );

    \I__1830\ : InMux
    port map (
            O => \N__7352\,
            I => \N__7349\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__7349\,
            I => \N__7346\
        );

    \I__1828\ : Sp12to4
    port map (
            O => \N__7346\,
            I => \N__7343\
        );

    \I__1827\ : Span12Mux_v
    port map (
            O => \N__7343\,
            I => \N__7340\
        );

    \I__1826\ : Span12Mux_h
    port map (
            O => \N__7340\,
            I => \N__7337\
        );

    \I__1825\ : Odrv12
    port map (
            O => \N__7337\,
            I => \D_UM_040_in_1\
        );

    \I__1824\ : IoInMux
    port map (
            O => \N__7334\,
            I => \N__7330\
        );

    \I__1823\ : InMux
    port map (
            O => \N__7333\,
            I => \N__7327\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__7330\,
            I => \N__7324\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__7327\,
            I => \N__7321\
        );

    \I__1820\ : Span4Mux_s3_h
    port map (
            O => \N__7324\,
            I => \N__7318\
        );

    \I__1819\ : Span4Mux_h
    port map (
            O => \N__7321\,
            I => \N__7315\
        );

    \I__1818\ : Sp12to4
    port map (
            O => \N__7318\,
            I => \N__7312\
        );

    \I__1817\ : Sp12to4
    port map (
            O => \N__7315\,
            I => \N__7309\
        );

    \I__1816\ : Span12Mux_v
    port map (
            O => \N__7312\,
            I => \N__7306\
        );

    \I__1815\ : Span12Mux_v
    port map (
            O => \N__7309\,
            I => \N__7303\
        );

    \I__1814\ : Span12Mux_h
    port map (
            O => \N__7306\,
            I => \N__7300\
        );

    \I__1813\ : Span12Mux_v
    port map (
            O => \N__7303\,
            I => \N__7297\
        );

    \I__1812\ : Span12Mux_h
    port map (
            O => \N__7300\,
            I => \N__7294\
        );

    \I__1811\ : Span12Mux_h
    port map (
            O => \N__7297\,
            I => \N__7291\
        );

    \I__1810\ : Odrv12
    port map (
            O => \N__7294\,
            I => \D_LL_040_in_1\
        );

    \I__1809\ : Odrv12
    port map (
            O => \N__7291\,
            I => \D_LL_040_in_1\
        );

    \I__1808\ : IoInMux
    port map (
            O => \N__7286\,
            I => \N__7283\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__7283\,
            I => \N__7280\
        );

    \I__1806\ : IoSpan4Mux
    port map (
            O => \N__7280\,
            I => \N__7277\
        );

    \I__1805\ : Sp12to4
    port map (
            O => \N__7277\,
            I => \N__7274\
        );

    \I__1804\ : Span12Mux_h
    port map (
            O => \N__7274\,
            I => \N__7271\
        );

    \I__1803\ : Odrv12
    port map (
            O => \N__7271\,
            I => \un1_D_UM_040_1\
        );

    \I__1802\ : InMux
    port map (
            O => \N__7268\,
            I => \N__7265\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__7265\,
            I => \N__7260\
        );

    \I__1800\ : InMux
    port map (
            O => \N__7264\,
            I => \N__7257\
        );

    \I__1799\ : InMux
    port map (
            O => \N__7263\,
            I => \N__7254\
        );

    \I__1798\ : Span4Mux_v
    port map (
            O => \N__7260\,
            I => \N__7251\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__7257\,
            I => \N__7246\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__7254\,
            I => \N__7246\
        );

    \I__1795\ : Span4Mux_v
    port map (
            O => \N__7251\,
            I => \N__7243\
        );

    \I__1794\ : Span4Mux_v
    port map (
            O => \N__7246\,
            I => \N__7240\
        );

    \I__1793\ : Sp12to4
    port map (
            O => \N__7243\,
            I => \N__7235\
        );

    \I__1792\ : Sp12to4
    port map (
            O => \N__7240\,
            I => \N__7235\
        );

    \I__1791\ : Span12Mux_h
    port map (
            O => \N__7235\,
            I => \N__7232\
        );

    \I__1790\ : Span12Mux_v
    port map (
            O => \N__7232\,
            I => \N__7229\
        );

    \I__1789\ : Odrv12
    port map (
            O => \N__7229\,
            I => \D_UM_AMIGA_in_6\
        );

    \I__1788\ : InMux
    port map (
            O => \N__7226\,
            I => \N__7223\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__7223\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\
        );

    \I__1786\ : InMux
    port map (
            O => \N__7220\,
            I => \N__7213\
        );

    \I__1785\ : InMux
    port map (
            O => \N__7219\,
            I => \N__7213\
        );

    \I__1784\ : InMux
    port map (
            O => \N__7218\,
            I => \N__7210\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__7213\,
            I => \N__7202\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__7210\,
            I => \N__7202\
        );

    \I__1781\ : InMux
    port map (
            O => \N__7209\,
            I => \N__7199\
        );

    \I__1780\ : InMux
    port map (
            O => \N__7208\,
            I => \N__7194\
        );

    \I__1779\ : InMux
    port map (
            O => \N__7207\,
            I => \N__7194\
        );

    \I__1778\ : Span4Mux_v
    port map (
            O => \N__7202\,
            I => \N__7180\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__7199\,
            I => \N__7180\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__7194\,
            I => \N__7180\
        );

    \I__1775\ : InMux
    port map (
            O => \N__7193\,
            I => \N__7173\
        );

    \I__1774\ : InMux
    port map (
            O => \N__7192\,
            I => \N__7173\
        );

    \I__1773\ : InMux
    port map (
            O => \N__7191\,
            I => \N__7173\
        );

    \I__1772\ : InMux
    port map (
            O => \N__7190\,
            I => \N__7168\
        );

    \I__1771\ : InMux
    port map (
            O => \N__7189\,
            I => \N__7165\
        );

    \I__1770\ : InMux
    port map (
            O => \N__7188\,
            I => \N__7162\
        );

    \I__1769\ : InMux
    port map (
            O => \N__7187\,
            I => \N__7159\
        );

    \I__1768\ : Span4Mux_v
    port map (
            O => \N__7180\,
            I => \N__7155\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__7173\,
            I => \N__7152\
        );

    \I__1766\ : InMux
    port map (
            O => \N__7172\,
            I => \N__7147\
        );

    \I__1765\ : InMux
    port map (
            O => \N__7171\,
            I => \N__7147\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__7168\,
            I => \N__7142\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__7165\,
            I => \N__7142\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__7162\,
            I => \N__7137\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__7159\,
            I => \N__7137\
        );

    \I__1760\ : CascadeMux
    port map (
            O => \N__7158\,
            I => \N__7133\
        );

    \I__1759\ : Span4Mux_v
    port map (
            O => \N__7155\,
            I => \N__7130\
        );

    \I__1758\ : Span12Mux_s8_v
    port map (
            O => \N__7152\,
            I => \N__7125\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__7147\,
            I => \N__7125\
        );

    \I__1756\ : Span4Mux_v
    port map (
            O => \N__7142\,
            I => \N__7120\
        );

    \I__1755\ : Span4Mux_v
    port map (
            O => \N__7137\,
            I => \N__7120\
        );

    \I__1754\ : InMux
    port map (
            O => \N__7136\,
            I => \N__7117\
        );

    \I__1753\ : InMux
    port map (
            O => \N__7133\,
            I => \N__7114\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__7130\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__1751\ : Odrv12
    port map (
            O => \N__7125\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__1750\ : Odrv4
    port map (
            O => \N__7120\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__7117\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__7114\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__1747\ : IoInMux
    port map (
            O => \N__7103\,
            I => \N__7100\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__7100\,
            I => \N__7097\
        );

    \I__1745\ : IoSpan4Mux
    port map (
            O => \N__7097\,
            I => \N__7094\
        );

    \I__1744\ : Span4Mux_s3_h
    port map (
            O => \N__7094\,
            I => \N__7091\
        );

    \I__1743\ : Span4Mux_h
    port map (
            O => \N__7091\,
            I => \N__7088\
        );

    \I__1742\ : Span4Mux_h
    port map (
            O => \N__7088\,
            I => \N__7085\
        );

    \I__1741\ : Odrv4
    port map (
            O => \N__7085\,
            I => \un1_D_UM_AMIGA_6\
        );

    \I__1740\ : InMux
    port map (
            O => \N__7082\,
            I => \N__7079\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__7079\,
            I => \N__7076\
        );

    \I__1738\ : Span12Mux_v
    port map (
            O => \N__7076\,
            I => \N__7073\
        );

    \I__1737\ : Span12Mux_h
    port map (
            O => \N__7073\,
            I => \N__7070\
        );

    \I__1736\ : Odrv12
    port map (
            O => \N__7070\,
            I => \D_UU_040_in_6\
        );

    \I__1735\ : IoInMux
    port map (
            O => \N__7067\,
            I => \N__7064\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__7064\,
            I => \N__7061\
        );

    \I__1733\ : Span4Mux_s2_h
    port map (
            O => \N__7061\,
            I => \N__7057\
        );

    \I__1732\ : InMux
    port map (
            O => \N__7060\,
            I => \N__7054\
        );

    \I__1731\ : Span4Mux_v
    port map (
            O => \N__7057\,
            I => \N__7051\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__7054\,
            I => \N__7048\
        );

    \I__1729\ : Sp12to4
    port map (
            O => \N__7051\,
            I => \N__7045\
        );

    \I__1728\ : Sp12to4
    port map (
            O => \N__7048\,
            I => \N__7042\
        );

    \I__1727\ : Span12Mux_h
    port map (
            O => \N__7045\,
            I => \N__7039\
        );

    \I__1726\ : Span12Mux_s11_v
    port map (
            O => \N__7042\,
            I => \N__7036\
        );

    \I__1725\ : Span12Mux_h
    port map (
            O => \N__7039\,
            I => \N__7033\
        );

    \I__1724\ : Span12Mux_h
    port map (
            O => \N__7036\,
            I => \N__7030\
        );

    \I__1723\ : Odrv12
    port map (
            O => \N__7033\,
            I => \D_LM_040_in_6\
        );

    \I__1722\ : Odrv12
    port map (
            O => \N__7030\,
            I => \D_LM_040_in_6\
        );

    \I__1721\ : IoInMux
    port map (
            O => \N__7025\,
            I => \N__7022\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__7022\,
            I => \N__7019\
        );

    \I__1719\ : IoSpan4Mux
    port map (
            O => \N__7019\,
            I => \N__7016\
        );

    \I__1718\ : IoSpan4Mux
    port map (
            O => \N__7016\,
            I => \N__7013\
        );

    \I__1717\ : Span4Mux_s2_v
    port map (
            O => \N__7013\,
            I => \N__7010\
        );

    \I__1716\ : Span4Mux_h
    port map (
            O => \N__7010\,
            I => \N__7007\
        );

    \I__1715\ : Span4Mux_v
    port map (
            O => \N__7007\,
            I => \N__7004\
        );

    \I__1714\ : Odrv4
    port map (
            O => \N__7004\,
            I => \un1_D_UU_040_6\
        );

    \I__1713\ : IoInMux
    port map (
            O => \N__7001\,
            I => \N__6998\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__6998\,
            I => \N__6995\
        );

    \I__1711\ : IoSpan4Mux
    port map (
            O => \N__6995\,
            I => \N__6992\
        );

    \I__1710\ : Span4Mux_s2_h
    port map (
            O => \N__6992\,
            I => \N__6988\
        );

    \I__1709\ : InMux
    port map (
            O => \N__6991\,
            I => \N__6985\
        );

    \I__1708\ : Span4Mux_v
    port map (
            O => \N__6988\,
            I => \N__6982\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__6985\,
            I => \N__6979\
        );

    \I__1706\ : Sp12to4
    port map (
            O => \N__6982\,
            I => \N__6976\
        );

    \I__1705\ : Sp12to4
    port map (
            O => \N__6979\,
            I => \N__6973\
        );

    \I__1704\ : Span12Mux_s9_h
    port map (
            O => \N__6976\,
            I => \N__6970\
        );

    \I__1703\ : Span12Mux_v
    port map (
            O => \N__6973\,
            I => \N__6967\
        );

    \I__1702\ : Span12Mux_h
    port map (
            O => \N__6970\,
            I => \N__6964\
        );

    \I__1701\ : Span12Mux_h
    port map (
            O => \N__6967\,
            I => \N__6961\
        );

    \I__1700\ : Odrv12
    port map (
            O => \N__6964\,
            I => \D_LM_040_in_5\
        );

    \I__1699\ : Odrv12
    port map (
            O => \N__6961\,
            I => \D_LM_040_in_5\
        );

    \I__1698\ : InMux
    port map (
            O => \N__6956\,
            I => \N__6950\
        );

    \I__1697\ : InMux
    port map (
            O => \N__6955\,
            I => \N__6950\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__6950\,
            I => \N__6941\
        );

    \I__1695\ : InMux
    port map (
            O => \N__6949\,
            I => \N__6938\
        );

    \I__1694\ : InMux
    port map (
            O => \N__6948\,
            I => \N__6927\
        );

    \I__1693\ : InMux
    port map (
            O => \N__6947\,
            I => \N__6927\
        );

    \I__1692\ : InMux
    port map (
            O => \N__6946\,
            I => \N__6922\
        );

    \I__1691\ : InMux
    port map (
            O => \N__6945\,
            I => \N__6922\
        );

    \I__1690\ : InMux
    port map (
            O => \N__6944\,
            I => \N__6912\
        );

    \I__1689\ : Span4Mux_v
    port map (
            O => \N__6941\,
            I => \N__6907\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__6938\,
            I => \N__6907\
        );

    \I__1687\ : InMux
    port map (
            O => \N__6937\,
            I => \N__6900\
        );

    \I__1686\ : InMux
    port map (
            O => \N__6936\,
            I => \N__6900\
        );

    \I__1685\ : InMux
    port map (
            O => \N__6935\,
            I => \N__6900\
        );

    \I__1684\ : InMux
    port map (
            O => \N__6934\,
            I => \N__6895\
        );

    \I__1683\ : InMux
    port map (
            O => \N__6933\,
            I => \N__6890\
        );

    \I__1682\ : InMux
    port map (
            O => \N__6932\,
            I => \N__6890\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__6927\,
            I => \N__6885\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__6922\,
            I => \N__6885\
        );

    \I__1679\ : InMux
    port map (
            O => \N__6921\,
            I => \N__6882\
        );

    \I__1678\ : InMux
    port map (
            O => \N__6920\,
            I => \N__6877\
        );

    \I__1677\ : InMux
    port map (
            O => \N__6919\,
            I => \N__6870\
        );

    \I__1676\ : InMux
    port map (
            O => \N__6918\,
            I => \N__6870\
        );

    \I__1675\ : InMux
    port map (
            O => \N__6917\,
            I => \N__6870\
        );

    \I__1674\ : InMux
    port map (
            O => \N__6916\,
            I => \N__6865\
        );

    \I__1673\ : InMux
    port map (
            O => \N__6915\,
            I => \N__6865\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__6912\,
            I => \N__6858\
        );

    \I__1671\ : Span4Mux_h
    port map (
            O => \N__6907\,
            I => \N__6858\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__6900\,
            I => \N__6858\
        );

    \I__1669\ : InMux
    port map (
            O => \N__6899\,
            I => \N__6855\
        );

    \I__1668\ : InMux
    port map (
            O => \N__6898\,
            I => \N__6852\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__6895\,
            I => \N__6847\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__6890\,
            I => \N__6847\
        );

    \I__1665\ : Span4Mux_v
    port map (
            O => \N__6885\,
            I => \N__6843\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__6882\,
            I => \N__6840\
        );

    \I__1663\ : InMux
    port map (
            O => \N__6881\,
            I => \N__6835\
        );

    \I__1662\ : InMux
    port map (
            O => \N__6880\,
            I => \N__6835\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__6877\,
            I => \N__6828\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__6870\,
            I => \N__6825\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__6865\,
            I => \N__6822\
        );

    \I__1658\ : Span4Mux_v
    port map (
            O => \N__6858\,
            I => \N__6815\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__6855\,
            I => \N__6815\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__6852\,
            I => \N__6815\
        );

    \I__1655\ : Span4Mux_v
    port map (
            O => \N__6847\,
            I => \N__6812\
        );

    \I__1654\ : InMux
    port map (
            O => \N__6846\,
            I => \N__6809\
        );

    \I__1653\ : Span4Mux_v
    port map (
            O => \N__6843\,
            I => \N__6802\
        );

    \I__1652\ : Span4Mux_h
    port map (
            O => \N__6840\,
            I => \N__6802\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__6835\,
            I => \N__6802\
        );

    \I__1650\ : InMux
    port map (
            O => \N__6834\,
            I => \N__6797\
        );

    \I__1649\ : InMux
    port map (
            O => \N__6833\,
            I => \N__6797\
        );

    \I__1648\ : InMux
    port map (
            O => \N__6832\,
            I => \N__6792\
        );

    \I__1647\ : InMux
    port map (
            O => \N__6831\,
            I => \N__6792\
        );

    \I__1646\ : Span12Mux_v
    port map (
            O => \N__6828\,
            I => \N__6784\
        );

    \I__1645\ : Span12Mux_v
    port map (
            O => \N__6825\,
            I => \N__6784\
        );

    \I__1644\ : Span12Mux_v
    port map (
            O => \N__6822\,
            I => \N__6781\
        );

    \I__1643\ : Span4Mux_v
    port map (
            O => \N__6815\,
            I => \N__6778\
        );

    \I__1642\ : Span4Mux_v
    port map (
            O => \N__6812\,
            I => \N__6773\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__6809\,
            I => \N__6773\
        );

    \I__1640\ : Span4Mux_v
    port map (
            O => \N__6802\,
            I => \N__6770\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__6797\,
            I => \N__6765\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__6792\,
            I => \N__6765\
        );

    \I__1637\ : InMux
    port map (
            O => \N__6791\,
            I => \N__6762\
        );

    \I__1636\ : InMux
    port map (
            O => \N__6790\,
            I => \N__6759\
        );

    \I__1635\ : InMux
    port map (
            O => \N__6789\,
            I => \N__6756\
        );

    \I__1634\ : Odrv12
    port map (
            O => \N__6784\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1633\ : Odrv12
    port map (
            O => \N__6781\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1632\ : Odrv4
    port map (
            O => \N__6778\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1631\ : Odrv4
    port map (
            O => \N__6773\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1630\ : Odrv4
    port map (
            O => \N__6770\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1629\ : Odrv12
    port map (
            O => \N__6765\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__6762\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__6759\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__6756\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1625\ : InMux
    port map (
            O => \N__6737\,
            I => \N__6734\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__6734\,
            I => \N__6731\
        );

    \I__1623\ : Odrv12
    port map (
            O => \N__6731\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\
        );

    \I__1622\ : InMux
    port map (
            O => \N__6728\,
            I => \N__6724\
        );

    \I__1621\ : InMux
    port map (
            O => \N__6727\,
            I => \N__6721\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__6724\,
            I => \N__6718\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__6721\,
            I => \N__6714\
        );

    \I__1618\ : Span4Mux_v
    port map (
            O => \N__6718\,
            I => \N__6711\
        );

    \I__1617\ : InMux
    port map (
            O => \N__6717\,
            I => \N__6708\
        );

    \I__1616\ : Span4Mux_v
    port map (
            O => \N__6714\,
            I => \N__6705\
        );

    \I__1615\ : Span4Mux_v
    port map (
            O => \N__6711\,
            I => \N__6700\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__6708\,
            I => \N__6700\
        );

    \I__1613\ : Span4Mux_v
    port map (
            O => \N__6705\,
            I => \N__6695\
        );

    \I__1612\ : Span4Mux_h
    port map (
            O => \N__6700\,
            I => \N__6695\
        );

    \I__1611\ : Span4Mux_v
    port map (
            O => \N__6695\,
            I => \N__6692\
        );

    \I__1610\ : Sp12to4
    port map (
            O => \N__6692\,
            I => \N__6689\
        );

    \I__1609\ : Span12Mux_h
    port map (
            O => \N__6689\,
            I => \N__6686\
        );

    \I__1608\ : Odrv12
    port map (
            O => \N__6686\,
            I => \D_UU_AMIGA_in_5\
        );

    \I__1607\ : IoInMux
    port map (
            O => \N__6683\,
            I => \N__6680\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__6680\,
            I => \N__6677\
        );

    \I__1605\ : IoSpan4Mux
    port map (
            O => \N__6677\,
            I => \N__6674\
        );

    \I__1604\ : IoSpan4Mux
    port map (
            O => \N__6674\,
            I => \N__6671\
        );

    \I__1603\ : Sp12to4
    port map (
            O => \N__6671\,
            I => \N__6668\
        );

    \I__1602\ : Span12Mux_s6_v
    port map (
            O => \N__6668\,
            I => \N__6665\
        );

    \I__1601\ : Odrv12
    port map (
            O => \N__6665\,
            I => \un1_D_UU_AMIGA_5\
        );

    \I__1600\ : IoInMux
    port map (
            O => \N__6662\,
            I => \N__6659\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__6659\,
            I => \N__6656\
        );

    \I__1598\ : IoSpan4Mux
    port map (
            O => \N__6656\,
            I => \N__6652\
        );

    \I__1597\ : InMux
    port map (
            O => \N__6655\,
            I => \N__6649\
        );

    \I__1596\ : IoSpan4Mux
    port map (
            O => \N__6652\,
            I => \N__6646\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__6649\,
            I => \N__6643\
        );

    \I__1594\ : Span4Mux_s2_h
    port map (
            O => \N__6646\,
            I => \N__6640\
        );

    \I__1593\ : Span4Mux_v
    port map (
            O => \N__6643\,
            I => \N__6637\
        );

    \I__1592\ : Sp12to4
    port map (
            O => \N__6640\,
            I => \N__6634\
        );

    \I__1591\ : Sp12to4
    port map (
            O => \N__6637\,
            I => \N__6631\
        );

    \I__1590\ : Span12Mux_h
    port map (
            O => \N__6634\,
            I => \N__6628\
        );

    \I__1589\ : Span12Mux_h
    port map (
            O => \N__6631\,
            I => \N__6625\
        );

    \I__1588\ : Span12Mux_h
    port map (
            O => \N__6628\,
            I => \N__6622\
        );

    \I__1587\ : Span12Mux_v
    port map (
            O => \N__6625\,
            I => \N__6619\
        );

    \I__1586\ : Odrv12
    port map (
            O => \N__6622\,
            I => \D_LM_040_in_3\
        );

    \I__1585\ : Odrv12
    port map (
            O => \N__6619\,
            I => \D_LM_040_in_3\
        );

    \I__1584\ : InMux
    port map (
            O => \N__6614\,
            I => \N__6611\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__6611\,
            I => \N__6608\
        );

    \I__1582\ : Span4Mux_v
    port map (
            O => \N__6608\,
            I => \N__6605\
        );

    \I__1581\ : Span4Mux_h
    port map (
            O => \N__6605\,
            I => \N__6602\
        );

    \I__1580\ : Sp12to4
    port map (
            O => \N__6602\,
            I => \N__6599\
        );

    \I__1579\ : Span12Mux_h
    port map (
            O => \N__6599\,
            I => \N__6596\
        );

    \I__1578\ : Odrv12
    port map (
            O => \N__6596\,
            I => \D_UU_040_in_3\
        );

    \I__1577\ : IoInMux
    port map (
            O => \N__6593\,
            I => \N__6590\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__6590\,
            I => \N__6587\
        );

    \I__1575\ : Span4Mux_s2_v
    port map (
            O => \N__6587\,
            I => \N__6584\
        );

    \I__1574\ : Span4Mux_v
    port map (
            O => \N__6584\,
            I => \N__6581\
        );

    \I__1573\ : Sp12to4
    port map (
            O => \N__6581\,
            I => \N__6578\
        );

    \I__1572\ : Span12Mux_h
    port map (
            O => \N__6578\,
            I => \N__6575\
        );

    \I__1571\ : Odrv12
    port map (
            O => \N__6575\,
            I => \un1_D_UU_040_3\
        );

    \I__1570\ : InMux
    port map (
            O => \N__6572\,
            I => \N__6569\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__6569\,
            I => \N__6566\
        );

    \I__1568\ : Odrv12
    port map (
            O => \N__6566\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\
        );

    \I__1567\ : InMux
    port map (
            O => \N__6563\,
            I => \N__6559\
        );

    \I__1566\ : InMux
    port map (
            O => \N__6562\,
            I => \N__6556\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__6559\,
            I => \N__6553\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__6556\,
            I => \N__6550\
        );

    \I__1563\ : Span4Mux_v
    port map (
            O => \N__6553\,
            I => \N__6546\
        );

    \I__1562\ : Span4Mux_v
    port map (
            O => \N__6550\,
            I => \N__6543\
        );

    \I__1561\ : InMux
    port map (
            O => \N__6549\,
            I => \N__6540\
        );

    \I__1560\ : Span4Mux_v
    port map (
            O => \N__6546\,
            I => \N__6537\
        );

    \I__1559\ : Span4Mux_v
    port map (
            O => \N__6543\,
            I => \N__6532\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__6540\,
            I => \N__6532\
        );

    \I__1557\ : Span4Mux_v
    port map (
            O => \N__6537\,
            I => \N__6527\
        );

    \I__1556\ : Span4Mux_v
    port map (
            O => \N__6532\,
            I => \N__6527\
        );

    \I__1555\ : Sp12to4
    port map (
            O => \N__6527\,
            I => \N__6524\
        );

    \I__1554\ : Span12Mux_h
    port map (
            O => \N__6524\,
            I => \N__6521\
        );

    \I__1553\ : Odrv12
    port map (
            O => \N__6521\,
            I => \D_UU_AMIGA_in_4\
        );

    \I__1552\ : IoInMux
    port map (
            O => \N__6518\,
            I => \N__6515\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__6515\,
            I => \N__6512\
        );

    \I__1550\ : IoSpan4Mux
    port map (
            O => \N__6512\,
            I => \N__6509\
        );

    \I__1549\ : Sp12to4
    port map (
            O => \N__6509\,
            I => \N__6506\
        );

    \I__1548\ : Span12Mux_s6_v
    port map (
            O => \N__6506\,
            I => \N__6503\
        );

    \I__1547\ : Odrv12
    port map (
            O => \N__6503\,
            I => \un1_D_UU_AMIGA_4\
        );

    \I__1546\ : InMux
    port map (
            O => \N__6500\,
            I => \N__6495\
        );

    \I__1545\ : InMux
    port map (
            O => \N__6499\,
            I => \N__6490\
        );

    \I__1544\ : InMux
    port map (
            O => \N__6498\,
            I => \N__6490\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__6495\,
            I => \N__6487\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__6490\,
            I => \U111_CYCLE_SM.LW_TRANSZ0\
        );

    \I__1541\ : Odrv4
    port map (
            O => \N__6487\,
            I => \U111_CYCLE_SM.LW_TRANSZ0\
        );

    \I__1540\ : CascadeMux
    port map (
            O => \N__6482\,
            I => \N__6478\
        );

    \I__1539\ : InMux
    port map (
            O => \N__6481\,
            I => \N__6474\
        );

    \I__1538\ : InMux
    port map (
            O => \N__6478\,
            I => \N__6471\
        );

    \I__1537\ : InMux
    port map (
            O => \N__6477\,
            I => \N__6467\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__6474\,
            I => \N__6464\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__6471\,
            I => \N__6460\
        );

    \I__1534\ : InMux
    port map (
            O => \N__6470\,
            I => \N__6457\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__6467\,
            I => \N__6454\
        );

    \I__1532\ : Span4Mux_h
    port map (
            O => \N__6464\,
            I => \N__6451\
        );

    \I__1531\ : InMux
    port map (
            O => \N__6463\,
            I => \N__6448\
        );

    \I__1530\ : Odrv4
    port map (
            O => \N__6460\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__6457\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1528\ : Odrv4
    port map (
            O => \N__6454\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1527\ : Odrv4
    port map (
            O => \N__6451\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__6448\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1525\ : InMux
    port map (
            O => \N__6437\,
            I => \N__6432\
        );

    \I__1524\ : InMux
    port map (
            O => \N__6436\,
            I => \N__6429\
        );

    \I__1523\ : InMux
    port map (
            O => \N__6435\,
            I => \N__6426\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__6432\,
            I => \N__6421\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__6429\,
            I => \N__6421\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__6426\,
            I => \N__6418\
        );

    \I__1519\ : Span12Mux_h
    port map (
            O => \N__6421\,
            I => \N__6415\
        );

    \I__1518\ : Span12Mux_h
    port map (
            O => \N__6418\,
            I => \N__6412\
        );

    \I__1517\ : Span12Mux_v
    port map (
            O => \N__6415\,
            I => \N__6409\
        );

    \I__1516\ : Span12Mux_v
    port map (
            O => \N__6412\,
            I => \N__6406\
        );

    \I__1515\ : Odrv12
    port map (
            O => \N__6409\,
            I => \PORTSIZE_c\
        );

    \I__1514\ : Odrv12
    port map (
            O => \N__6406\,
            I => \PORTSIZE_c\
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__6401\,
            I => \N__6398\
        );

    \I__1512\ : InMux
    port map (
            O => \N__6398\,
            I => \N__6392\
        );

    \I__1511\ : InMux
    port map (
            O => \N__6397\,
            I => \N__6392\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__6392\,
            I => \N__6389\
        );

    \I__1509\ : Span12Mux_h
    port map (
            O => \N__6389\,
            I => \N__6386\
        );

    \I__1508\ : Span12Mux_v
    port map (
            O => \N__6386\,
            I => \N__6383\
        );

    \I__1507\ : Odrv12
    port map (
            O => \N__6383\,
            I => \SIZ_c_1\
        );

    \I__1506\ : CascadeMux
    port map (
            O => \N__6380\,
            I => \N__6376\
        );

    \I__1505\ : InMux
    port map (
            O => \N__6379\,
            I => \N__6371\
        );

    \I__1504\ : InMux
    port map (
            O => \N__6376\,
            I => \N__6371\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__6371\,
            I => \N__6368\
        );

    \I__1502\ : Span12Mux_h
    port map (
            O => \N__6368\,
            I => \N__6365\
        );

    \I__1501\ : Span12Mux_v
    port map (
            O => \N__6365\,
            I => \N__6362\
        );

    \I__1500\ : Odrv12
    port map (
            O => \N__6362\,
            I => \SIZ_c_0\
        );

    \I__1499\ : CascadeMux
    port map (
            O => \N__6359\,
            I => \N__6354\
        );

    \I__1498\ : InMux
    port map (
            O => \N__6358\,
            I => \N__6343\
        );

    \I__1497\ : InMux
    port map (
            O => \N__6357\,
            I => \N__6343\
        );

    \I__1496\ : InMux
    port map (
            O => \N__6354\,
            I => \N__6343\
        );

    \I__1495\ : InMux
    port map (
            O => \N__6353\,
            I => \N__6343\
        );

    \I__1494\ : InMux
    port map (
            O => \N__6352\,
            I => \N__6340\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__6343\,
            I => \N__6337\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__6340\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\
        );

    \I__1491\ : Odrv4
    port map (
            O => \N__6337\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\
        );

    \I__1490\ : InMux
    port map (
            O => \N__6332\,
            I => \N__6323\
        );

    \I__1489\ : InMux
    port map (
            O => \N__6331\,
            I => \N__6323\
        );

    \I__1488\ : InMux
    port map (
            O => \N__6330\,
            I => \N__6320\
        );

    \I__1487\ : InMux
    port map (
            O => \N__6329\,
            I => \N__6315\
        );

    \I__1486\ : InMux
    port map (
            O => \N__6328\,
            I => \N__6315\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__6323\,
            I => \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__6320\,
            I => \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__6315\,
            I => \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa\
        );

    \I__1482\ : CEMux
    port map (
            O => \N__6308\,
            I => \N__6303\
        );

    \I__1481\ : CEMux
    port map (
            O => \N__6307\,
            I => \N__6299\
        );

    \I__1480\ : CEMux
    port map (
            O => \N__6306\,
            I => \N__6296\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__6303\,
            I => \N__6292\
        );

    \I__1478\ : CEMux
    port map (
            O => \N__6302\,
            I => \N__6289\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__6299\,
            I => \N__6285\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__6296\,
            I => \N__6282\
        );

    \I__1475\ : CEMux
    port map (
            O => \N__6295\,
            I => \N__6279\
        );

    \I__1474\ : Span4Mux_h
    port map (
            O => \N__6292\,
            I => \N__6274\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__6289\,
            I => \N__6274\
        );

    \I__1472\ : CEMux
    port map (
            O => \N__6288\,
            I => \N__6271\
        );

    \I__1471\ : Span4Mux_v
    port map (
            O => \N__6285\,
            I => \N__6266\
        );

    \I__1470\ : Span4Mux_v
    port map (
            O => \N__6282\,
            I => \N__6266\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__6279\,
            I => \N__6263\
        );

    \I__1468\ : Span4Mux_h
    port map (
            O => \N__6274\,
            I => \N__6260\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__6271\,
            I => \N__6257\
        );

    \I__1466\ : Odrv4
    port map (
            O => \N__6266\,
            I => \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0\
        );

    \I__1465\ : Odrv4
    port map (
            O => \N__6263\,
            I => \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0\
        );

    \I__1464\ : Odrv4
    port map (
            O => \N__6260\,
            I => \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0\
        );

    \I__1463\ : Odrv4
    port map (
            O => \N__6257\,
            I => \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0\
        );

    \I__1462\ : SRMux
    port map (
            O => \N__6248\,
            I => \N__6240\
        );

    \I__1461\ : SRMux
    port map (
            O => \N__6247\,
            I => \N__6237\
        );

    \I__1460\ : SRMux
    port map (
            O => \N__6246\,
            I => \N__6234\
        );

    \I__1459\ : SRMux
    port map (
            O => \N__6245\,
            I => \N__6231\
        );

    \I__1458\ : SRMux
    port map (
            O => \N__6244\,
            I => \N__6228\
        );

    \I__1457\ : SRMux
    port map (
            O => \N__6243\,
            I => \N__6225\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__6240\,
            I => \N__6222\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__6237\,
            I => \N__6215\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__6234\,
            I => \N__6215\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__6231\,
            I => \N__6215\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__6228\,
            I => \N__6210\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__6225\,
            I => \N__6210\
        );

    \I__1450\ : Odrv4
    port map (
            O => \N__6222\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81\
        );

    \I__1449\ : Odrv4
    port map (
            O => \N__6215\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81\
        );

    \I__1448\ : Odrv4
    port map (
            O => \N__6210\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81\
        );

    \I__1447\ : InMux
    port map (
            O => \N__6203\,
            I => \N__6200\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__6200\,
            I => \N__6197\
        );

    \I__1445\ : Span4Mux_v
    port map (
            O => \N__6197\,
            I => \N__6194\
        );

    \I__1444\ : Span4Mux_v
    port map (
            O => \N__6194\,
            I => \N__6190\
        );

    \I__1443\ : InMux
    port map (
            O => \N__6193\,
            I => \N__6187\
        );

    \I__1442\ : Span4Mux_v
    port map (
            O => \N__6190\,
            I => \N__6181\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__6187\,
            I => \N__6181\
        );

    \I__1440\ : InMux
    port map (
            O => \N__6186\,
            I => \N__6178\
        );

    \I__1439\ : Span4Mux_h
    port map (
            O => \N__6181\,
            I => \N__6173\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__6178\,
            I => \N__6173\
        );

    \I__1437\ : Span4Mux_v
    port map (
            O => \N__6173\,
            I => \N__6170\
        );

    \I__1436\ : Span4Mux_v
    port map (
            O => \N__6170\,
            I => \N__6167\
        );

    \I__1435\ : Sp12to4
    port map (
            O => \N__6167\,
            I => \N__6164\
        );

    \I__1434\ : Span12Mux_h
    port map (
            O => \N__6164\,
            I => \N__6161\
        );

    \I__1433\ : Odrv12
    port map (
            O => \N__6161\,
            I => \D_UM_AMIGA_in_4\
        );

    \I__1432\ : InMux
    port map (
            O => \N__6158\,
            I => \N__6155\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__6155\,
            I => \N__6152\
        );

    \I__1430\ : Odrv4
    port map (
            O => \N__6152\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\
        );

    \I__1429\ : IoInMux
    port map (
            O => \N__6149\,
            I => \N__6146\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__6146\,
            I => \N__6143\
        );

    \I__1427\ : IoSpan4Mux
    port map (
            O => \N__6143\,
            I => \N__6140\
        );

    \I__1426\ : Sp12to4
    port map (
            O => \N__6140\,
            I => \N__6137\
        );

    \I__1425\ : Span12Mux_s6_v
    port map (
            O => \N__6137\,
            I => \N__6134\
        );

    \I__1424\ : Span12Mux_h
    port map (
            O => \N__6134\,
            I => \N__6131\
        );

    \I__1423\ : Odrv12
    port map (
            O => \N__6131\,
            I => \un1_D_UM_AMIGA_4\
        );

    \I__1422\ : InMux
    port map (
            O => \N__6128\,
            I => \N__6125\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__6125\,
            I => \N__6122\
        );

    \I__1420\ : Odrv4
    port map (
            O => \N__6122\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\
        );

    \I__1419\ : InMux
    port map (
            O => \N__6119\,
            I => \N__6115\
        );

    \I__1418\ : InMux
    port map (
            O => \N__6118\,
            I => \N__6112\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__6115\,
            I => \N__6109\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__6112\,
            I => \N__6105\
        );

    \I__1415\ : Span4Mux_v
    port map (
            O => \N__6109\,
            I => \N__6102\
        );

    \I__1414\ : InMux
    port map (
            O => \N__6108\,
            I => \N__6099\
        );

    \I__1413\ : Span4Mux_v
    port map (
            O => \N__6105\,
            I => \N__6096\
        );

    \I__1412\ : Span4Mux_v
    port map (
            O => \N__6102\,
            I => \N__6093\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__6099\,
            I => \N__6090\
        );

    \I__1410\ : Sp12to4
    port map (
            O => \N__6096\,
            I => \N__6083\
        );

    \I__1409\ : Sp12to4
    port map (
            O => \N__6093\,
            I => \N__6083\
        );

    \I__1408\ : Span12Mux_h
    port map (
            O => \N__6090\,
            I => \N__6083\
        );

    \I__1407\ : Span12Mux_h
    port map (
            O => \N__6083\,
            I => \N__6080\
        );

    \I__1406\ : Odrv12
    port map (
            O => \N__6080\,
            I => \D_UU_AMIGA_in_3\
        );

    \I__1405\ : IoInMux
    port map (
            O => \N__6077\,
            I => \N__6074\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__6074\,
            I => \N__6071\
        );

    \I__1403\ : Span12Mux_s9_v
    port map (
            O => \N__6071\,
            I => \N__6068\
        );

    \I__1402\ : Span12Mux_h
    port map (
            O => \N__6068\,
            I => \N__6065\
        );

    \I__1401\ : Odrv12
    port map (
            O => \N__6065\,
            I => \un1_D_UU_AMIGA_3\
        );

    \I__1400\ : InMux
    port map (
            O => \N__6062\,
            I => \N__6059\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__6059\,
            I => \N__6056\
        );

    \I__1398\ : Odrv12
    port map (
            O => \N__6056\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\
        );

    \I__1397\ : InMux
    port map (
            O => \N__6053\,
            I => \N__6049\
        );

    \I__1396\ : InMux
    port map (
            O => \N__6052\,
            I => \N__6046\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__6049\,
            I => \N__6042\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__6046\,
            I => \N__6039\
        );

    \I__1393\ : InMux
    port map (
            O => \N__6045\,
            I => \N__6036\
        );

    \I__1392\ : Span4Mux_h
    port map (
            O => \N__6042\,
            I => \N__6033\
        );

    \I__1391\ : Span4Mux_v
    port map (
            O => \N__6039\,
            I => \N__6028\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__6036\,
            I => \N__6028\
        );

    \I__1389\ : Span4Mux_v
    port map (
            O => \N__6033\,
            I => \N__6025\
        );

    \I__1388\ : Span4Mux_v
    port map (
            O => \N__6028\,
            I => \N__6022\
        );

    \I__1387\ : Sp12to4
    port map (
            O => \N__6025\,
            I => \N__6019\
        );

    \I__1386\ : Sp12to4
    port map (
            O => \N__6022\,
            I => \N__6016\
        );

    \I__1385\ : Span12Mux_v
    port map (
            O => \N__6019\,
            I => \N__6013\
        );

    \I__1384\ : Span12Mux_h
    port map (
            O => \N__6016\,
            I => \N__6010\
        );

    \I__1383\ : Odrv12
    port map (
            O => \N__6013\,
            I => \D_UM_AMIGA_in_3\
        );

    \I__1382\ : Odrv12
    port map (
            O => \N__6010\,
            I => \D_UM_AMIGA_in_3\
        );

    \I__1381\ : IoInMux
    port map (
            O => \N__6005\,
            I => \N__6002\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__6002\,
            I => \N__5999\
        );

    \I__1379\ : Span4Mux_s3_h
    port map (
            O => \N__5999\,
            I => \N__5996\
        );

    \I__1378\ : Span4Mux_h
    port map (
            O => \N__5996\,
            I => \N__5993\
        );

    \I__1377\ : Span4Mux_h
    port map (
            O => \N__5993\,
            I => \N__5990\
        );

    \I__1376\ : Span4Mux_h
    port map (
            O => \N__5990\,
            I => \N__5987\
        );

    \I__1375\ : Span4Mux_v
    port map (
            O => \N__5987\,
            I => \N__5984\
        );

    \I__1374\ : Odrv4
    port map (
            O => \N__5984\,
            I => \un1_D_UM_AMIGA_3\
        );

    \I__1373\ : InMux
    port map (
            O => \N__5981\,
            I => \N__5978\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__5978\,
            I => \N__5975\
        );

    \I__1371\ : Span4Mux_v
    port map (
            O => \N__5975\,
            I => \N__5972\
        );

    \I__1370\ : Span4Mux_v
    port map (
            O => \N__5972\,
            I => \N__5969\
        );

    \I__1369\ : Sp12to4
    port map (
            O => \N__5969\,
            I => \N__5966\
        );

    \I__1368\ : Span12Mux_h
    port map (
            O => \N__5966\,
            I => \N__5963\
        );

    \I__1367\ : Odrv12
    port map (
            O => \N__5963\,
            I => \D_UM_040_in_3\
        );

    \I__1366\ : IoInMux
    port map (
            O => \N__5960\,
            I => \N__5957\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__5957\,
            I => \N__5953\
        );

    \I__1364\ : InMux
    port map (
            O => \N__5956\,
            I => \N__5950\
        );

    \I__1363\ : Span4Mux_s3_h
    port map (
            O => \N__5953\,
            I => \N__5947\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__5950\,
            I => \N__5944\
        );

    \I__1361\ : Sp12to4
    port map (
            O => \N__5947\,
            I => \N__5941\
        );

    \I__1360\ : Span12Mux_v
    port map (
            O => \N__5944\,
            I => \N__5938\
        );

    \I__1359\ : Span12Mux_v
    port map (
            O => \N__5941\,
            I => \N__5935\
        );

    \I__1358\ : Span12Mux_v
    port map (
            O => \N__5938\,
            I => \N__5930\
        );

    \I__1357\ : Span12Mux_h
    port map (
            O => \N__5935\,
            I => \N__5930\
        );

    \I__1356\ : Span12Mux_h
    port map (
            O => \N__5930\,
            I => \N__5927\
        );

    \I__1355\ : Odrv12
    port map (
            O => \N__5927\,
            I => \D_LL_040_in_3\
        );

    \I__1354\ : IoInMux
    port map (
            O => \N__5924\,
            I => \N__5921\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__5921\,
            I => \N__5918\
        );

    \I__1352\ : Span4Mux_s3_h
    port map (
            O => \N__5918\,
            I => \N__5915\
        );

    \I__1351\ : Span4Mux_h
    port map (
            O => \N__5915\,
            I => \N__5912\
        );

    \I__1350\ : Span4Mux_h
    port map (
            O => \N__5912\,
            I => \N__5909\
        );

    \I__1349\ : Span4Mux_h
    port map (
            O => \N__5909\,
            I => \N__5906\
        );

    \I__1348\ : Odrv4
    port map (
            O => \N__5906\,
            I => \un1_D_UM_040_3\
        );

    \I__1347\ : InMux
    port map (
            O => \N__5903\,
            I => \N__5899\
        );

    \I__1346\ : InMux
    port map (
            O => \N__5902\,
            I => \N__5896\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__5899\,
            I => \N__5893\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__5896\,
            I => \N__5889\
        );

    \I__1343\ : Span4Mux_h
    port map (
            O => \N__5893\,
            I => \N__5886\
        );

    \I__1342\ : InMux
    port map (
            O => \N__5892\,
            I => \N__5883\
        );

    \I__1341\ : Span4Mux_v
    port map (
            O => \N__5889\,
            I => \N__5880\
        );

    \I__1340\ : Span4Mux_v
    port map (
            O => \N__5886\,
            I => \N__5875\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__5883\,
            I => \N__5875\
        );

    \I__1338\ : Sp12to4
    port map (
            O => \N__5880\,
            I => \N__5872\
        );

    \I__1337\ : Span4Mux_v
    port map (
            O => \N__5875\,
            I => \N__5869\
        );

    \I__1336\ : Span12Mux_h
    port map (
            O => \N__5872\,
            I => \N__5866\
        );

    \I__1335\ : Sp12to4
    port map (
            O => \N__5869\,
            I => \N__5863\
        );

    \I__1334\ : Span12Mux_v
    port map (
            O => \N__5866\,
            I => \N__5858\
        );

    \I__1333\ : Span12Mux_h
    port map (
            O => \N__5863\,
            I => \N__5858\
        );

    \I__1332\ : Odrv12
    port map (
            O => \N__5858\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__1331\ : InMux
    port map (
            O => \N__5855\,
            I => \N__5852\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__5852\,
            I => \N__5849\
        );

    \I__1329\ : Span4Mux_v
    port map (
            O => \N__5849\,
            I => \N__5846\
        );

    \I__1328\ : Odrv4
    port map (
            O => \N__5846\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\
        );

    \I__1327\ : IoInMux
    port map (
            O => \N__5843\,
            I => \N__5840\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__5840\,
            I => \N__5837\
        );

    \I__1325\ : IoSpan4Mux
    port map (
            O => \N__5837\,
            I => \N__5834\
        );

    \I__1324\ : Span4Mux_s3_h
    port map (
            O => \N__5834\,
            I => \N__5831\
        );

    \I__1323\ : Span4Mux_h
    port map (
            O => \N__5831\,
            I => \N__5828\
        );

    \I__1322\ : Span4Mux_h
    port map (
            O => \N__5828\,
            I => \N__5825\
        );

    \I__1321\ : Span4Mux_h
    port map (
            O => \N__5825\,
            I => \N__5822\
        );

    \I__1320\ : Odrv4
    port map (
            O => \N__5822\,
            I => \un1_D_UM_AMIGA_7\
        );

    \I__1319\ : InMux
    port map (
            O => \N__5819\,
            I => \N__5816\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__5816\,
            I => \N__5813\
        );

    \I__1317\ : Span4Mux_h
    port map (
            O => \N__5813\,
            I => \N__5810\
        );

    \I__1316\ : Sp12to4
    port map (
            O => \N__5810\,
            I => \N__5807\
        );

    \I__1315\ : Span12Mux_v
    port map (
            O => \N__5807\,
            I => \N__5804\
        );

    \I__1314\ : Span12Mux_h
    port map (
            O => \N__5804\,
            I => \N__5801\
        );

    \I__1313\ : Odrv12
    port map (
            O => \N__5801\,
            I => \D_UM_040_in_4\
        );

    \I__1312\ : InMux
    port map (
            O => \N__5798\,
            I => \N__5794\
        );

    \I__1311\ : IoInMux
    port map (
            O => \N__5797\,
            I => \N__5791\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__5794\,
            I => \N__5788\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__5791\,
            I => \N__5785\
        );

    \I__1308\ : Span4Mux_v
    port map (
            O => \N__5788\,
            I => \N__5782\
        );

    \I__1307\ : Span4Mux_s2_h
    port map (
            O => \N__5785\,
            I => \N__5779\
        );

    \I__1306\ : Sp12to4
    port map (
            O => \N__5782\,
            I => \N__5776\
        );

    \I__1305\ : Span4Mux_v
    port map (
            O => \N__5779\,
            I => \N__5773\
        );

    \I__1304\ : Span12Mux_h
    port map (
            O => \N__5776\,
            I => \N__5770\
        );

    \I__1303\ : Sp12to4
    port map (
            O => \N__5773\,
            I => \N__5767\
        );

    \I__1302\ : Span12Mux_v
    port map (
            O => \N__5770\,
            I => \N__5764\
        );

    \I__1301\ : Span12Mux_h
    port map (
            O => \N__5767\,
            I => \N__5761\
        );

    \I__1300\ : Span12Mux_v
    port map (
            O => \N__5764\,
            I => \N__5756\
        );

    \I__1299\ : Span12Mux_h
    port map (
            O => \N__5761\,
            I => \N__5756\
        );

    \I__1298\ : Odrv12
    port map (
            O => \N__5756\,
            I => \D_LL_040_in_4\
        );

    \I__1297\ : IoInMux
    port map (
            O => \N__5753\,
            I => \N__5750\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__5750\,
            I => \N__5747\
        );

    \I__1295\ : Span4Mux_s3_h
    port map (
            O => \N__5747\,
            I => \N__5744\
        );

    \I__1294\ : Span4Mux_h
    port map (
            O => \N__5744\,
            I => \N__5741\
        );

    \I__1293\ : Span4Mux_h
    port map (
            O => \N__5741\,
            I => \N__5738\
        );

    \I__1292\ : Span4Mux_h
    port map (
            O => \N__5738\,
            I => \N__5735\
        );

    \I__1291\ : Odrv4
    port map (
            O => \N__5735\,
            I => \un1_D_UM_040_4\
        );

    \I__1290\ : InMux
    port map (
            O => \N__5732\,
            I => \N__5729\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__5729\,
            I => \N__5726\
        );

    \I__1288\ : Span4Mux_v
    port map (
            O => \N__5726\,
            I => \N__5723\
        );

    \I__1287\ : Span4Mux_v
    port map (
            O => \N__5723\,
            I => \N__5720\
        );

    \I__1286\ : Sp12to4
    port map (
            O => \N__5720\,
            I => \N__5717\
        );

    \I__1285\ : Span12Mux_h
    port map (
            O => \N__5717\,
            I => \N__5714\
        );

    \I__1284\ : Odrv12
    port map (
            O => \N__5714\,
            I => \D_UM_040_in_7\
        );

    \I__1283\ : IoInMux
    port map (
            O => \N__5711\,
            I => \N__5708\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__5708\,
            I => \N__5705\
        );

    \I__1281\ : IoSpan4Mux
    port map (
            O => \N__5705\,
            I => \N__5702\
        );

    \I__1280\ : Span4Mux_s3_h
    port map (
            O => \N__5702\,
            I => \N__5698\
        );

    \I__1279\ : InMux
    port map (
            O => \N__5701\,
            I => \N__5695\
        );

    \I__1278\ : Sp12to4
    port map (
            O => \N__5698\,
            I => \N__5692\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__5695\,
            I => \N__5689\
        );

    \I__1276\ : Span12Mux_v
    port map (
            O => \N__5692\,
            I => \N__5686\
        );

    \I__1275\ : Span12Mux_v
    port map (
            O => \N__5689\,
            I => \N__5683\
        );

    \I__1274\ : Span12Mux_h
    port map (
            O => \N__5686\,
            I => \N__5678\
        );

    \I__1273\ : Span12Mux_v
    port map (
            O => \N__5683\,
            I => \N__5678\
        );

    \I__1272\ : Span12Mux_h
    port map (
            O => \N__5678\,
            I => \N__5675\
        );

    \I__1271\ : Odrv12
    port map (
            O => \N__5675\,
            I => \D_LL_040_in_7\
        );

    \I__1270\ : IoInMux
    port map (
            O => \N__5672\,
            I => \N__5669\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__5669\,
            I => \N__5666\
        );

    \I__1268\ : Span12Mux_s3_h
    port map (
            O => \N__5666\,
            I => \N__5663\
        );

    \I__1267\ : Span12Mux_h
    port map (
            O => \N__5663\,
            I => \N__5660\
        );

    \I__1266\ : Odrv12
    port map (
            O => \N__5660\,
            I => \un1_D_UM_040_7\
        );

    \I__1265\ : InMux
    port map (
            O => \N__5657\,
            I => \N__5651\
        );

    \I__1264\ : InMux
    port map (
            O => \N__5656\,
            I => \N__5648\
        );

    \I__1263\ : InMux
    port map (
            O => \N__5655\,
            I => \N__5645\
        );

    \I__1262\ : InMux
    port map (
            O => \N__5654\,
            I => \N__5642\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__5651\,
            I => \N__5628\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__5648\,
            I => \N__5628\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__5645\,
            I => \N__5628\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__5642\,
            I => \N__5628\
        );

    \I__1257\ : InMux
    port map (
            O => \N__5641\,
            I => \N__5625\
        );

    \I__1256\ : InMux
    port map (
            O => \N__5640\,
            I => \N__5620\
        );

    \I__1255\ : InMux
    port map (
            O => \N__5639\,
            I => \N__5620\
        );

    \I__1254\ : InMux
    port map (
            O => \N__5638\,
            I => \N__5615\
        );

    \I__1253\ : InMux
    port map (
            O => \N__5637\,
            I => \N__5615\
        );

    \I__1252\ : Span4Mux_v
    port map (
            O => \N__5628\,
            I => \N__5606\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__5625\,
            I => \N__5606\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__5620\,
            I => \N__5606\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__5615\,
            I => \N__5606\
        );

    \I__1248\ : Span4Mux_v
    port map (
            O => \N__5606\,
            I => \N__5603\
        );

    \I__1247\ : Span4Mux_h
    port map (
            O => \N__5603\,
            I => \N__5600\
        );

    \I__1246\ : Sp12to4
    port map (
            O => \N__5600\,
            I => \N__5597\
        );

    \I__1245\ : Span12Mux_v
    port map (
            O => \N__5597\,
            I => \N__5594\
        );

    \I__1244\ : Odrv12
    port map (
            O => \N__5594\,
            I => \RESETn_c\
        );

    \I__1243\ : CascadeMux
    port map (
            O => \N__5591\,
            I => \U111_CYCLE_SM.CYCLE_STATE_srsts_i_1_2_cascade_\
        );

    \I__1242\ : InMux
    port map (
            O => \N__5588\,
            I => \N__5585\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__5585\,
            I => \N__5582\
        );

    \I__1240\ : Glb2LocalMux
    port map (
            O => \N__5582\,
            I => \N__5579\
        );

    \I__1239\ : GlobalMux
    port map (
            O => \N__5579\,
            I => \CLK80\
        );

    \I__1238\ : IoInMux
    port map (
            O => \N__5576\,
            I => \N__5573\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__5573\,
            I => \N__5569\
        );

    \I__1236\ : IoInMux
    port map (
            O => \N__5572\,
            I => \N__5566\
        );

    \I__1235\ : Span4Mux_s1_v
    port map (
            O => \N__5569\,
            I => \N__5563\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__5566\,
            I => \N__5560\
        );

    \I__1233\ : Span4Mux_v
    port map (
            O => \N__5563\,
            I => \N__5557\
        );

    \I__1232\ : IoSpan4Mux
    port map (
            O => \N__5560\,
            I => \N__5554\
        );

    \I__1231\ : Span4Mux_v
    port map (
            O => \N__5557\,
            I => \N__5551\
        );

    \I__1230\ : Span4Mux_s3_h
    port map (
            O => \N__5554\,
            I => \N__5548\
        );

    \I__1229\ : Span4Mux_v
    port map (
            O => \N__5551\,
            I => \N__5545\
        );

    \I__1228\ : Sp12to4
    port map (
            O => \N__5548\,
            I => \N__5542\
        );

    \I__1227\ : Odrv4
    port map (
            O => \N__5545\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__1226\ : Odrv12
    port map (
            O => \N__5542\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__1225\ : InMux
    port map (
            O => \N__5537\,
            I => \N__5534\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__5534\,
            I => \N__5531\
        );

    \I__1223\ : Span12Mux_h
    port map (
            O => \N__5531\,
            I => \N__5528\
        );

    \I__1222\ : Odrv12
    port map (
            O => \N__5528\,
            I => \D_LM_AMIGA_in_2\
        );

    \I__1221\ : InMux
    port map (
            O => \N__5525\,
            I => \N__5521\
        );

    \I__1220\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5518\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__5521\,
            I => \N__5515\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__5518\,
            I => \N__5512\
        );

    \I__1217\ : Span4Mux_v
    port map (
            O => \N__5515\,
            I => \N__5508\
        );

    \I__1216\ : Span4Mux_v
    port map (
            O => \N__5512\,
            I => \N__5505\
        );

    \I__1215\ : InMux
    port map (
            O => \N__5511\,
            I => \N__5502\
        );

    \I__1214\ : Span4Mux_v
    port map (
            O => \N__5508\,
            I => \N__5499\
        );

    \I__1213\ : Span4Mux_v
    port map (
            O => \N__5505\,
            I => \N__5494\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__5502\,
            I => \N__5494\
        );

    \I__1211\ : Span4Mux_v
    port map (
            O => \N__5499\,
            I => \N__5491\
        );

    \I__1210\ : Span4Mux_v
    port map (
            O => \N__5494\,
            I => \N__5488\
        );

    \I__1209\ : Sp12to4
    port map (
            O => \N__5491\,
            I => \N__5483\
        );

    \I__1208\ : Sp12to4
    port map (
            O => \N__5488\,
            I => \N__5483\
        );

    \I__1207\ : Span12Mux_h
    port map (
            O => \N__5483\,
            I => \N__5480\
        );

    \I__1206\ : Odrv12
    port map (
            O => \N__5480\,
            I => \D_UU_AMIGA_in_2\
        );

    \I__1205\ : IoInMux
    port map (
            O => \N__5477\,
            I => \N__5474\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__5474\,
            I => \N__5471\
        );

    \I__1203\ : Span12Mux_s7_h
    port map (
            O => \N__5471\,
            I => \N__5468\
        );

    \I__1202\ : Span12Mux_v
    port map (
            O => \N__5468\,
            I => \N__5465\
        );

    \I__1201\ : Odrv12
    port map (
            O => \N__5465\,
            I => \un1_D_LM_AMIGA_2\
        );

    \I__1200\ : CascadeMux
    port map (
            O => \N__5462\,
            I => \N__5458\
        );

    \I__1199\ : InMux
    port map (
            O => \N__5461\,
            I => \N__5453\
        );

    \I__1198\ : InMux
    port map (
            O => \N__5458\,
            I => \N__5453\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__5453\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\
        );

    \I__1196\ : CascadeMux
    port map (
            O => \N__5450\,
            I => \U111_CYCLE_SM.CYCLE_STATE_srsts_i_o2_0_5_cascade_\
        );

    \I__1195\ : InMux
    port map (
            O => \N__5447\,
            I => \N__5443\
        );

    \I__1194\ : InMux
    port map (
            O => \N__5446\,
            I => \N__5439\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__5443\,
            I => \N__5436\
        );

    \I__1192\ : InMux
    port map (
            O => \N__5442\,
            I => \N__5433\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__5439\,
            I => \N__5429\
        );

    \I__1190\ : Span4Mux_h
    port map (
            O => \N__5436\,
            I => \N__5423\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5433\,
            I => \N__5423\
        );

    \I__1188\ : InMux
    port map (
            O => \N__5432\,
            I => \N__5420\
        );

    \I__1187\ : Span4Mux_v
    port map (
            O => \N__5429\,
            I => \N__5417\
        );

    \I__1186\ : InMux
    port map (
            O => \N__5428\,
            I => \N__5414\
        );

    \I__1185\ : Sp12to4
    port map (
            O => \N__5423\,
            I => \N__5409\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__5420\,
            I => \N__5409\
        );

    \I__1183\ : Span4Mux_v
    port map (
            O => \N__5417\,
            I => \N__5404\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__5414\,
            I => \N__5404\
        );

    \I__1181\ : Span12Mux_v
    port map (
            O => \N__5409\,
            I => \N__5401\
        );

    \I__1180\ : Span4Mux_v
    port map (
            O => \N__5404\,
            I => \N__5398\
        );

    \I__1179\ : Odrv12
    port map (
            O => \N__5401\,
            I => \LBENn_c\
        );

    \I__1178\ : Odrv4
    port map (
            O => \N__5398\,
            I => \LBENn_c\
        );

    \I__1177\ : InMux
    port map (
            O => \N__5393\,
            I => \N__5390\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__5390\,
            I => \N__5386\
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__5389\,
            I => \N__5383\
        );

    \I__1174\ : Span4Mux_h
    port map (
            O => \N__5386\,
            I => \N__5380\
        );

    \I__1173\ : InMux
    port map (
            O => \N__5383\,
            I => \N__5377\
        );

    \I__1172\ : Odrv4
    port map (
            O => \N__5380\,
            I => \U111_CYCLE_SM.TA_DISZ0\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__5377\,
            I => \U111_CYCLE_SM.TA_DISZ0\
        );

    \I__1170\ : IoInMux
    port map (
            O => \N__5372\,
            I => \N__5369\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__5369\,
            I => \N__5366\
        );

    \I__1168\ : Span4Mux_s3_v
    port map (
            O => \N__5366\,
            I => \N__5363\
        );

    \I__1167\ : Span4Mux_v
    port map (
            O => \N__5363\,
            I => \N__5360\
        );

    \I__1166\ : Span4Mux_v
    port map (
            O => \N__5360\,
            I => \N__5357\
        );

    \I__1165\ : Span4Mux_v
    port map (
            O => \N__5357\,
            I => \N__5354\
        );

    \I__1164\ : Odrv4
    port map (
            O => \N__5354\,
            I => \TAn_1_i\
        );

    \I__1163\ : InMux
    port map (
            O => \N__5351\,
            I => \N__5342\
        );

    \I__1162\ : InMux
    port map (
            O => \N__5350\,
            I => \N__5342\
        );

    \I__1161\ : InMux
    port map (
            O => \N__5349\,
            I => \N__5339\
        );

    \I__1160\ : InMux
    port map (
            O => \N__5348\,
            I => \N__5334\
        );

    \I__1159\ : InMux
    port map (
            O => \N__5347\,
            I => \N__5334\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__5342\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__5339\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__5334\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__5327\,
            I => \U111_CYCLE_SM.N_135_cascade_\
        );

    \I__1154\ : InMux
    port map (
            O => \N__5324\,
            I => \N__5321\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__5321\,
            I => \U111_CYCLE_SM.N_128_0\
        );

    \I__1152\ : CascadeMux
    port map (
            O => \N__5318\,
            I => \U111_CYCLE_SM.CYCLE_STATE_srsts_0_1_0_cascade_\
        );

    \I__1151\ : InMux
    port map (
            O => \N__5315\,
            I => \N__5310\
        );

    \I__1150\ : InMux
    port map (
            O => \N__5314\,
            I => \N__5307\
        );

    \I__1149\ : InMux
    port map (
            O => \N__5313\,
            I => \N__5301\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__5310\,
            I => \N__5298\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__5307\,
            I => \N__5295\
        );

    \I__1146\ : InMux
    port map (
            O => \N__5306\,
            I => \N__5292\
        );

    \I__1145\ : InMux
    port map (
            O => \N__5305\,
            I => \N__5287\
        );

    \I__1144\ : InMux
    port map (
            O => \N__5304\,
            I => \N__5287\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__5301\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1142\ : Odrv4
    port map (
            O => \N__5298\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1141\ : Odrv4
    port map (
            O => \N__5295\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__5292\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__5287\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1138\ : IoInMux
    port map (
            O => \N__5276\,
            I => \N__5273\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__5273\,
            I => \N__5270\
        );

    \I__1136\ : Span4Mux_s1_v
    port map (
            O => \N__5270\,
            I => \N__5261\
        );

    \I__1135\ : InMux
    port map (
            O => \N__5269\,
            I => \N__5256\
        );

    \I__1134\ : InMux
    port map (
            O => \N__5268\,
            I => \N__5256\
        );

    \I__1133\ : InMux
    port map (
            O => \N__5267\,
            I => \N__5253\
        );

    \I__1132\ : InMux
    port map (
            O => \N__5266\,
            I => \N__5250\
        );

    \I__1131\ : InMux
    port map (
            O => \N__5265\,
            I => \N__5245\
        );

    \I__1130\ : InMux
    port map (
            O => \N__5264\,
            I => \N__5245\
        );

    \I__1129\ : Span4Mux_v
    port map (
            O => \N__5261\,
            I => \N__5242\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__5256\,
            I => \N__5239\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__5253\,
            I => \N__5232\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__5250\,
            I => \N__5232\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__5245\,
            I => \N__5232\
        );

    \I__1124\ : Sp12to4
    port map (
            O => \N__5242\,
            I => \N__5229\
        );

    \I__1123\ : Span4Mux_v
    port map (
            O => \N__5239\,
            I => \N__5226\
        );

    \I__1122\ : Span4Mux_v
    port map (
            O => \N__5232\,
            I => \N__5223\
        );

    \I__1121\ : Span12Mux_h
    port map (
            O => \N__5229\,
            I => \N__5220\
        );

    \I__1120\ : Sp12to4
    port map (
            O => \N__5226\,
            I => \N__5215\
        );

    \I__1119\ : Sp12to4
    port map (
            O => \N__5223\,
            I => \N__5215\
        );

    \I__1118\ : Span12Mux_v
    port map (
            O => \N__5220\,
            I => \N__5210\
        );

    \I__1117\ : Span12Mux_h
    port map (
            O => \N__5215\,
            I => \N__5210\
        );

    \I__1116\ : Span12Mux_v
    port map (
            O => \N__5210\,
            I => \N__5207\
        );

    \I__1115\ : Odrv12
    port map (
            O => \N__5207\,
            I => \TEAn_c\
        );

    \I__1114\ : InMux
    port map (
            O => \N__5204\,
            I => \N__5201\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__5201\,
            I => \N__5198\
        );

    \I__1112\ : Span4Mux_v
    port map (
            O => \N__5198\,
            I => \N__5195\
        );

    \I__1111\ : Odrv4
    port map (
            O => \N__5195\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\
        );

    \I__1110\ : InMux
    port map (
            O => \N__5192\,
            I => \N__5188\
        );

    \I__1109\ : InMux
    port map (
            O => \N__5191\,
            I => \N__5185\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__5188\,
            I => \N__5182\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__5185\,
            I => \N__5178\
        );

    \I__1106\ : Span4Mux_v
    port map (
            O => \N__5182\,
            I => \N__5175\
        );

    \I__1105\ : InMux
    port map (
            O => \N__5181\,
            I => \N__5172\
        );

    \I__1104\ : Span4Mux_v
    port map (
            O => \N__5178\,
            I => \N__5169\
        );

    \I__1103\ : Sp12to4
    port map (
            O => \N__5175\,
            I => \N__5164\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__5172\,
            I => \N__5164\
        );

    \I__1101\ : Sp12to4
    port map (
            O => \N__5169\,
            I => \N__5161\
        );

    \I__1100\ : Span12Mux_h
    port map (
            O => \N__5164\,
            I => \N__5158\
        );

    \I__1099\ : Span12Mux_h
    port map (
            O => \N__5161\,
            I => \N__5155\
        );

    \I__1098\ : Odrv12
    port map (
            O => \N__5158\,
            I => \D_UU_AMIGA_in_7\
        );

    \I__1097\ : Odrv12
    port map (
            O => \N__5155\,
            I => \D_UU_AMIGA_in_7\
        );

    \I__1096\ : IoInMux
    port map (
            O => \N__5150\,
            I => \N__5147\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__5147\,
            I => \N__5144\
        );

    \I__1094\ : IoSpan4Mux
    port map (
            O => \N__5144\,
            I => \N__5141\
        );

    \I__1093\ : Span4Mux_s2_v
    port map (
            O => \N__5141\,
            I => \N__5138\
        );

    \I__1092\ : Span4Mux_v
    port map (
            O => \N__5138\,
            I => \N__5135\
        );

    \I__1091\ : Sp12to4
    port map (
            O => \N__5135\,
            I => \N__5132\
        );

    \I__1090\ : Odrv12
    port map (
            O => \N__5132\,
            I => \un1_D_UU_AMIGA_7\
        );

    \I__1089\ : InMux
    port map (
            O => \N__5129\,
            I => \N__5126\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__5126\,
            I => \N__5123\
        );

    \I__1087\ : Span4Mux_v
    port map (
            O => \N__5123\,
            I => \N__5120\
        );

    \I__1086\ : Sp12to4
    port map (
            O => \N__5120\,
            I => \N__5117\
        );

    \I__1085\ : Span12Mux_h
    port map (
            O => \N__5117\,
            I => \N__5114\
        );

    \I__1084\ : Odrv12
    port map (
            O => \N__5114\,
            I => \D_LL_AMIGA_in_2\
        );

    \I__1083\ : IoInMux
    port map (
            O => \N__5111\,
            I => \N__5108\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__5108\,
            I => \N__5105\
        );

    \I__1081\ : Span4Mux_s3_h
    port map (
            O => \N__5105\,
            I => \N__5102\
        );

    \I__1080\ : Span4Mux_v
    port map (
            O => \N__5102\,
            I => \N__5099\
        );

    \I__1079\ : Span4Mux_h
    port map (
            O => \N__5099\,
            I => \N__5096\
        );

    \I__1078\ : Span4Mux_h
    port map (
            O => \N__5096\,
            I => \N__5093\
        );

    \I__1077\ : Span4Mux_h
    port map (
            O => \N__5093\,
            I => \N__5090\
        );

    \I__1076\ : Odrv4
    port map (
            O => \N__5090\,
            I => \un1_D_LL_AMIGA_2\
        );

    \I__1075\ : InMux
    port map (
            O => \N__5087\,
            I => \N__5084\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__5084\,
            I => \N__5081\
        );

    \I__1073\ : Span12Mux_v
    port map (
            O => \N__5081\,
            I => \N__5078\
        );

    \I__1072\ : Span12Mux_h
    port map (
            O => \N__5078\,
            I => \N__5075\
        );

    \I__1071\ : Odrv12
    port map (
            O => \N__5075\,
            I => \D_LL_AMIGA_in_4\
        );

    \I__1070\ : IoInMux
    port map (
            O => \N__5072\,
            I => \N__5069\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__5069\,
            I => \N__5066\
        );

    \I__1068\ : Span4Mux_s3_h
    port map (
            O => \N__5066\,
            I => \N__5063\
        );

    \I__1067\ : Span4Mux_h
    port map (
            O => \N__5063\,
            I => \N__5060\
        );

    \I__1066\ : Sp12to4
    port map (
            O => \N__5060\,
            I => \N__5057\
        );

    \I__1065\ : Span12Mux_s8_v
    port map (
            O => \N__5057\,
            I => \N__5054\
        );

    \I__1064\ : Odrv12
    port map (
            O => \N__5054\,
            I => \un1_D_LL_AMIGA_4\
        );

    \I__1063\ : InMux
    port map (
            O => \N__5051\,
            I => \N__5045\
        );

    \I__1062\ : InMux
    port map (
            O => \N__5050\,
            I => \N__5045\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__5045\,
            I => \N__5042\
        );

    \I__1060\ : Span4Mux_v
    port map (
            O => \N__5042\,
            I => \N__5039\
        );

    \I__1059\ : Sp12to4
    port map (
            O => \N__5039\,
            I => \N__5036\
        );

    \I__1058\ : Span12Mux_h
    port map (
            O => \N__5036\,
            I => \N__5032\
        );

    \I__1057\ : InMux
    port map (
            O => \N__5035\,
            I => \N__5029\
        );

    \I__1056\ : Odrv12
    port map (
            O => \N__5032\,
            I => \U111_CYCLE_SM.A2_ENZ0\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__5029\,
            I => \U111_CYCLE_SM.A2_ENZ0\
        );

    \I__1054\ : InMux
    port map (
            O => \N__5024\,
            I => \N__5021\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__5021\,
            I => \U111_CYCLE_SM.N_148\
        );

    \I__1052\ : CascadeMux
    port map (
            O => \N__5018\,
            I => \U111_CYCLE_SM.N_148_cascade_\
        );

    \I__1051\ : InMux
    port map (
            O => \N__5015\,
            I => \N__5012\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__5012\,
            I => \U111_CYCLE_SM.TS_EN_6\
        );

    \I__1049\ : InMux
    port map (
            O => \N__5009\,
            I => \N__5006\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__5006\,
            I => \N__5003\
        );

    \I__1047\ : Odrv4
    port map (
            O => \N__5003\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\
        );

    \I__1046\ : InMux
    port map (
            O => \N__5000\,
            I => \N__4995\
        );

    \I__1045\ : InMux
    port map (
            O => \N__4999\,
            I => \N__4992\
        );

    \I__1044\ : InMux
    port map (
            O => \N__4998\,
            I => \N__4989\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__4995\,
            I => \N__4984\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__4992\,
            I => \N__4984\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__4989\,
            I => \N__4981\
        );

    \I__1040\ : Span4Mux_v
    port map (
            O => \N__4984\,
            I => \N__4978\
        );

    \I__1039\ : Span4Mux_v
    port map (
            O => \N__4981\,
            I => \N__4975\
        );

    \I__1038\ : Sp12to4
    port map (
            O => \N__4978\,
            I => \N__4970\
        );

    \I__1037\ : Sp12to4
    port map (
            O => \N__4975\,
            I => \N__4970\
        );

    \I__1036\ : Span12Mux_h
    port map (
            O => \N__4970\,
            I => \N__4967\
        );

    \I__1035\ : Odrv12
    port map (
            O => \N__4967\,
            I => \D_UU_AMIGA_in_6\
        );

    \I__1034\ : IoInMux
    port map (
            O => \N__4964\,
            I => \N__4961\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__4961\,
            I => \N__4958\
        );

    \I__1032\ : Span4Mux_s3_v
    port map (
            O => \N__4958\,
            I => \N__4955\
        );

    \I__1031\ : Span4Mux_v
    port map (
            O => \N__4955\,
            I => \N__4952\
        );

    \I__1030\ : Sp12to4
    port map (
            O => \N__4952\,
            I => \N__4949\
        );

    \I__1029\ : Span12Mux_h
    port map (
            O => \N__4949\,
            I => \N__4946\
        );

    \I__1028\ : Odrv12
    port map (
            O => \N__4946\,
            I => \un1_D_UU_AMIGA_6\
        );

    \I__1027\ : InMux
    port map (
            O => \N__4943\,
            I => \N__4940\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__4940\,
            I => \N__4937\
        );

    \I__1025\ : Span4Mux_v
    port map (
            O => \N__4937\,
            I => \N__4932\
        );

    \I__1024\ : InMux
    port map (
            O => \N__4936\,
            I => \N__4929\
        );

    \I__1023\ : InMux
    port map (
            O => \N__4935\,
            I => \N__4926\
        );

    \I__1022\ : Span4Mux_v
    port map (
            O => \N__4932\,
            I => \N__4919\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__4929\,
            I => \N__4919\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__4926\,
            I => \N__4919\
        );

    \I__1019\ : Span4Mux_v
    port map (
            O => \N__4919\,
            I => \N__4916\
        );

    \I__1018\ : Sp12to4
    port map (
            O => \N__4916\,
            I => \N__4913\
        );

    \I__1017\ : Span12Mux_h
    port map (
            O => \N__4913\,
            I => \N__4910\
        );

    \I__1016\ : Odrv12
    port map (
            O => \N__4910\,
            I => \D_UU_AMIGA_in_0\
        );

    \I__1015\ : InMux
    port map (
            O => \N__4907\,
            I => \N__4904\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__4904\,
            I => \N__4901\
        );

    \I__1013\ : Odrv4
    port map (
            O => \N__4901\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\
        );

    \I__1012\ : IoInMux
    port map (
            O => \N__4898\,
            I => \N__4895\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__4895\,
            I => \N__4892\
        );

    \I__1010\ : Span4Mux_s2_v
    port map (
            O => \N__4892\,
            I => \N__4889\
        );

    \I__1009\ : Span4Mux_v
    port map (
            O => \N__4889\,
            I => \N__4886\
        );

    \I__1008\ : Span4Mux_v
    port map (
            O => \N__4886\,
            I => \N__4883\
        );

    \I__1007\ : Sp12to4
    port map (
            O => \N__4883\,
            I => \N__4880\
        );

    \I__1006\ : Odrv12
    port map (
            O => \N__4880\,
            I => \un1_D_UU_AMIGA_0\
        );

    \I__1005\ : InMux
    port map (
            O => \N__4877\,
            I => \N__4874\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__4874\,
            I => \N__4871\
        );

    \I__1003\ : Odrv12
    port map (
            O => \N__4871\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\
        );

    \I__1002\ : IoInMux
    port map (
            O => \N__4868\,
            I => \N__4865\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__4865\,
            I => \N__4862\
        );

    \I__1000\ : Span12Mux_s9_v
    port map (
            O => \N__4862\,
            I => \N__4859\
        );

    \I__999\ : Span12Mux_h
    port map (
            O => \N__4859\,
            I => \N__4856\
        );

    \I__998\ : Odrv12
    port map (
            O => \N__4856\,
            I => \un1_D_UU_AMIGA_2\
        );

    \I__997\ : InMux
    port map (
            O => \N__4853\,
            I => \N__4850\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__4850\,
            I => \N__4847\
        );

    \I__995\ : Odrv12
    port map (
            O => \N__4847\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\
        );

    \I__994\ : InMux
    port map (
            O => \N__4844\,
            I => \N__4841\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__4841\,
            I => \N__4838\
        );

    \I__992\ : Span4Mux_v
    port map (
            O => \N__4838\,
            I => \N__4834\
        );

    \I__991\ : InMux
    port map (
            O => \N__4837\,
            I => \N__4831\
        );

    \I__990\ : Span4Mux_v
    port map (
            O => \N__4834\,
            I => \N__4828\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__4831\,
            I => \N__4825\
        );

    \I__988\ : Span4Mux_v
    port map (
            O => \N__4828\,
            I => \N__4819\
        );

    \I__987\ : Span4Mux_v
    port map (
            O => \N__4825\,
            I => \N__4819\
        );

    \I__986\ : InMux
    port map (
            O => \N__4824\,
            I => \N__4816\
        );

    \I__985\ : Span4Mux_v
    port map (
            O => \N__4819\,
            I => \N__4811\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__4816\,
            I => \N__4811\
        );

    \I__983\ : Span4Mux_v
    port map (
            O => \N__4811\,
            I => \N__4808\
        );

    \I__982\ : IoSpan4Mux
    port map (
            O => \N__4808\,
            I => \N__4805\
        );

    \I__981\ : IoSpan4Mux
    port map (
            O => \N__4805\,
            I => \N__4802\
        );

    \I__980\ : IoSpan4Mux
    port map (
            O => \N__4802\,
            I => \N__4799\
        );

    \I__979\ : Odrv4
    port map (
            O => \N__4799\,
            I => \D_UM_AMIGA_in_5\
        );

    \I__978\ : IoInMux
    port map (
            O => \N__4796\,
            I => \N__4793\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__4793\,
            I => \N__4790\
        );

    \I__976\ : Span4Mux_s2_v
    port map (
            O => \N__4790\,
            I => \N__4787\
        );

    \I__975\ : Span4Mux_v
    port map (
            O => \N__4787\,
            I => \N__4784\
        );

    \I__974\ : Sp12to4
    port map (
            O => \N__4784\,
            I => \N__4781\
        );

    \I__973\ : Span12Mux_h
    port map (
            O => \N__4781\,
            I => \N__4778\
        );

    \I__972\ : Odrv12
    port map (
            O => \N__4778\,
            I => \un1_D_UM_AMIGA_5\
        );

    \I__971\ : InMux
    port map (
            O => \N__4775\,
            I => \N__4772\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__4772\,
            I => \U111_CYCLE_SM.PORT_MISMATCH_2\
        );

    \I__969\ : CascadeMux
    port map (
            O => \N__4769\,
            I => \U111_CYCLE_SM.N_123_0_cascade_\
        );

    \I__968\ : InMux
    port map (
            O => \N__4766\,
            I => \N__4763\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__4763\,
            I => \U111_CYCLE_SM.N_121_0\
        );

    \I__966\ : InMux
    port map (
            O => \N__4760\,
            I => \N__4754\
        );

    \I__965\ : InMux
    port map (
            O => \N__4759\,
            I => \N__4754\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__4754\,
            I => \U111_CYCLE_SM.un1_CYCLE_STATE_0\
        );

    \I__963\ : IoInMux
    port map (
            O => \N__4751\,
            I => \N__4747\
        );

    \I__962\ : IoInMux
    port map (
            O => \N__4750\,
            I => \N__4744\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__4747\,
            I => \N__4737\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4744\,
            I => \N__4737\
        );

    \I__959\ : IoInMux
    port map (
            O => \N__4743\,
            I => \N__4734\
        );

    \I__958\ : IoInMux
    port map (
            O => \N__4742\,
            I => \N__4731\
        );

    \I__957\ : IoSpan4Mux
    port map (
            O => \N__4737\,
            I => \N__4719\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__4734\,
            I => \N__4719\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__4731\,
            I => \N__4719\
        );

    \I__954\ : IoInMux
    port map (
            O => \N__4730\,
            I => \N__4716\
        );

    \I__953\ : IoInMux
    port map (
            O => \N__4729\,
            I => \N__4713\
        );

    \I__952\ : IoInMux
    port map (
            O => \N__4728\,
            I => \N__4710\
        );

    \I__951\ : IoInMux
    port map (
            O => \N__4727\,
            I => \N__4707\
        );

    \I__950\ : IoInMux
    port map (
            O => \N__4726\,
            I => \N__4704\
        );

    \I__949\ : IoSpan4Mux
    port map (
            O => \N__4719\,
            I => \N__4688\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__4716\,
            I => \N__4688\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4713\,
            I => \N__4688\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__4710\,
            I => \N__4688\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__4707\,
            I => \N__4688\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4704\,
            I => \N__4688\
        );

    \I__943\ : IoInMux
    port map (
            O => \N__4703\,
            I => \N__4685\
        );

    \I__942\ : IoInMux
    port map (
            O => \N__4702\,
            I => \N__4682\
        );

    \I__941\ : IoInMux
    port map (
            O => \N__4701\,
            I => \N__4679\
        );

    \I__940\ : IoSpan4Mux
    port map (
            O => \N__4688\,
            I => \N__4675\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__4685\,
            I => \N__4667\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4682\,
            I => \N__4667\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__4679\,
            I => \N__4667\
        );

    \I__936\ : IoInMux
    port map (
            O => \N__4678\,
            I => \N__4664\
        );

    \I__935\ : IoSpan4Mux
    port map (
            O => \N__4675\,
            I => \N__4654\
        );

    \I__934\ : IoInMux
    port map (
            O => \N__4674\,
            I => \N__4651\
        );

    \I__933\ : IoSpan4Mux
    port map (
            O => \N__4667\,
            I => \N__4643\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4664\,
            I => \N__4643\
        );

    \I__931\ : IoInMux
    port map (
            O => \N__4663\,
            I => \N__4640\
        );

    \I__930\ : IoInMux
    port map (
            O => \N__4662\,
            I => \N__4633\
        );

    \I__929\ : IoInMux
    port map (
            O => \N__4661\,
            I => \N__4630\
        );

    \I__928\ : IoInMux
    port map (
            O => \N__4660\,
            I => \N__4627\
        );

    \I__927\ : IoInMux
    port map (
            O => \N__4659\,
            I => \N__4624\
        );

    \I__926\ : IoInMux
    port map (
            O => \N__4658\,
            I => \N__4621\
        );

    \I__925\ : IoInMux
    port map (
            O => \N__4657\,
            I => \N__4618\
        );

    \I__924\ : IoSpan4Mux
    port map (
            O => \N__4654\,
            I => \N__4613\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__4651\,
            I => \N__4613\
        );

    \I__922\ : IoInMux
    port map (
            O => \N__4650\,
            I => \N__4610\
        );

    \I__921\ : IoInMux
    port map (
            O => \N__4649\,
            I => \N__4607\
        );

    \I__920\ : IoInMux
    port map (
            O => \N__4648\,
            I => \N__4604\
        );

    \I__919\ : IoSpan4Mux
    port map (
            O => \N__4643\,
            I => \N__4599\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__4640\,
            I => \N__4599\
        );

    \I__917\ : IoInMux
    port map (
            O => \N__4639\,
            I => \N__4596\
        );

    \I__916\ : IoInMux
    port map (
            O => \N__4638\,
            I => \N__4593\
        );

    \I__915\ : IoInMux
    port map (
            O => \N__4637\,
            I => \N__4589\
        );

    \I__914\ : IoInMux
    port map (
            O => \N__4636\,
            I => \N__4586\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__4633\,
            I => \N__4575\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__4630\,
            I => \N__4575\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__4627\,
            I => \N__4575\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__4624\,
            I => \N__4575\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__4621\,
            I => \N__4571\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__4618\,
            I => \N__4568\
        );

    \I__907\ : IoSpan4Mux
    port map (
            O => \N__4613\,
            I => \N__4559\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__4610\,
            I => \N__4559\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__4607\,
            I => \N__4559\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__4604\,
            I => \N__4559\
        );

    \I__903\ : IoSpan4Mux
    port map (
            O => \N__4599\,
            I => \N__4552\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__4596\,
            I => \N__4552\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__4593\,
            I => \N__4552\
        );

    \I__900\ : IoInMux
    port map (
            O => \N__4592\,
            I => \N__4549\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__4589\,
            I => \N__4544\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__4586\,
            I => \N__4544\
        );

    \I__897\ : IoInMux
    port map (
            O => \N__4585\,
            I => \N__4541\
        );

    \I__896\ : IoInMux
    port map (
            O => \N__4584\,
            I => \N__4538\
        );

    \I__895\ : IoSpan4Mux
    port map (
            O => \N__4575\,
            I => \N__4535\
        );

    \I__894\ : IoInMux
    port map (
            O => \N__4574\,
            I => \N__4532\
        );

    \I__893\ : Span4Mux_s2_v
    port map (
            O => \N__4571\,
            I => \N__4529\
        );

    \I__892\ : Span4Mux_s2_v
    port map (
            O => \N__4568\,
            I => \N__4526\
        );

    \I__891\ : IoSpan4Mux
    port map (
            O => \N__4559\,
            I => \N__4521\
        );

    \I__890\ : IoSpan4Mux
    port map (
            O => \N__4552\,
            I => \N__4521\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__4549\,
            I => \N__4518\
        );

    \I__888\ : Span12Mux_s5_h
    port map (
            O => \N__4544\,
            I => \N__4515\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__4541\,
            I => \N__4510\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__4538\,
            I => \N__4510\
        );

    \I__885\ : Span4Mux_s2_v
    port map (
            O => \N__4535\,
            I => \N__4507\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__4532\,
            I => \N__4504\
        );

    \I__883\ : Sp12to4
    port map (
            O => \N__4529\,
            I => \N__4499\
        );

    \I__882\ : Sp12to4
    port map (
            O => \N__4526\,
            I => \N__4499\
        );

    \I__881\ : Span4Mux_s2_h
    port map (
            O => \N__4521\,
            I => \N__4496\
        );

    \I__880\ : Span12Mux_s5_h
    port map (
            O => \N__4518\,
            I => \N__4493\
        );

    \I__879\ : Span12Mux_h
    port map (
            O => \N__4515\,
            I => \N__4490\
        );

    \I__878\ : Span12Mux_s5_h
    port map (
            O => \N__4510\,
            I => \N__4481\
        );

    \I__877\ : Sp12to4
    port map (
            O => \N__4507\,
            I => \N__4481\
        );

    \I__876\ : Span12Mux_s2_v
    port map (
            O => \N__4504\,
            I => \N__4481\
        );

    \I__875\ : Span12Mux_h
    port map (
            O => \N__4499\,
            I => \N__4481\
        );

    \I__874\ : Span4Mux_h
    port map (
            O => \N__4496\,
            I => \N__4478\
        );

    \I__873\ : Span12Mux_h
    port map (
            O => \N__4493\,
            I => \N__4475\
        );

    \I__872\ : Span12Mux_v
    port map (
            O => \N__4490\,
            I => \N__4468\
        );

    \I__871\ : Span12Mux_v
    port map (
            O => \N__4481\,
            I => \N__4468\
        );

    \I__870\ : Sp12to4
    port map (
            O => \N__4478\,
            I => \N__4468\
        );

    \I__869\ : Odrv12
    port map (
            O => \N__4475\,
            I => \D_UU_040_1_i\
        );

    \I__868\ : Odrv12
    port map (
            O => \N__4468\,
            I => \D_UU_040_1_i\
        );

    \I__867\ : InMux
    port map (
            O => \N__4463\,
            I => \N__4458\
        );

    \I__866\ : InMux
    port map (
            O => \N__4462\,
            I => \N__4452\
        );

    \I__865\ : InMux
    port map (
            O => \N__4461\,
            I => \N__4452\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__4458\,
            I => \N__4449\
        );

    \I__863\ : InMux
    port map (
            O => \N__4457\,
            I => \N__4446\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4452\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__861\ : Odrv4
    port map (
            O => \N__4449\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__4446\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__859\ : CascadeMux
    port map (
            O => \N__4439\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81_cascade_\
        );

    \I__858\ : InMux
    port map (
            O => \N__4436\,
            I => \N__4433\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__4433\,
            I => \N__4430\
        );

    \I__856\ : Span4Mux_v
    port map (
            O => \N__4430\,
            I => \N__4427\
        );

    \I__855\ : Sp12to4
    port map (
            O => \N__4427\,
            I => \N__4424\
        );

    \I__854\ : Span12Mux_h
    port map (
            O => \N__4424\,
            I => \N__4421\
        );

    \I__853\ : Odrv12
    port map (
            O => \N__4421\,
            I => \D_LM_AMIGA_in_0\
        );

    \I__852\ : IoInMux
    port map (
            O => \N__4418\,
            I => \N__4415\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__4415\,
            I => \N__4412\
        );

    \I__850\ : Span4Mux_s2_h
    port map (
            O => \N__4412\,
            I => \N__4409\
        );

    \I__849\ : Span4Mux_v
    port map (
            O => \N__4409\,
            I => \N__4406\
        );

    \I__848\ : Span4Mux_v
    port map (
            O => \N__4406\,
            I => \N__4403\
        );

    \I__847\ : Span4Mux_h
    port map (
            O => \N__4403\,
            I => \N__4400\
        );

    \I__846\ : Sp12to4
    port map (
            O => \N__4400\,
            I => \N__4397\
        );

    \I__845\ : Odrv12
    port map (
            O => \N__4397\,
            I => \un1_D_LM_AMIGA_0\
        );

    \I__844\ : IoInMux
    port map (
            O => \N__4394\,
            I => \N__4391\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__4391\,
            I => \N__4388\
        );

    \I__842\ : IoSpan4Mux
    port map (
            O => \N__4388\,
            I => \N__4385\
        );

    \I__841\ : Sp12to4
    port map (
            O => \N__4385\,
            I => \N__4382\
        );

    \I__840\ : Span12Mux_s7_v
    port map (
            O => \N__4382\,
            I => \N__4379\
        );

    \I__839\ : Odrv12
    port map (
            O => \N__4379\,
            I => \TSn_c\
        );

    \I__838\ : IoInMux
    port map (
            O => \N__4376\,
            I => \N__4369\
        );

    \I__837\ : IoInMux
    port map (
            O => \N__4375\,
            I => \N__4366\
        );

    \I__836\ : IoInMux
    port map (
            O => \N__4374\,
            I => \N__4363\
        );

    \I__835\ : IoInMux
    port map (
            O => \N__4373\,
            I => \N__4360\
        );

    \I__834\ : IoInMux
    port map (
            O => \N__4372\,
            I => \N__4357\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__4369\,
            I => \N__4342\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4366\,
            I => \N__4342\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__4363\,
            I => \N__4342\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__4360\,
            I => \N__4342\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__4357\,
            I => \N__4342\
        );

    \I__828\ : IoInMux
    port map (
            O => \N__4356\,
            I => \N__4333\
        );

    \I__827\ : IoInMux
    port map (
            O => \N__4355\,
            I => \N__4330\
        );

    \I__826\ : IoInMux
    port map (
            O => \N__4354\,
            I => \N__4327\
        );

    \I__825\ : IoInMux
    port map (
            O => \N__4353\,
            I => \N__4324\
        );

    \I__824\ : IoSpan4Mux
    port map (
            O => \N__4342\,
            I => \N__4317\
        );

    \I__823\ : IoInMux
    port map (
            O => \N__4341\,
            I => \N__4314\
        );

    \I__822\ : IoInMux
    port map (
            O => \N__4340\,
            I => \N__4311\
        );

    \I__821\ : IoInMux
    port map (
            O => \N__4339\,
            I => \N__4308\
        );

    \I__820\ : IoInMux
    port map (
            O => \N__4338\,
            I => \N__4305\
        );

    \I__819\ : IoInMux
    port map (
            O => \N__4337\,
            I => \N__4299\
        );

    \I__818\ : IoInMux
    port map (
            O => \N__4336\,
            I => \N__4296\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__4333\,
            I => \N__4287\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__4330\,
            I => \N__4287\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__4327\,
            I => \N__4287\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__4324\,
            I => \N__4287\
        );

    \I__813\ : IoInMux
    port map (
            O => \N__4323\,
            I => \N__4283\
        );

    \I__812\ : IoInMux
    port map (
            O => \N__4322\,
            I => \N__4280\
        );

    \I__811\ : IoInMux
    port map (
            O => \N__4321\,
            I => \N__4276\
        );

    \I__810\ : IoInMux
    port map (
            O => \N__4320\,
            I => \N__4273\
        );

    \I__809\ : IoSpan4Mux
    port map (
            O => \N__4317\,
            I => \N__4262\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__4314\,
            I => \N__4262\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__4311\,
            I => \N__4262\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__4308\,
            I => \N__4262\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__4305\,
            I => \N__4262\
        );

    \I__804\ : IoInMux
    port map (
            O => \N__4304\,
            I => \N__4259\
        );

    \I__803\ : IoInMux
    port map (
            O => \N__4303\,
            I => \N__4250\
        );

    \I__802\ : IoInMux
    port map (
            O => \N__4302\,
            I => \N__4247\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__4299\,
            I => \N__4240\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__4296\,
            I => \N__4240\
        );

    \I__799\ : IoSpan4Mux
    port map (
            O => \N__4287\,
            I => \N__4237\
        );

    \I__798\ : IoInMux
    port map (
            O => \N__4286\,
            I => \N__4234\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__4283\,
            I => \N__4229\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__4280\,
            I => \N__4229\
        );

    \I__795\ : IoInMux
    port map (
            O => \N__4279\,
            I => \N__4226\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__4276\,
            I => \N__4217\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__4273\,
            I => \N__4217\
        );

    \I__792\ : IoSpan4Mux
    port map (
            O => \N__4262\,
            I => \N__4217\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__4259\,
            I => \N__4217\
        );

    \I__790\ : IoInMux
    port map (
            O => \N__4258\,
            I => \N__4214\
        );

    \I__789\ : IoInMux
    port map (
            O => \N__4257\,
            I => \N__4211\
        );

    \I__788\ : IoInMux
    port map (
            O => \N__4256\,
            I => \N__4208\
        );

    \I__787\ : IoInMux
    port map (
            O => \N__4255\,
            I => \N__4205\
        );

    \I__786\ : IoInMux
    port map (
            O => \N__4254\,
            I => \N__4202\
        );

    \I__785\ : IoInMux
    port map (
            O => \N__4253\,
            I => \N__4199\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__4250\,
            I => \N__4196\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__4247\,
            I => \N__4193\
        );

    \I__782\ : IoInMux
    port map (
            O => \N__4246\,
            I => \N__4190\
        );

    \I__781\ : IoInMux
    port map (
            O => \N__4245\,
            I => \N__4187\
        );

    \I__780\ : Span4Mux_s3_h
    port map (
            O => \N__4240\,
            I => \N__4182\
        );

    \I__779\ : Span4Mux_s2_v
    port map (
            O => \N__4237\,
            I => \N__4182\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__4234\,
            I => \N__4179\
        );

    \I__777\ : IoSpan4Mux
    port map (
            O => \N__4229\,
            I => \N__4174\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__4226\,
            I => \N__4174\
        );

    \I__775\ : IoSpan4Mux
    port map (
            O => \N__4217\,
            I => \N__4171\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__4214\,
            I => \N__4166\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__4211\,
            I => \N__4166\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__4208\,
            I => \N__4163\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__4205\,
            I => \N__4160\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__4202\,
            I => \N__4155\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__4199\,
            I => \N__4155\
        );

    \I__768\ : Span4Mux_s3_h
    port map (
            O => \N__4196\,
            I => \N__4150\
        );

    \I__767\ : Span4Mux_s3_h
    port map (
            O => \N__4193\,
            I => \N__4150\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__4190\,
            I => \N__4145\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__4187\,
            I => \N__4145\
        );

    \I__764\ : Span4Mux_v
    port map (
            O => \N__4182\,
            I => \N__4142\
        );

    \I__763\ : Span4Mux_s3_h
    port map (
            O => \N__4179\,
            I => \N__4135\
        );

    \I__762\ : Span4Mux_s3_h
    port map (
            O => \N__4174\,
            I => \N__4135\
        );

    \I__761\ : Span4Mux_s3_h
    port map (
            O => \N__4171\,
            I => \N__4135\
        );

    \I__760\ : Span4Mux_s3_h
    port map (
            O => \N__4166\,
            I => \N__4130\
        );

    \I__759\ : Span4Mux_s3_h
    port map (
            O => \N__4163\,
            I => \N__4130\
        );

    \I__758\ : Span12Mux_s10_v
    port map (
            O => \N__4160\,
            I => \N__4127\
        );

    \I__757\ : Span12Mux_s5_v
    port map (
            O => \N__4155\,
            I => \N__4114\
        );

    \I__756\ : Sp12to4
    port map (
            O => \N__4150\,
            I => \N__4114\
        );

    \I__755\ : Span12Mux_s3_h
    port map (
            O => \N__4145\,
            I => \N__4114\
        );

    \I__754\ : Sp12to4
    port map (
            O => \N__4142\,
            I => \N__4114\
        );

    \I__753\ : Sp12to4
    port map (
            O => \N__4135\,
            I => \N__4114\
        );

    \I__752\ : Sp12to4
    port map (
            O => \N__4130\,
            I => \N__4114\
        );

    \I__751\ : Span12Mux_h
    port map (
            O => \N__4127\,
            I => \N__4111\
        );

    \I__750\ : Span12Mux_v
    port map (
            O => \N__4114\,
            I => \N__4108\
        );

    \I__749\ : Odrv12
    port map (
            O => \N__4111\,
            I => \D_UU_AMIGA_1_i\
        );

    \I__748\ : Odrv12
    port map (
            O => \N__4108\,
            I => \D_UU_AMIGA_1_i\
        );

    \I__747\ : CascadeMux
    port map (
            O => \N__4103\,
            I => \N__4100\
        );

    \I__746\ : InMux
    port map (
            O => \N__4100\,
            I => \N__4097\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__4097\,
            I => \N__4093\
        );

    \I__744\ : InMux
    port map (
            O => \N__4096\,
            I => \N__4090\
        );

    \I__743\ : Odrv4
    port map (
            O => \N__4093\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__4090\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__741\ : CascadeMux
    port map (
            O => \N__4085\,
            I => \N__4082\
        );

    \I__740\ : InMux
    port map (
            O => \N__4082\,
            I => \N__4079\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__4079\,
            I => \N__4076\
        );

    \I__738\ : Odrv12
    port map (
            O => \N__4076\,
            I => \U111_CYCLE_SM.FLIP_WORD_2\
        );

    \I__737\ : InMux
    port map (
            O => \N__4073\,
            I => \N__4070\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__4070\,
            I => \N__4067\
        );

    \I__735\ : Span4Mux_v
    port map (
            O => \N__4067\,
            I => \N__4064\
        );

    \I__734\ : Sp12to4
    port map (
            O => \N__4064\,
            I => \N__4061\
        );

    \I__733\ : Span12Mux_h
    port map (
            O => \N__4061\,
            I => \N__4058\
        );

    \I__732\ : Odrv12
    port map (
            O => \N__4058\,
            I => \D_UM_040_in_2\
        );

    \I__731\ : IoInMux
    port map (
            O => \N__4055\,
            I => \N__4052\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__4052\,
            I => \N__4048\
        );

    \I__729\ : InMux
    port map (
            O => \N__4051\,
            I => \N__4045\
        );

    \I__728\ : IoSpan4Mux
    port map (
            O => \N__4048\,
            I => \N__4042\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__4045\,
            I => \N__4039\
        );

    \I__726\ : Span4Mux_s2_h
    port map (
            O => \N__4042\,
            I => \N__4036\
        );

    \I__725\ : Span4Mux_v
    port map (
            O => \N__4039\,
            I => \N__4033\
        );

    \I__724\ : Sp12to4
    port map (
            O => \N__4036\,
            I => \N__4030\
        );

    \I__723\ : Sp12to4
    port map (
            O => \N__4033\,
            I => \N__4027\
        );

    \I__722\ : Span12Mux_h
    port map (
            O => \N__4030\,
            I => \N__4024\
        );

    \I__721\ : Span12Mux_h
    port map (
            O => \N__4027\,
            I => \N__4021\
        );

    \I__720\ : Span12Mux_h
    port map (
            O => \N__4024\,
            I => \N__4016\
        );

    \I__719\ : Span12Mux_v
    port map (
            O => \N__4021\,
            I => \N__4016\
        );

    \I__718\ : Odrv12
    port map (
            O => \N__4016\,
            I => \D_LL_040_in_2\
        );

    \I__717\ : IoInMux
    port map (
            O => \N__4013\,
            I => \N__4010\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__4010\,
            I => \N__4007\
        );

    \I__715\ : IoSpan4Mux
    port map (
            O => \N__4007\,
            I => \N__4004\
        );

    \I__714\ : Span4Mux_s1_h
    port map (
            O => \N__4004\,
            I => \N__4001\
        );

    \I__713\ : Sp12to4
    port map (
            O => \N__4001\,
            I => \N__3998\
        );

    \I__712\ : Span12Mux_s9_h
    port map (
            O => \N__3998\,
            I => \N__3995\
        );

    \I__711\ : Odrv12
    port map (
            O => \N__3995\,
            I => \un1_D_UM_040_2\
        );

    \I__710\ : IoInMux
    port map (
            O => \N__3992\,
            I => \N__3989\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__3989\,
            I => \N__3985\
        );

    \I__708\ : IoInMux
    port map (
            O => \N__3988\,
            I => \N__3980\
        );

    \I__707\ : Span4Mux_s3_v
    port map (
            O => \N__3985\,
            I => \N__3977\
        );

    \I__706\ : IoInMux
    port map (
            O => \N__3984\,
            I => \N__3974\
        );

    \I__705\ : IoInMux
    port map (
            O => \N__3983\,
            I => \N__3971\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__3980\,
            I => \N__3968\
        );

    \I__703\ : Span4Mux_h
    port map (
            O => \N__3977\,
            I => \N__3965\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__3974\,
            I => \N__3962\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__3971\,
            I => \N__3959\
        );

    \I__700\ : IoSpan4Mux
    port map (
            O => \N__3968\,
            I => \N__3956\
        );

    \I__699\ : Span4Mux_h
    port map (
            O => \N__3965\,
            I => \N__3951\
        );

    \I__698\ : Span4Mux_s3_v
    port map (
            O => \N__3962\,
            I => \N__3951\
        );

    \I__697\ : Span4Mux_s2_h
    port map (
            O => \N__3959\,
            I => \N__3948\
        );

    \I__696\ : Span4Mux_s2_h
    port map (
            O => \N__3956\,
            I => \N__3945\
        );

    \I__695\ : Span4Mux_v
    port map (
            O => \N__3951\,
            I => \N__3942\
        );

    \I__694\ : Span4Mux_h
    port map (
            O => \N__3948\,
            I => \N__3939\
        );

    \I__693\ : Sp12to4
    port map (
            O => \N__3945\,
            I => \N__3936\
        );

    \I__692\ : Span4Mux_v
    port map (
            O => \N__3942\,
            I => \N__3933\
        );

    \I__691\ : Span4Mux_h
    port map (
            O => \N__3939\,
            I => \N__3930\
        );

    \I__690\ : Span12Mux_s11_h
    port map (
            O => \N__3936\,
            I => \N__3927\
        );

    \I__689\ : Span4Mux_v
    port map (
            O => \N__3933\,
            I => \N__3924\
        );

    \I__688\ : Span4Mux_h
    port map (
            O => \N__3930\,
            I => \N__3921\
        );

    \I__687\ : Odrv12
    port map (
            O => \N__3927\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__686\ : Odrv4
    port map (
            O => \N__3924\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__685\ : Odrv4
    port map (
            O => \N__3921\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__684\ : InMux
    port map (
            O => \N__3914\,
            I => \N__3911\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__3911\,
            I => \N__3906\
        );

    \I__682\ : InMux
    port map (
            O => \N__3910\,
            I => \N__3901\
        );

    \I__681\ : InMux
    port map (
            O => \N__3909\,
            I => \N__3901\
        );

    \I__680\ : Span4Mux_v
    port map (
            O => \N__3906\,
            I => \N__3896\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__3901\,
            I => \N__3896\
        );

    \I__678\ : Span4Mux_v
    port map (
            O => \N__3896\,
            I => \N__3893\
        );

    \I__677\ : Span4Mux_v
    port map (
            O => \N__3893\,
            I => \N__3890\
        );

    \I__676\ : Sp12to4
    port map (
            O => \N__3890\,
            I => \N__3887\
        );

    \I__675\ : Span12Mux_h
    port map (
            O => \N__3887\,
            I => \N__3884\
        );

    \I__674\ : Odrv12
    port map (
            O => \N__3884\,
            I => \D_UU_AMIGA_in_1\
        );

    \I__673\ : InMux
    port map (
            O => \N__3881\,
            I => \N__3878\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__3878\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\
        );

    \I__671\ : InMux
    port map (
            O => \N__3875\,
            I => \N__3872\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__3872\,
            I => \N__3869\
        );

    \I__669\ : Span4Mux_v
    port map (
            O => \N__3869\,
            I => \N__3866\
        );

    \I__668\ : Sp12to4
    port map (
            O => \N__3866\,
            I => \N__3863\
        );

    \I__667\ : Span12Mux_h
    port map (
            O => \N__3863\,
            I => \N__3860\
        );

    \I__666\ : Odrv12
    port map (
            O => \N__3860\,
            I => \D_UU_040_in_2\
        );

    \I__665\ : IoInMux
    port map (
            O => \N__3857\,
            I => \N__3853\
        );

    \I__664\ : InMux
    port map (
            O => \N__3856\,
            I => \N__3850\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__3853\,
            I => \N__3847\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__3850\,
            I => \N__3844\
        );

    \I__661\ : Span12Mux_s9_h
    port map (
            O => \N__3847\,
            I => \N__3841\
        );

    \I__660\ : Span12Mux_v
    port map (
            O => \N__3844\,
            I => \N__3838\
        );

    \I__659\ : Span12Mux_v
    port map (
            O => \N__3841\,
            I => \N__3835\
        );

    \I__658\ : Span12Mux_v
    port map (
            O => \N__3838\,
            I => \N__3832\
        );

    \I__657\ : Span12Mux_h
    port map (
            O => \N__3835\,
            I => \N__3829\
        );

    \I__656\ : Span12Mux_h
    port map (
            O => \N__3832\,
            I => \N__3826\
        );

    \I__655\ : Odrv12
    port map (
            O => \N__3829\,
            I => \D_LM_040_in_2\
        );

    \I__654\ : Odrv12
    port map (
            O => \N__3826\,
            I => \D_LM_040_in_2\
        );

    \I__653\ : IoInMux
    port map (
            O => \N__3821\,
            I => \N__3818\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__3818\,
            I => \N__3815\
        );

    \I__651\ : IoSpan4Mux
    port map (
            O => \N__3815\,
            I => \N__3812\
        );

    \I__650\ : Sp12to4
    port map (
            O => \N__3812\,
            I => \N__3809\
        );

    \I__649\ : Span12Mux_s6_v
    port map (
            O => \N__3809\,
            I => \N__3806\
        );

    \I__648\ : Odrv12
    port map (
            O => \N__3806\,
            I => \un1_D_UU_040_2\
        );

    \I__647\ : IoInMux
    port map (
            O => \N__3803\,
            I => \N__3799\
        );

    \I__646\ : InMux
    port map (
            O => \N__3802\,
            I => \N__3796\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__3799\,
            I => \N__3793\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__3796\,
            I => \N__3790\
        );

    \I__643\ : IoSpan4Mux
    port map (
            O => \N__3793\,
            I => \N__3787\
        );

    \I__642\ : Span4Mux_h
    port map (
            O => \N__3790\,
            I => \N__3784\
        );

    \I__641\ : Span4Mux_s3_h
    port map (
            O => \N__3787\,
            I => \N__3781\
        );

    \I__640\ : Sp12to4
    port map (
            O => \N__3784\,
            I => \N__3778\
        );

    \I__639\ : Sp12to4
    port map (
            O => \N__3781\,
            I => \N__3775\
        );

    \I__638\ : Span12Mux_v
    port map (
            O => \N__3778\,
            I => \N__3772\
        );

    \I__637\ : Span12Mux_v
    port map (
            O => \N__3775\,
            I => \N__3769\
        );

    \I__636\ : Span12Mux_v
    port map (
            O => \N__3772\,
            I => \N__3764\
        );

    \I__635\ : Span12Mux_h
    port map (
            O => \N__3769\,
            I => \N__3764\
        );

    \I__634\ : Span12Mux_h
    port map (
            O => \N__3764\,
            I => \N__3761\
        );

    \I__633\ : Odrv12
    port map (
            O => \N__3761\,
            I => \D_LL_040_in_5\
        );

    \I__632\ : InMux
    port map (
            O => \N__3758\,
            I => \N__3755\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__3755\,
            I => \N__3752\
        );

    \I__630\ : Span4Mux_v
    port map (
            O => \N__3752\,
            I => \N__3749\
        );

    \I__629\ : Span4Mux_h
    port map (
            O => \N__3749\,
            I => \N__3746\
        );

    \I__628\ : Sp12to4
    port map (
            O => \N__3746\,
            I => \N__3743\
        );

    \I__627\ : Span12Mux_h
    port map (
            O => \N__3743\,
            I => \N__3740\
        );

    \I__626\ : Odrv12
    port map (
            O => \N__3740\,
            I => \D_UM_040_in_5\
        );

    \I__625\ : IoInMux
    port map (
            O => \N__3737\,
            I => \N__3734\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3734\,
            I => \N__3731\
        );

    \I__623\ : Span4Mux_s0_v
    port map (
            O => \N__3731\,
            I => \N__3728\
        );

    \I__622\ : Sp12to4
    port map (
            O => \N__3728\,
            I => \N__3725\
        );

    \I__621\ : Span12Mux_h
    port map (
            O => \N__3725\,
            I => \N__3722\
        );

    \I__620\ : Odrv12
    port map (
            O => \N__3722\,
            I => \un1_D_UM_040_5\
        );

    \I__619\ : IoInMux
    port map (
            O => \N__3719\,
            I => \N__3716\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__3716\,
            I => \N__3713\
        );

    \I__617\ : Odrv12
    port map (
            O => \N__3713\,
            I => \LBENn_c_i_0\
        );

    \I__616\ : InMux
    port map (
            O => \N__3710\,
            I => \N__3707\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__3707\,
            I => \N__3704\
        );

    \I__614\ : Span4Mux_v
    port map (
            O => \N__3704\,
            I => \N__3701\
        );

    \I__613\ : Sp12to4
    port map (
            O => \N__3701\,
            I => \N__3698\
        );

    \I__612\ : Span12Mux_h
    port map (
            O => \N__3698\,
            I => \N__3695\
        );

    \I__611\ : Odrv12
    port map (
            O => \N__3695\,
            I => \D_LL_AMIGA_in_6\
        );

    \I__610\ : IoInMux
    port map (
            O => \N__3692\,
            I => \N__3689\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__3689\,
            I => \N__3686\
        );

    \I__608\ : IoSpan4Mux
    port map (
            O => \N__3686\,
            I => \N__3683\
        );

    \I__607\ : Span4Mux_s3_h
    port map (
            O => \N__3683\,
            I => \N__3680\
        );

    \I__606\ : Sp12to4
    port map (
            O => \N__3680\,
            I => \N__3677\
        );

    \I__605\ : Span12Mux_h
    port map (
            O => \N__3677\,
            I => \N__3674\
        );

    \I__604\ : Odrv12
    port map (
            O => \N__3674\,
            I => \un1_D_LL_AMIGA_6\
        );

    \I__603\ : InMux
    port map (
            O => \N__3671\,
            I => \N__3668\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__3668\,
            I => \N__3665\
        );

    \I__601\ : Span4Mux_v
    port map (
            O => \N__3665\,
            I => \N__3662\
        );

    \I__600\ : Sp12to4
    port map (
            O => \N__3662\,
            I => \N__3659\
        );

    \I__599\ : Span12Mux_h
    port map (
            O => \N__3659\,
            I => \N__3656\
        );

    \I__598\ : Odrv12
    port map (
            O => \N__3656\,
            I => \D_LL_AMIGA_in_5\
        );

    \I__597\ : IoInMux
    port map (
            O => \N__3653\,
            I => \N__3650\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3650\,
            I => \N__3647\
        );

    \I__595\ : IoSpan4Mux
    port map (
            O => \N__3647\,
            I => \N__3644\
        );

    \I__594\ : Span4Mux_s3_h
    port map (
            O => \N__3644\,
            I => \N__3641\
        );

    \I__593\ : Sp12to4
    port map (
            O => \N__3641\,
            I => \N__3638\
        );

    \I__592\ : Span12Mux_h
    port map (
            O => \N__3638\,
            I => \N__3635\
        );

    \I__591\ : Odrv12
    port map (
            O => \N__3635\,
            I => \un1_D_LL_AMIGA_5\
        );

    \I__590\ : InMux
    port map (
            O => \N__3632\,
            I => \N__3629\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3629\,
            I => \N__3626\
        );

    \I__588\ : Sp12to4
    port map (
            O => \N__3626\,
            I => \N__3622\
        );

    \I__587\ : InMux
    port map (
            O => \N__3625\,
            I => \N__3619\
        );

    \I__586\ : Span12Mux_v
    port map (
            O => \N__3622\,
            I => \N__3614\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__3619\,
            I => \N__3614\
        );

    \I__584\ : Span12Mux_h
    port map (
            O => \N__3614\,
            I => \N__3611\
        );

    \I__583\ : Odrv12
    port map (
            O => \N__3611\,
            I => \A_040_c_1\
        );

    \I__582\ : InMux
    port map (
            O => \N__3608\,
            I => \N__3605\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__3605\,
            I => \N__3602\
        );

    \I__580\ : Span4Mux_v
    port map (
            O => \N__3602\,
            I => \N__3599\
        );

    \I__579\ : Sp12to4
    port map (
            O => \N__3599\,
            I => \N__3596\
        );

    \I__578\ : Span12Mux_h
    port map (
            O => \N__3596\,
            I => \N__3593\
        );

    \I__577\ : Odrv12
    port map (
            O => \N__3593\,
            I => \D_LL_AMIGA_in_7\
        );

    \I__576\ : IoInMux
    port map (
            O => \N__3590\,
            I => \N__3587\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__3587\,
            I => \N__3584\
        );

    \I__574\ : IoSpan4Mux
    port map (
            O => \N__3584\,
            I => \N__3581\
        );

    \I__573\ : Span4Mux_s3_h
    port map (
            O => \N__3581\,
            I => \N__3578\
        );

    \I__572\ : Sp12to4
    port map (
            O => \N__3578\,
            I => \N__3575\
        );

    \I__571\ : Span12Mux_h
    port map (
            O => \N__3575\,
            I => \N__3572\
        );

    \I__570\ : Odrv12
    port map (
            O => \N__3572\,
            I => \un1_D_LL_AMIGA_7\
        );

    \I__569\ : InMux
    port map (
            O => \N__3569\,
            I => \N__3566\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__3566\,
            I => \N__3563\
        );

    \I__567\ : Span4Mux_v
    port map (
            O => \N__3563\,
            I => \N__3560\
        );

    \I__566\ : Sp12to4
    port map (
            O => \N__3560\,
            I => \N__3557\
        );

    \I__565\ : Span12Mux_h
    port map (
            O => \N__3557\,
            I => \N__3554\
        );

    \I__564\ : Odrv12
    port map (
            O => \N__3554\,
            I => \D_UU_040_in_4\
        );

    \I__563\ : IoInMux
    port map (
            O => \N__3551\,
            I => \N__3548\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3548\,
            I => \N__3545\
        );

    \I__561\ : Span4Mux_s1_h
    port map (
            O => \N__3545\,
            I => \N__3542\
        );

    \I__560\ : Sp12to4
    port map (
            O => \N__3542\,
            I => \N__3538\
        );

    \I__559\ : InMux
    port map (
            O => \N__3541\,
            I => \N__3535\
        );

    \I__558\ : Span12Mux_v
    port map (
            O => \N__3538\,
            I => \N__3532\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__3535\,
            I => \N__3529\
        );

    \I__556\ : Span12Mux_h
    port map (
            O => \N__3532\,
            I => \N__3526\
        );

    \I__555\ : Span12Mux_h
    port map (
            O => \N__3529\,
            I => \N__3523\
        );

    \I__554\ : Span12Mux_h
    port map (
            O => \N__3526\,
            I => \N__3520\
        );

    \I__553\ : Span12Mux_v
    port map (
            O => \N__3523\,
            I => \N__3517\
        );

    \I__552\ : Odrv12
    port map (
            O => \N__3520\,
            I => \D_LM_040_in_4\
        );

    \I__551\ : Odrv12
    port map (
            O => \N__3517\,
            I => \D_LM_040_in_4\
        );

    \I__550\ : IoInMux
    port map (
            O => \N__3512\,
            I => \N__3509\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3509\,
            I => \N__3506\
        );

    \I__548\ : Span4Mux_s2_v
    port map (
            O => \N__3506\,
            I => \N__3503\
        );

    \I__547\ : Span4Mux_h
    port map (
            O => \N__3503\,
            I => \N__3500\
        );

    \I__546\ : Span4Mux_v
    port map (
            O => \N__3500\,
            I => \N__3497\
        );

    \I__545\ : Odrv4
    port map (
            O => \N__3497\,
            I => \un1_D_UU_040_4\
        );

    \I__544\ : InMux
    port map (
            O => \N__3494\,
            I => \N__3491\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__3491\,
            I => \N__3488\
        );

    \I__542\ : Span4Mux_v
    port map (
            O => \N__3488\,
            I => \N__3485\
        );

    \I__541\ : Span4Mux_h
    port map (
            O => \N__3485\,
            I => \N__3482\
        );

    \I__540\ : Sp12to4
    port map (
            O => \N__3482\,
            I => \N__3479\
        );

    \I__539\ : Span12Mux_h
    port map (
            O => \N__3479\,
            I => \N__3476\
        );

    \I__538\ : Odrv12
    port map (
            O => \N__3476\,
            I => \D_UU_040_in_0\
        );

    \I__537\ : IoInMux
    port map (
            O => \N__3473\,
            I => \N__3470\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__3470\,
            I => \N__3466\
        );

    \I__535\ : InMux
    port map (
            O => \N__3469\,
            I => \N__3463\
        );

    \I__534\ : IoSpan4Mux
    port map (
            O => \N__3466\,
            I => \N__3460\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3463\,
            I => \N__3457\
        );

    \I__532\ : IoSpan4Mux
    port map (
            O => \N__3460\,
            I => \N__3454\
        );

    \I__531\ : Sp12to4
    port map (
            O => \N__3457\,
            I => \N__3451\
        );

    \I__530\ : Span4Mux_s2_h
    port map (
            O => \N__3454\,
            I => \N__3448\
        );

    \I__529\ : Span12Mux_v
    port map (
            O => \N__3451\,
            I => \N__3445\
        );

    \I__528\ : Sp12to4
    port map (
            O => \N__3448\,
            I => \N__3442\
        );

    \I__527\ : Span12Mux_v
    port map (
            O => \N__3445\,
            I => \N__3437\
        );

    \I__526\ : Span12Mux_h
    port map (
            O => \N__3442\,
            I => \N__3437\
        );

    \I__525\ : Span12Mux_h
    port map (
            O => \N__3437\,
            I => \N__3434\
        );

    \I__524\ : Odrv12
    port map (
            O => \N__3434\,
            I => \D_LM_040_in_0\
        );

    \I__523\ : IoInMux
    port map (
            O => \N__3431\,
            I => \N__3428\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__3428\,
            I => \N__3425\
        );

    \I__521\ : IoSpan4Mux
    port map (
            O => \N__3425\,
            I => \N__3422\
        );

    \I__520\ : Span4Mux_s2_v
    port map (
            O => \N__3422\,
            I => \N__3419\
        );

    \I__519\ : Span4Mux_v
    port map (
            O => \N__3419\,
            I => \N__3416\
        );

    \I__518\ : Odrv4
    port map (
            O => \N__3416\,
            I => \un1_D_UU_040_0\
        );

    \I__517\ : IoInMux
    port map (
            O => \N__3413\,
            I => \N__3410\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__3410\,
            I => \N__3407\
        );

    \I__515\ : IoSpan4Mux
    port map (
            O => \N__3407\,
            I => \N__3404\
        );

    \I__514\ : Sp12to4
    port map (
            O => \N__3404\,
            I => \N__3401\
        );

    \I__513\ : Span12Mux_s7_h
    port map (
            O => \N__3401\,
            I => \N__3398\
        );

    \I__512\ : Odrv12
    port map (
            O => \N__3398\,
            I => \un1_D_UM_AMIGA_0\
        );

    \I__511\ : InMux
    port map (
            O => \N__3395\,
            I => \N__3392\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__3392\,
            I => \N__3389\
        );

    \I__509\ : Span12Mux_h
    port map (
            O => \N__3389\,
            I => \N__3386\
        );

    \I__508\ : Odrv12
    port map (
            O => \N__3386\,
            I => \D_LM_AMIGA_in_1\
        );

    \I__507\ : IoInMux
    port map (
            O => \N__3383\,
            I => \N__3380\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__3380\,
            I => \N__3377\
        );

    \I__505\ : Span4Mux_s0_h
    port map (
            O => \N__3377\,
            I => \N__3374\
        );

    \I__504\ : Span4Mux_h
    port map (
            O => \N__3374\,
            I => \N__3371\
        );

    \I__503\ : Span4Mux_h
    port map (
            O => \N__3371\,
            I => \N__3368\
        );

    \I__502\ : Sp12to4
    port map (
            O => \N__3368\,
            I => \N__3365\
        );

    \I__501\ : Span12Mux_v
    port map (
            O => \N__3365\,
            I => \N__3362\
        );

    \I__500\ : Odrv12
    port map (
            O => \N__3362\,
            I => \un1_D_LM_AMIGA_1\
        );

    \I__499\ : InMux
    port map (
            O => \N__3359\,
            I => \N__3356\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3356\,
            I => \N__3353\
        );

    \I__497\ : Span4Mux_v
    port map (
            O => \N__3353\,
            I => \N__3349\
        );

    \I__496\ : InMux
    port map (
            O => \N__3352\,
            I => \N__3346\
        );

    \I__495\ : Span4Mux_v
    port map (
            O => \N__3349\,
            I => \N__3343\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__3346\,
            I => \N__3340\
        );

    \I__493\ : Span4Mux_v
    port map (
            O => \N__3343\,
            I => \N__3336\
        );

    \I__492\ : Span4Mux_v
    port map (
            O => \N__3340\,
            I => \N__3333\
        );

    \I__491\ : InMux
    port map (
            O => \N__3339\,
            I => \N__3330\
        );

    \I__490\ : Sp12to4
    port map (
            O => \N__3336\,
            I => \N__3323\
        );

    \I__489\ : Sp12to4
    port map (
            O => \N__3333\,
            I => \N__3323\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__3330\,
            I => \N__3323\
        );

    \I__487\ : Span12Mux_h
    port map (
            O => \N__3323\,
            I => \N__3320\
        );

    \I__486\ : Odrv12
    port map (
            O => \N__3320\,
            I => \D_UM_AMIGA_in_0\
        );

    \I__485\ : InMux
    port map (
            O => \N__3317\,
            I => \N__3314\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__3314\,
            I => \N__3311\
        );

    \I__483\ : Odrv4
    port map (
            O => \N__3311\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\
        );

    \I__482\ : IoInMux
    port map (
            O => \N__3308\,
            I => \N__3305\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__3305\,
            I => \N__3302\
        );

    \I__480\ : Span4Mux_s2_h
    port map (
            O => \N__3302\,
            I => \N__3299\
        );

    \I__479\ : Span4Mux_h
    port map (
            O => \N__3299\,
            I => \N__3296\
        );

    \I__478\ : Sp12to4
    port map (
            O => \N__3296\,
            I => \N__3293\
        );

    \I__477\ : Span12Mux_v
    port map (
            O => \N__3293\,
            I => \N__3290\
        );

    \I__476\ : Span12Mux_h
    port map (
            O => \N__3290\,
            I => \N__3287\
        );

    \I__475\ : Odrv12
    port map (
            O => \N__3287\,
            I => \un1_D_UM_AMIGA_1\
        );

    \I__474\ : InMux
    port map (
            O => \N__3284\,
            I => \N__3281\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__3281\,
            I => \N__3278\
        );

    \I__472\ : Span4Mux_v
    port map (
            O => \N__3278\,
            I => \N__3273\
        );

    \I__471\ : InMux
    port map (
            O => \N__3277\,
            I => \N__3268\
        );

    \I__470\ : InMux
    port map (
            O => \N__3276\,
            I => \N__3268\
        );

    \I__469\ : Sp12to4
    port map (
            O => \N__3273\,
            I => \N__3265\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__3268\,
            I => \N__3262\
        );

    \I__467\ : Span12Mux_h
    port map (
            O => \N__3265\,
            I => \N__3259\
        );

    \I__466\ : Span12Mux_v
    port map (
            O => \N__3262\,
            I => \N__3256\
        );

    \I__465\ : Span12Mux_v
    port map (
            O => \N__3259\,
            I => \N__3253\
        );

    \I__464\ : Span12Mux_h
    port map (
            O => \N__3256\,
            I => \N__3250\
        );

    \I__463\ : Odrv12
    port map (
            O => \N__3253\,
            I => \D_UM_AMIGA_in_1\
        );

    \I__462\ : Odrv12
    port map (
            O => \N__3250\,
            I => \D_UM_AMIGA_in_1\
        );

    \I__461\ : InMux
    port map (
            O => \N__3245\,
            I => \N__3242\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__3242\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\
        );

    \I__459\ : IoInMux
    port map (
            O => \N__3239\,
            I => \N__3236\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__3236\,
            I => \N__3233\
        );

    \I__457\ : IoSpan4Mux
    port map (
            O => \N__3233\,
            I => \N__3230\
        );

    \I__456\ : Span4Mux_s3_h
    port map (
            O => \N__3230\,
            I => \N__3227\
        );

    \I__455\ : Sp12to4
    port map (
            O => \N__3227\,
            I => \N__3224\
        );

    \I__454\ : Span12Mux_s8_h
    port map (
            O => \N__3224\,
            I => \N__3221\
        );

    \I__453\ : Span12Mux_v
    port map (
            O => \N__3221\,
            I => \N__3218\
        );

    \I__452\ : Odrv12
    port map (
            O => \N__3218\,
            I => \un1_D_UU_AMIGA_1\
        );

    \I__451\ : InMux
    port map (
            O => \N__3215\,
            I => \N__3212\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__3212\,
            I => \N__3209\
        );

    \I__449\ : Span12Mux_v
    port map (
            O => \N__3209\,
            I => \N__3206\
        );

    \I__448\ : Odrv12
    port map (
            O => \N__3206\,
            I => \D_LM_AMIGA_in_5\
        );

    \I__447\ : IoInMux
    port map (
            O => \N__3203\,
            I => \N__3200\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__3200\,
            I => \N__3197\
        );

    \I__445\ : IoSpan4Mux
    port map (
            O => \N__3197\,
            I => \N__3194\
        );

    \I__444\ : Span4Mux_s3_h
    port map (
            O => \N__3194\,
            I => \N__3191\
        );

    \I__443\ : Sp12to4
    port map (
            O => \N__3191\,
            I => \N__3188\
        );

    \I__442\ : Span12Mux_s8_h
    port map (
            O => \N__3188\,
            I => \N__3185\
        );

    \I__441\ : Span12Mux_h
    port map (
            O => \N__3185\,
            I => \N__3182\
        );

    \I__440\ : Odrv12
    port map (
            O => \N__3182\,
            I => \un1_D_LM_AMIGA_5\
        );

    \I__439\ : InMux
    port map (
            O => \N__3179\,
            I => \N__3176\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__3176\,
            I => \N__3173\
        );

    \I__437\ : Span12Mux_v
    port map (
            O => \N__3173\,
            I => \N__3170\
        );

    \I__436\ : Odrv12
    port map (
            O => \N__3170\,
            I => \D_LM_AMIGA_in_7\
        );

    \I__435\ : IoInMux
    port map (
            O => \N__3167\,
            I => \N__3164\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__3164\,
            I => \N__3161\
        );

    \I__433\ : Span12Mux_s8_h
    port map (
            O => \N__3161\,
            I => \N__3158\
        );

    \I__432\ : Span12Mux_h
    port map (
            O => \N__3158\,
            I => \N__3155\
        );

    \I__431\ : Odrv12
    port map (
            O => \N__3155\,
            I => \un1_D_LM_AMIGA_7\
        );

    \I__430\ : InMux
    port map (
            O => \N__3152\,
            I => \N__3149\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__3149\,
            I => \N__3146\
        );

    \I__428\ : Span4Mux_h
    port map (
            O => \N__3146\,
            I => \N__3143\
        );

    \I__427\ : Span4Mux_v
    port map (
            O => \N__3143\,
            I => \N__3140\
        );

    \I__426\ : Sp12to4
    port map (
            O => \N__3140\,
            I => \N__3137\
        );

    \I__425\ : Odrv12
    port map (
            O => \N__3137\,
            I => \D_LM_AMIGA_in_6\
        );

    \I__424\ : IoInMux
    port map (
            O => \N__3134\,
            I => \N__3131\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__3131\,
            I => \N__3128\
        );

    \I__422\ : Span12Mux_s9_h
    port map (
            O => \N__3128\,
            I => \N__3125\
        );

    \I__421\ : Odrv12
    port map (
            O => \N__3125\,
            I => \un1_D_LM_AMIGA_6\
        );

    \I__420\ : IoInMux
    port map (
            O => \N__3122\,
            I => \N__3118\
        );

    \I__419\ : IoInMux
    port map (
            O => \N__3121\,
            I => \N__3115\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__3118\,
            I => \N__3112\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__3115\,
            I => \N__3109\
        );

    \I__416\ : Span4Mux_s2_v
    port map (
            O => \N__3112\,
            I => \N__3106\
        );

    \I__415\ : Span4Mux_s2_v
    port map (
            O => \N__3109\,
            I => \N__3103\
        );

    \I__414\ : Span4Mux_h
    port map (
            O => \N__3106\,
            I => \N__3100\
        );

    \I__413\ : Span4Mux_h
    port map (
            O => \N__3103\,
            I => \N__3097\
        );

    \I__412\ : Span4Mux_v
    port map (
            O => \N__3100\,
            I => \N__3092\
        );

    \I__411\ : Span4Mux_v
    port map (
            O => \N__3097\,
            I => \N__3092\
        );

    \I__410\ : Odrv4
    port map (
            O => \N__3092\,
            I => \CONSTANT_ONE_NET\
        );

    \I__409\ : IoInMux
    port map (
            O => \N__3089\,
            I => \N__3086\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__3086\,
            I => \N__3083\
        );

    \I__407\ : IoSpan4Mux
    port map (
            O => \N__3083\,
            I => \N__3079\
        );

    \I__406\ : InMux
    port map (
            O => \N__3082\,
            I => \N__3076\
        );

    \I__405\ : Span4Mux_s2_h
    port map (
            O => \N__3079\,
            I => \N__3073\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__3076\,
            I => \N__3070\
        );

    \I__403\ : Sp12to4
    port map (
            O => \N__3073\,
            I => \N__3067\
        );

    \I__402\ : Span4Mux_v
    port map (
            O => \N__3070\,
            I => \N__3064\
        );

    \I__401\ : Span12Mux_h
    port map (
            O => \N__3067\,
            I => \N__3059\
        );

    \I__400\ : Sp12to4
    port map (
            O => \N__3064\,
            I => \N__3059\
        );

    \I__399\ : Span12Mux_h
    port map (
            O => \N__3059\,
            I => \N__3056\
        );

    \I__398\ : Odrv12
    port map (
            O => \N__3056\,
            I => \D_LM_040_in_7\
        );

    \I__397\ : InMux
    port map (
            O => \N__3053\,
            I => \N__3050\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__3050\,
            I => \N__3047\
        );

    \I__395\ : Span4Mux_v
    port map (
            O => \N__3047\,
            I => \N__3044\
        );

    \I__394\ : Span4Mux_h
    port map (
            O => \N__3044\,
            I => \N__3041\
        );

    \I__393\ : Sp12to4
    port map (
            O => \N__3041\,
            I => \N__3038\
        );

    \I__392\ : Span12Mux_h
    port map (
            O => \N__3038\,
            I => \N__3035\
        );

    \I__391\ : Odrv12
    port map (
            O => \N__3035\,
            I => \D_UU_040_in_7\
        );

    \I__390\ : IoInMux
    port map (
            O => \N__3032\,
            I => \N__3029\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__3029\,
            I => \N__3026\
        );

    \I__388\ : Span4Mux_s3_v
    port map (
            O => \N__3026\,
            I => \N__3023\
        );

    \I__387\ : Sp12to4
    port map (
            O => \N__3023\,
            I => \N__3020\
        );

    \I__386\ : Span12Mux_s11_h
    port map (
            O => \N__3020\,
            I => \N__3017\
        );

    \I__385\ : Odrv12
    port map (
            O => \N__3017\,
            I => \un1_D_UU_040_7\
        );

    \I__384\ : InMux
    port map (
            O => \N__3014\,
            I => \N__3011\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__3011\,
            I => \N__3008\
        );

    \I__382\ : Span12Mux_h
    port map (
            O => \N__3008\,
            I => \N__3005\
        );

    \I__381\ : Odrv12
    port map (
            O => \N__3005\,
            I => \D_LM_AMIGA_in_3\
        );

    \I__380\ : IoInMux
    port map (
            O => \N__3002\,
            I => \N__2999\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__2999\,
            I => \N__2996\
        );

    \I__378\ : Span4Mux_s0_h
    port map (
            O => \N__2996\,
            I => \N__2993\
        );

    \I__377\ : Sp12to4
    port map (
            O => \N__2993\,
            I => \N__2990\
        );

    \I__376\ : Span12Mux_v
    port map (
            O => \N__2990\,
            I => \N__2987\
        );

    \I__375\ : Span12Mux_h
    port map (
            O => \N__2987\,
            I => \N__2984\
        );

    \I__374\ : Odrv12
    port map (
            O => \N__2984\,
            I => \un1_D_LM_AMIGA_3\
        );

    \I__373\ : InMux
    port map (
            O => \N__2981\,
            I => \N__2978\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__2978\,
            I => \N__2975\
        );

    \I__371\ : Span4Mux_v
    port map (
            O => \N__2975\,
            I => \N__2972\
        );

    \I__370\ : Sp12to4
    port map (
            O => \N__2972\,
            I => \N__2969\
        );

    \I__369\ : Span12Mux_h
    port map (
            O => \N__2969\,
            I => \N__2966\
        );

    \I__368\ : Odrv12
    port map (
            O => \N__2966\,
            I => \D_UM_040_in_0\
        );

    \I__367\ : IoInMux
    port map (
            O => \N__2963\,
            I => \N__2959\
        );

    \I__366\ : InMux
    port map (
            O => \N__2962\,
            I => \N__2956\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__2959\,
            I => \N__2953\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__2956\,
            I => \N__2950\
        );

    \I__363\ : IoSpan4Mux
    port map (
            O => \N__2953\,
            I => \N__2947\
        );

    \I__362\ : Span4Mux_v
    port map (
            O => \N__2950\,
            I => \N__2944\
        );

    \I__361\ : Span4Mux_s2_h
    port map (
            O => \N__2947\,
            I => \N__2941\
        );

    \I__360\ : Sp12to4
    port map (
            O => \N__2944\,
            I => \N__2938\
        );

    \I__359\ : Sp12to4
    port map (
            O => \N__2941\,
            I => \N__2935\
        );

    \I__358\ : Span12Mux_v
    port map (
            O => \N__2938\,
            I => \N__2930\
        );

    \I__357\ : Span12Mux_h
    port map (
            O => \N__2935\,
            I => \N__2930\
        );

    \I__356\ : Span12Mux_h
    port map (
            O => \N__2930\,
            I => \N__2927\
        );

    \I__355\ : Odrv12
    port map (
            O => \N__2927\,
            I => \D_LL_040_in_0\
        );

    \I__354\ : IoInMux
    port map (
            O => \N__2924\,
            I => \N__2921\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__2921\,
            I => \N__2918\
        );

    \I__352\ : Span4Mux_s3_h
    port map (
            O => \N__2918\,
            I => \N__2915\
        );

    \I__351\ : Sp12to4
    port map (
            O => \N__2915\,
            I => \N__2912\
        );

    \I__350\ : Span12Mux_v
    port map (
            O => \N__2912\,
            I => \N__2909\
        );

    \I__349\ : Odrv12
    port map (
            O => \N__2909\,
            I => \un1_D_UM_040_0\
        );

    \I__348\ : InMux
    port map (
            O => \N__2906\,
            I => \N__2903\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__2903\,
            I => \N__2900\
        );

    \I__346\ : Span4Mux_v
    port map (
            O => \N__2900\,
            I => \N__2897\
        );

    \I__345\ : Span4Mux_v
    port map (
            O => \N__2897\,
            I => \N__2894\
        );

    \I__344\ : Sp12to4
    port map (
            O => \N__2894\,
            I => \N__2891\
        );

    \I__343\ : Span12Mux_h
    port map (
            O => \N__2891\,
            I => \N__2888\
        );

    \I__342\ : Odrv12
    port map (
            O => \N__2888\,
            I => \D_UU_040_in_1\
        );

    \I__341\ : IoInMux
    port map (
            O => \N__2885\,
            I => \N__2882\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__2882\,
            I => \N__2878\
        );

    \I__339\ : InMux
    port map (
            O => \N__2881\,
            I => \N__2875\
        );

    \I__338\ : Span4Mux_s3_h
    port map (
            O => \N__2878\,
            I => \N__2872\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__2875\,
            I => \N__2869\
        );

    \I__336\ : Span4Mux_h
    port map (
            O => \N__2872\,
            I => \N__2866\
        );

    \I__335\ : Span4Mux_h
    port map (
            O => \N__2869\,
            I => \N__2863\
        );

    \I__334\ : Span4Mux_h
    port map (
            O => \N__2866\,
            I => \N__2860\
        );

    \I__333\ : Sp12to4
    port map (
            O => \N__2863\,
            I => \N__2857\
        );

    \I__332\ : Sp12to4
    port map (
            O => \N__2860\,
            I => \N__2852\
        );

    \I__331\ : Span12Mux_v
    port map (
            O => \N__2857\,
            I => \N__2852\
        );

    \I__330\ : Span12Mux_v
    port map (
            O => \N__2852\,
            I => \N__2849\
        );

    \I__329\ : Span12Mux_h
    port map (
            O => \N__2849\,
            I => \N__2846\
        );

    \I__328\ : Odrv12
    port map (
            O => \N__2846\,
            I => \D_LM_040_in_1\
        );

    \I__327\ : IoInMux
    port map (
            O => \N__2843\,
            I => \N__2840\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__2840\,
            I => \N__2837\
        );

    \I__325\ : Span4Mux_s3_h
    port map (
            O => \N__2837\,
            I => \N__2834\
        );

    \I__324\ : Sp12to4
    port map (
            O => \N__2834\,
            I => \N__2831\
        );

    \I__323\ : Span12Mux_s8_v
    port map (
            O => \N__2831\,
            I => \N__2828\
        );

    \I__322\ : Odrv12
    port map (
            O => \N__2828\,
            I => \un1_D_UU_040_1\
        );

    \I__321\ : InMux
    port map (
            O => \N__2825\,
            I => \N__2822\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__2822\,
            I => \N__2819\
        );

    \I__319\ : Span4Mux_h
    port map (
            O => \N__2819\,
            I => \N__2816\
        );

    \I__318\ : Span4Mux_v
    port map (
            O => \N__2816\,
            I => \N__2813\
        );

    \I__317\ : Odrv4
    port map (
            O => \N__2813\,
            I => \A_040_c_0\
        );

    \I__316\ : IoInMux
    port map (
            O => \N__2810\,
            I => \N__2807\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__2807\,
            I => \N__2804\
        );

    \I__314\ : Span4Mux_s2_v
    port map (
            O => \N__2804\,
            I => \N__2801\
        );

    \I__313\ : Span4Mux_v
    port map (
            O => \N__2801\,
            I => \N__2798\
        );

    \I__312\ : Odrv4
    port map (
            O => \N__2798\,
            I => \A_AMIGA_c_0\
        );

    \I__311\ : IoInMux
    port map (
            O => \N__2795\,
            I => \N__2792\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__2792\,
            I => \N__2789\
        );

    \I__309\ : Span4Mux_s3_v
    port map (
            O => \N__2789\,
            I => \N__2786\
        );

    \I__308\ : Odrv4
    port map (
            O => \N__2786\,
            I => \U111_CYCLE_SM_A_AMIGA_0_i_1\
        );

    \I__307\ : InMux
    port map (
            O => \N__2783\,
            I => \N__2780\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__2780\,
            I => \N__2777\
        );

    \I__305\ : Span4Mux_v
    port map (
            O => \N__2777\,
            I => \N__2774\
        );

    \I__304\ : Span4Mux_h
    port map (
            O => \N__2774\,
            I => \N__2771\
        );

    \I__303\ : Span4Mux_h
    port map (
            O => \N__2771\,
            I => \N__2768\
        );

    \I__302\ : Span4Mux_v
    port map (
            O => \N__2768\,
            I => \N__2765\
        );

    \I__301\ : Odrv4
    port map (
            O => \N__2765\,
            I => \D_LL_AMIGA_in_0\
        );

    \I__300\ : IoInMux
    port map (
            O => \N__2762\,
            I => \N__2759\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__2759\,
            I => \N__2756\
        );

    \I__298\ : Span4Mux_s0_h
    port map (
            O => \N__2756\,
            I => \N__2753\
        );

    \I__297\ : Sp12to4
    port map (
            O => \N__2753\,
            I => \N__2750\
        );

    \I__296\ : Span12Mux_s8_v
    port map (
            O => \N__2750\,
            I => \N__2747\
        );

    \I__295\ : Span12Mux_h
    port map (
            O => \N__2747\,
            I => \N__2744\
        );

    \I__294\ : Odrv12
    port map (
            O => \N__2744\,
            I => \un1_D_LL_AMIGA_0\
        );

    \I__293\ : InMux
    port map (
            O => \N__2741\,
            I => \N__2738\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__2738\,
            I => \N__2735\
        );

    \I__291\ : Span4Mux_v
    port map (
            O => \N__2735\,
            I => \N__2732\
        );

    \I__290\ : Sp12to4
    port map (
            O => \N__2732\,
            I => \N__2729\
        );

    \I__289\ : Span12Mux_h
    port map (
            O => \N__2729\,
            I => \N__2726\
        );

    \I__288\ : Odrv12
    port map (
            O => \N__2726\,
            I => \D_LL_AMIGA_in_1\
        );

    \I__287\ : IoInMux
    port map (
            O => \N__2723\,
            I => \N__2720\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__2720\,
            I => \N__2717\
        );

    \I__285\ : Span4Mux_s3_h
    port map (
            O => \N__2717\,
            I => \N__2714\
        );

    \I__284\ : Sp12to4
    port map (
            O => \N__2714\,
            I => \N__2711\
        );

    \I__283\ : Span12Mux_s8_v
    port map (
            O => \N__2711\,
            I => \N__2708\
        );

    \I__282\ : Span12Mux_h
    port map (
            O => \N__2708\,
            I => \N__2705\
        );

    \I__281\ : Odrv12
    port map (
            O => \N__2705\,
            I => \un1_D_LL_AMIGA_1\
        );

    \I__280\ : InMux
    port map (
            O => \N__2702\,
            I => \N__2699\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__2699\,
            I => \N__2696\
        );

    \I__278\ : Span12Mux_v
    port map (
            O => \N__2696\,
            I => \N__2693\
        );

    \I__277\ : Odrv12
    port map (
            O => \N__2693\,
            I => \D_LL_AMIGA_in_3\
        );

    \I__276\ : IoInMux
    port map (
            O => \N__2690\,
            I => \N__2687\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2687\,
            I => \N__2684\
        );

    \I__274\ : Span12Mux_s8_h
    port map (
            O => \N__2684\,
            I => \N__2681\
        );

    \I__273\ : Span12Mux_h
    port map (
            O => \N__2681\,
            I => \N__2678\
        );

    \I__272\ : Odrv12
    port map (
            O => \N__2678\,
            I => \un1_D_LL_AMIGA_3\
        );

    \I__271\ : InMux
    port map (
            O => \N__2675\,
            I => \N__2672\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2672\,
            I => \N__2669\
        );

    \I__269\ : Span4Mux_v
    port map (
            O => \N__2669\,
            I => \N__2666\
        );

    \I__268\ : Sp12to4
    port map (
            O => \N__2666\,
            I => \N__2663\
        );

    \I__267\ : Span12Mux_h
    port map (
            O => \N__2663\,
            I => \N__2660\
        );

    \I__266\ : Odrv12
    port map (
            O => \N__2660\,
            I => \D_UM_040_in_6\
        );

    \I__265\ : IoInMux
    port map (
            O => \N__2657\,
            I => \N__2654\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__2654\,
            I => \N__2651\
        );

    \I__263\ : IoSpan4Mux
    port map (
            O => \N__2651\,
            I => \N__2647\
        );

    \I__262\ : InMux
    port map (
            O => \N__2650\,
            I => \N__2644\
        );

    \I__261\ : IoSpan4Mux
    port map (
            O => \N__2647\,
            I => \N__2641\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__2644\,
            I => \N__2638\
        );

    \I__259\ : Span4Mux_s2_h
    port map (
            O => \N__2641\,
            I => \N__2635\
        );

    \I__258\ : Span4Mux_v
    port map (
            O => \N__2638\,
            I => \N__2632\
        );

    \I__257\ : Sp12to4
    port map (
            O => \N__2635\,
            I => \N__2629\
        );

    \I__256\ : Sp12to4
    port map (
            O => \N__2632\,
            I => \N__2626\
        );

    \I__255\ : Span12Mux_h
    port map (
            O => \N__2629\,
            I => \N__2623\
        );

    \I__254\ : Span12Mux_h
    port map (
            O => \N__2626\,
            I => \N__2620\
        );

    \I__253\ : Span12Mux_h
    port map (
            O => \N__2623\,
            I => \N__2615\
        );

    \I__252\ : Span12Mux_v
    port map (
            O => \N__2620\,
            I => \N__2615\
        );

    \I__251\ : Odrv12
    port map (
            O => \N__2615\,
            I => \D_LL_040_in_6\
        );

    \I__250\ : IoInMux
    port map (
            O => \N__2612\,
            I => \N__2609\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__2609\,
            I => \N__2606\
        );

    \I__248\ : Span12Mux_s8_h
    port map (
            O => \N__2606\,
            I => \N__2603\
        );

    \I__247\ : Span12Mux_v
    port map (
            O => \N__2603\,
            I => \N__2600\
        );

    \I__246\ : Odrv12
    port map (
            O => \N__2600\,
            I => \un1_D_UM_040_6\
        );

    \I__245\ : IoInMux
    port map (
            O => \N__2597\,
            I => \N__2594\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__2594\,
            I => \N__2591\
        );

    \I__243\ : Span4Mux_s3_v
    port map (
            O => \N__2591\,
            I => \N__2588\
        );

    \I__242\ : Span4Mux_h
    port map (
            O => \N__2588\,
            I => \N__2585\
        );

    \I__241\ : Sp12to4
    port map (
            O => \N__2585\,
            I => \N__2582\
        );

    \I__240\ : Odrv12
    port map (
            O => \N__2582\,
            I => \LBENn_c_i\
        );

    \I__239\ : InMux
    port map (
            O => \N__2579\,
            I => \N__2576\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__2576\,
            I => \N__2573\
        );

    \I__237\ : Span12Mux_v
    port map (
            O => \N__2573\,
            I => \N__2570\
        );

    \I__236\ : Odrv12
    port map (
            O => \N__2570\,
            I => \D_LM_AMIGA_in_4\
        );

    \I__235\ : IoInMux
    port map (
            O => \N__2567\,
            I => \N__2564\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__2564\,
            I => \N__2561\
        );

    \I__233\ : IoSpan4Mux
    port map (
            O => \N__2561\,
            I => \N__2558\
        );

    \I__232\ : IoSpan4Mux
    port map (
            O => \N__2558\,
            I => \N__2555\
        );

    \I__231\ : Sp12to4
    port map (
            O => \N__2555\,
            I => \N__2552\
        );

    \I__230\ : Span12Mux_s9_h
    port map (
            O => \N__2552\,
            I => \N__2549\
        );

    \I__229\ : Odrv12
    port map (
            O => \N__2549\,
            I => \un1_D_LM_AMIGA_4\
        );

    \I__228\ : IoInMux
    port map (
            O => \N__2546\,
            I => \N__2543\
        );

    \I__227\ : LocalMux
    port map (
            O => \N__2543\,
            I => \N__2540\
        );

    \I__226\ : Span4Mux_s0_v
    port map (
            O => \N__2540\,
            I => \N__2537\
        );

    \I__225\ : Sp12to4
    port map (
            O => \N__2537\,
            I => \N__2534\
        );

    \I__224\ : Span12Mux_h
    port map (
            O => \N__2534\,
            I => \N__2531\
        );

    \I__223\ : Span12Mux_v
    port map (
            O => \N__2531\,
            I => \N__2528\
        );

    \I__222\ : Span12Mux_v
    port map (
            O => \N__2528\,
            I => \N__2525\
        );

    \I__221\ : Odrv12
    port map (
            O => \N__2525\,
            I => \TAn_in\
        );

    \I__220\ : IoInMux
    port map (
            O => \N__2522\,
            I => \N__2519\
        );

    \I__219\ : LocalMux
    port map (
            O => \N__2519\,
            I => \N__2516\
        );

    \I__218\ : Span4Mux_s0_h
    port map (
            O => \N__2516\,
            I => \N__2513\
        );

    \I__217\ : Span4Mux_h
    port map (
            O => \N__2513\,
            I => \N__2510\
        );

    \I__216\ : Span4Mux_h
    port map (
            O => \N__2510\,
            I => \N__2507\
        );

    \I__215\ : Sp12to4
    port map (
            O => \N__2507\,
            I => \N__2504\
        );

    \I__214\ : Span12Mux_v
    port map (
            O => \N__2504\,
            I => \N__2501\
        );

    \I__213\ : Span12Mux_v
    port map (
            O => \N__2501\,
            I => \N__2498\
        );

    \I__212\ : Span12Mux_h
    port map (
            O => \N__2498\,
            I => \N__2495\
        );

    \I__211\ : Odrv12
    port map (
            O => \N__2495\,
            I => \TCIn_c\
        );

    \INVU111_CYCLE_SM.TSnC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.TSnC_net\,
            I => \N__7753\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__5050\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2825\,
            lcout => \A_AMIGA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3625\,
            in2 => \_gnd_net_\,
            in3 => \N__5051\,
            lcout => \U111_CYCLE_SM_A_AMIGA_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6919\,
            in1 => \N__3359\,
            in2 => \_gnd_net_\,
            in3 => \N__2783\,
            lcout => \un1_D_LL_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__2741\,
            in1 => \N__3284\,
            in2 => \_gnd_net_\,
            in3 => \N__6917\,
            lcout => \un1_D_LL_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6918\,
            in1 => \N__6053\,
            in2 => \_gnd_net_\,
            in3 => \N__2702\,
            lcout => \un1_D_LL_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6898\,
            in1 => \N__2675\,
            in2 => \_gnd_net_\,
            in3 => \N__2650\,
            lcout => \un1_D_UM_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \BUFENn_obuf_RNO_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5447\,
            lcout => \LBENn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6899\,
            in1 => \N__6563\,
            in2 => \_gnd_net_\,
            in3 => \N__2579\,
            lcout => \un1_D_LM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6935\,
            in1 => \N__6727\,
            in2 => \_gnd_net_\,
            in3 => \N__3215\,
            lcout => \un1_D_LM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6937\,
            in1 => \N__5181\,
            in2 => \_gnd_net_\,
            in3 => \N__3179\,
            lcout => \un1_D_LM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3152\,
            in1 => \N__4998\,
            in2 => \_gnd_net_\,
            in3 => \N__6936\,
            lcout => \un1_D_LM_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__3082\,
            in1 => \N__3053\,
            in2 => \_gnd_net_\,
            in3 => \N__6920\,
            lcout => \un1_D_UU_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6881\,
            in1 => \N__6119\,
            in2 => \_gnd_net_\,
            in3 => \N__3014\,
            lcout => \un1_D_LM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6880\,
            in1 => \N__2981\,
            in2 => \_gnd_net_\,
            in3 => \N__2962\,
            lcout => \un1_D_UM_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6944\,
            in1 => \N__2906\,
            in2 => \_gnd_net_\,
            in3 => \N__2881\,
            lcout => \un1_D_UU_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6948\,
            in1 => \N__3569\,
            in2 => \_gnd_net_\,
            in3 => \N__3541\,
            lcout => \un1_D_UU_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6947\,
            in1 => \N__3494\,
            in2 => \_gnd_net_\,
            in3 => \N__3469\,
            lcout => \un1_D_UU_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7136\,
            in1 => \N__3317\,
            in2 => \_gnd_net_\,
            in3 => \N__3352\,
            lcout => \un1_D_UM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3395\,
            in1 => \N__3914\,
            in2 => \_gnd_net_\,
            in3 => \N__6790\,
            lcout => \un1_D_LM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_DIS_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__5315\,
            in1 => \N__6481\,
            in2 => \N__5389\,
            in3 => \N__4775\,
            lcout => \U111_CYCLE_SM.TA_DISZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7751\,
            ce => 'H',
            sr => \N__7695\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__3339\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7748\,
            ce => \N__6306\,
            sr => \N__6246\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__3277\,
            in1 => \N__7187\,
            in2 => \_gnd_net_\,
            in3 => \N__3245\,
            lcout => \un1_D_UM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3276\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7742\,
            ce => \N__6288\,
            sr => \N__6243\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNIUR6Q_1_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7188\,
            in1 => \N__3881\,
            in2 => \_gnd_net_\,
            in3 => \N__3910\,
            lcout => \un1_D_UU_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_1_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__3909\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7740\,
            ce => \N__6307\,
            sr => \N__6247\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6946\,
            in1 => \N__3875\,
            in2 => \_gnd_net_\,
            in3 => \N__3856\,
            lcout => \un1_D_UU_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__3802\,
            in1 => \N__3758\,
            in2 => \_gnd_net_\,
            in3 => \N__6945\,
            lcout => \un1_D_UM_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LBENn_c_sbtinv_LC_11_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5428\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \LBENn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3710\,
            in1 => \N__7268\,
            in2 => \_gnd_net_\,
            in3 => \N__6834\,
            lcout => \un1_D_LL_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3671\,
            in1 => \N__4844\,
            in2 => \_gnd_net_\,
            in3 => \N__6833\,
            lcout => \un1_D_LL_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6435\,
            in2 => \_gnd_net_\,
            in3 => \N__3632\,
            lcout => \U111_CYCLE_SM.FLIP_WORD_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3608\,
            in1 => \N__5902\,
            in2 => \_gnd_net_\,
            in3 => \N__6832\,
            lcout => \un1_D_LL_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4436\,
            in1 => \N__4943\,
            in2 => \_gnd_net_\,
            in3 => \N__6831\,
            lcout => \un1_D_LM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5637\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TSn_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5638\,
            in2 => \_gnd_net_\,
            in3 => \N__4096\,
            lcout => \TSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TSnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_RNIDDAN_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7775\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5446\,
            lcout => \D_UU_AMIGA_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LATCH_EN_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__4759\,
            in1 => \N__7809\,
            in2 => \N__7158\,
            in3 => \N__4463\,
            lcout => \U111_CYCLE_SM.LATCH_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7752\,
            ce => 'H',
            sr => \N__7691\
        );

    \U111_CYCLE_SM.TS_EN_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011111111"
        )
    port map (
            in0 => \N__4766\,
            in1 => \N__5015\,
            in2 => \N__4103\,
            in3 => \N__4760\,
            lcout => \U111_CYCLE_SM.TS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7752\,
            ce => 'H',
            sr => \N__7691\
        );

    \U111_CYCLE_SM.FLIP_WORD_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011101110"
        )
    port map (
            in0 => \N__6789\,
            in1 => \N__5313\,
            in2 => \N__4085\,
            in3 => \N__6470\,
            lcout => \U111_CYCLE_SM.FLIP_WORDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7752\,
            ce => 'H',
            sr => \N__7691\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4073\,
            in1 => \N__4051\,
            in2 => \_gnd_net_\,
            in3 => \N__6791\,
            lcout => \un1_D_UM_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK40_THRU_LUT4_0_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7757\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_CLK40_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_DIS_RNO_0_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6436\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6500\,
            lcout => \U111_CYCLE_SM.PORT_MISMATCH_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_2_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5266\,
            in2 => \_gnd_net_\,
            in3 => \N__7496\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.N_123_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010001"
        )
    port map (
            in0 => \N__7805\,
            in1 => \N__5349\,
            in2 => \N__4769\,
            in3 => \N__7443\,
            lcout => \U111_CYCLE_SM.N_121_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNISO2G_3_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__7806\,
            in1 => \N__7921\,
            in2 => \_gnd_net_\,
            in3 => \N__5306\,
            lcout => \U111_CYCLE_SM.un1_CYCLE_STATE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__7922\,
            in1 => \N__7811\,
            in2 => \N__7872\,
            in3 => \N__4461\,
            lcout => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7743\,
            ce => 'H',
            sr => \N__7684\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIUBHI_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4462\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5442\,
            lcout => \D_UU_040_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTO81_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__5657\,
            in1 => \N__4457\,
            in2 => \_gnd_net_\,
            in3 => \N__6328\,
            lcout => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81\,
            ltout => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNIGTOZ0Z81_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNI0BVS1_2_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__6329\,
            in1 => \_gnd_net_\,
            in2 => \N__4439\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5903\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7738\,
            ce => \N__6302\,
            sr => \N__6245\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_2_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5524\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7738\,
            ce => \N__6302\,
            sr => \N__6245\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4837\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7738\,
            ce => \N__6302\,
            sr => \N__6245\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_6_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5000\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7738\,
            ce => \N__6302\,
            sr => \N__6245\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_7_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5192\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7738\,
            ce => \N__6302\,
            sr => \N__6245\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_0_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4936\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7738\,
            ce => \N__6302\,
            sr => \N__6245\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNI867Q_6_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7171\,
            in1 => \N__5009\,
            in2 => \_gnd_net_\,
            in3 => \N__4999\,
            lcout => \un1_D_UU_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNISP6Q_0_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4935\,
            in1 => \N__4907\,
            in2 => \_gnd_net_\,
            in3 => \N__7172\,
            lcout => \un1_D_UU_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNI0U6Q_2_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7192\,
            in1 => \N__4877\,
            in2 => \_gnd_net_\,
            in3 => \N__5511\,
            lcout => \un1_D_UU_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7191\,
            in1 => \N__4853\,
            in2 => \_gnd_net_\,
            in3 => \N__4824\,
            lcout => \un1_D_UM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNIA87Q_7_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7193\,
            in1 => \N__5204\,
            in2 => \_gnd_net_\,
            in3 => \N__5191\,
            lcout => \un1_D_UU_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7406\,
            in1 => \N__5129\,
            in2 => \_gnd_net_\,
            in3 => \N__6915\,
            lcout => \un1_D_LL_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6916\,
            in1 => \N__6203\,
            in2 => \_gnd_net_\,
            in3 => \N__5087\,
            lcout => \un1_D_LL_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A2_EN_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__5035\,
            in1 => \N__5024\,
            in2 => \_gnd_net_\,
            in3 => \N__5314\,
            lcout => \U111_CYCLE_SM.A2_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7750\,
            ce => 'H',
            sr => \N__7699\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__7541\,
            in1 => \N__5264\,
            in2 => \_gnd_net_\,
            in3 => \N__5350\,
            lcout => \U111_CYCLE_SM.N_148\,
            ltout => \U111_CYCLE_SM.N_148_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_1_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__7585\,
            in1 => \N__6352\,
            in2 => \N__5018\,
            in3 => \N__5639\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7744\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_1_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__5304\,
            in1 => \N__6463\,
            in2 => \N__5462\,
            in3 => \N__7584\,
            lcout => \U111_CYCLE_SM.TS_EN_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_4_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5640\,
            in2 => \_gnd_net_\,
            in3 => \N__5305\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7744\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5265\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7542\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_srsts_i_o2_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_5_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__5461\,
            in1 => \N__5641\,
            in2 => \N__5450\,
            in3 => \N__5351\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7744\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNITIC9_0_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7916\,
            in2 => \_gnd_net_\,
            in3 => \N__7807\,
            lcout => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5348\,
            in2 => \_gnd_net_\,
            in3 => \N__7444\,
            lcout => \U111_CYCLE_SM.N_128_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__5432\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5393\,
            lcout => \TAn_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_3_0_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__7543\,
            in1 => \N__5347\,
            in2 => \_gnd_net_\,
            in3 => \N__7582\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.N_135_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001010"
        )
    port map (
            in0 => \N__5655\,
            in1 => \N__7917\,
            in2 => \N__5327\,
            in3 => \N__7808\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_srsts_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100011111"
        )
    port map (
            in0 => \N__5267\,
            in1 => \N__5324\,
            in2 => \N__5318\,
            in3 => \N__7418\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7741\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_3_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5654\,
            in1 => \N__6330\,
            in2 => \_gnd_net_\,
            in3 => \N__7472\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7741\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__7544\,
            in1 => \N__5268\,
            in2 => \_gnd_net_\,
            in3 => \N__7441\,
            lcout => \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110101011111"
        )
    port map (
            in0 => \N__5269\,
            in1 => \N__7470\,
            in2 => \N__7552\,
            in3 => \N__7559\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_srsts_i_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_2_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010001000"
        )
    port map (
            in0 => \N__5656\,
            in1 => \N__6477\,
            in2 => \N__5591\,
            in3 => \N__7442\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7739\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5588\,
            lcout => \GB_BUFFER_CLK80_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5537\,
            in1 => \N__5525\,
            in2 => \_gnd_net_\,
            in3 => \N__6846\,
            lcout => \un1_D_LM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7398\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7737\,
            ce => \N__6295\,
            sr => \N__6244\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7263\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7736\,
            ce => \N__6308\,
            sr => \N__6248\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_4_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6562\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7736\,
            ce => \N__6308\,
            sr => \N__6248\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_5_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6728\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7736\,
            ce => \N__6308\,
            sr => \N__6248\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6052\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7736\,
            ce => \N__6308\,
            sr => \N__6248\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_3_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6118\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7736\,
            ce => \N__6308\,
            sr => \N__6248\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6193\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7736\,
            ce => \N__6308\,
            sr => \N__6248\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6186\,
            in1 => \N__6158\,
            in2 => \_gnd_net_\,
            in3 => \N__7207\,
            lcout => \un1_D_UM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNI207Q_3_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6128\,
            in1 => \N__6108\,
            in2 => \_gnd_net_\,
            in3 => \N__7208\,
            lcout => \un1_D_UU_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7209\,
            in1 => \N__6062\,
            in2 => \_gnd_net_\,
            in3 => \N__6045\,
            lcout => \un1_D_UM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5981\,
            in1 => \N__5956\,
            in2 => \_gnd_net_\,
            in3 => \N__6949\,
            lcout => \un1_D_UM_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5892\,
            in1 => \N__5855\,
            in2 => \_gnd_net_\,
            in3 => \N__7218\,
            lcout => \un1_D_UM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6932\,
            in1 => \N__5819\,
            in2 => \_gnd_net_\,
            in3 => \N__5798\,
            lcout => \un1_D_UM_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5732\,
            in1 => \N__5701\,
            in2 => \_gnd_net_\,
            in3 => \N__6933\,
            lcout => \un1_D_UM_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNI647Q_5_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7220\,
            in1 => \N__6737\,
            in2 => \_gnd_net_\,
            in3 => \N__6717\,
            lcout => \un1_D_UU_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6655\,
            in1 => \N__6934\,
            in2 => \_gnd_net_\,
            in3 => \N__6614\,
            lcout => \un1_D_UU_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNI427Q_4_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7219\,
            in1 => \N__6572\,
            in2 => \_gnd_net_\,
            in3 => \N__6549\,
            lcout => \un1_D_UU_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.BURST_COUNT_1_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001010"
        )
    port map (
            in0 => \N__7649\,
            in1 => \N__7637\,
            in2 => \N__6359\,
            in3 => \N__6332\,
            lcout => \U111_CYCLE_SM.BURST_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7749\,
            ce => 'H',
            sr => \N__7700\
        );

    \U111_CYCLE_SM.LW_TRANS_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__6379\,
            in1 => \N__6498\,
            in2 => \N__6401\,
            in3 => \N__6358\,
            lcout => \U111_CYCLE_SM.LW_TRANSZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7749\,
            ce => 'H',
            sr => \N__7700\
        );

    \U111_CYCLE_SM.PORT_MISMATCH_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__6499\,
            in1 => \N__7471\,
            in2 => \N__6482\,
            in3 => \N__6437\,
            lcout => \U111_CYCLE_SM.PORT_MISMATCHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7749\,
            ce => 'H',
            sr => \N__7700\
        );

    \U111_CYCLE_SM.BURST_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__6397\,
            in1 => \N__6357\,
            in2 => \N__6380\,
            in3 => \N__7586\,
            lcout => \U111_CYCLE_SM.BURSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7749\,
            ce => 'H',
            sr => \N__7700\
        );

    \U111_CYCLE_SM.BURST_COUNT_0_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6353\,
            in1 => \N__7636\,
            in2 => \_gnd_net_\,
            in3 => \N__6331\,
            lcout => \U111_CYCLE_SM.BURST_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7749\,
            ce => 'H',
            sr => \N__7700\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001100"
        )
    port map (
            in0 => \N__7915\,
            in1 => \N__7768\,
            in2 => \N__7873\,
            in3 => \N__7810\,
            lcout => \U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7749\,
            ce => 'H',
            sr => \N__7700\
        );

    \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__7648\,
            in1 => \N__7635\,
            in2 => \N__7622\,
            in3 => \N__7583\,
            lcout => \U111_CYCLE_SM.un7_CYCLE_STATE_0\,
            ltout => \U111_CYCLE_SM.un7_CYCLE_STATE_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__7548\,
            in1 => \N__7469\,
            in2 => \N__7448\,
            in3 => \N__7445\,
            lcout => \U111_CYCLE_SM.N_136\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7412\,
            in1 => \N__7399\,
            in2 => \_gnd_net_\,
            in3 => \N__7189\,
            lcout => \un1_D_UM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__7352\,
            in1 => \N__6921\,
            in2 => \_gnd_net_\,
            in3 => \N__7333\,
            lcout => \un1_D_UM_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7264\,
            in1 => \N__7226\,
            in2 => \_gnd_net_\,
            in3 => \N__7190\,
            lcout => \un1_D_UM_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__7082\,
            in1 => \N__6956\,
            in2 => \_gnd_net_\,
            in3 => \N__7060\,
            lcout => \un1_D_UU_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6991\,
            in1 => \N__6955\,
            in2 => \_gnd_net_\,
            in3 => \N__7961\,
            lcout => \un1_D_UU_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

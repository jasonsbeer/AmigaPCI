-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 14 2024 10:36:48

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U111_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U111_TOP
entity U111_TOP is
port (
    D_LL_AMIGA : inout std_logic_vector(7 downto 0);
    D_LM_AMIGA : inout std_logic_vector(7 downto 0);
    D_UU_AMIGA : inout std_logic_vector(7 downto 0);
    D_UM_AMIGA : inout std_logic_vector(7 downto 0);
    D_UU_040 : inout std_logic_vector(7 downto 0);
    D_LL_040 : inout std_logic_vector(7 downto 0);
    D_LM_040 : inout std_logic_vector(7 downto 0);
    D_UM_040 : inout std_logic_vector(7 downto 0);
    A_AMIGA : out std_logic_vector(1 downto 0);
    A_040 : in std_logic_vector(1 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    TSn : out std_logic;
    RESETn : in std_logic;
    CLKRAMA : out std_logic;
    PORTSIZE : in std_logic;
    CLK40B : out std_logic;
    TBI_CPUn : out std_logic;
    TAn : out std_logic;
    CPUBGn : out std_logic;
    BUFENn : out std_logic;
    RnW : in std_logic;
    CLK80_CPU : out std_logic;
    BUFDIR : out std_logic;
    TCI_CPUn : out std_logic;
    TS_CPUn : in std_logic;
    CLKRAMB : out std_logic;
    CLK40A : out std_logic;
    DMAn : out std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    TACKn : in std_logic;
    BGn : in std_logic);
end U111_TOP;

-- Architecture of U111_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U111_TOP is

signal \N__7843\ : std_logic;
signal \N__7827\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7260\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4018\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4012\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3938\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3779\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3760\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3622\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3618\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3587\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3548\ : std_logic;
signal \N__3545\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3482\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3476\ : std_logic;
signal \N__3473\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3442\ : std_logic;
signal \N__3439\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3404\ : std_logic;
signal \N__3401\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3392\ : std_logic;
signal \N__3389\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3383\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3353\ : std_logic;
signal \N__3350\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3263\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3254\ : std_logic;
signal \N__3251\ : std_logic;
signal \N__3248\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3209\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3176\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3056\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2987\ : std_logic;
signal \N__2984\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2951\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2875\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2863\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2854\ : std_logic;
signal \N__2851\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2845\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2794\ : std_logic;
signal \N__2791\ : std_logic;
signal \N__2788\ : std_logic;
signal \N__2785\ : std_logic;
signal \N__2782\ : std_logic;
signal \N__2779\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2747\ : std_logic;
signal \N__2744\ : std_logic;
signal \N__2741\ : std_logic;
signal \N__2738\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2705\ : std_logic;
signal \N__2702\ : std_logic;
signal \N__2699\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2672\ : std_logic;
signal \N__2669\ : std_logic;
signal \N__2666\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2639\ : std_logic;
signal \N__2636\ : std_logic;
signal \N__2635\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2617\ : std_logic;
signal \N__2614\ : std_logic;
signal \N__2611\ : std_logic;
signal \N__2608\ : std_logic;
signal \N__2605\ : std_logic;
signal \N__2600\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2579\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2546\ : std_logic;
signal \N__2543\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2524\ : std_logic;
signal \N__2523\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2521\ : std_logic;
signal \N__2520\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2518\ : std_logic;
signal \N__2517\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2515\ : std_logic;
signal \N__2512\ : std_logic;
signal \N__2509\ : std_logic;
signal \N__2506\ : std_logic;
signal \N__2503\ : std_logic;
signal \N__2502\ : std_logic;
signal \N__2501\ : std_logic;
signal \N__2500\ : std_logic;
signal \N__2499\ : std_logic;
signal \N__2496\ : std_logic;
signal \N__2493\ : std_logic;
signal \N__2490\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2488\ : std_logic;
signal \N__2487\ : std_logic;
signal \N__2484\ : std_logic;
signal \N__2481\ : std_logic;
signal \N__2478\ : std_logic;
signal \N__2475\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2463\ : std_logic;
signal \N__2460\ : std_logic;
signal \N__2457\ : std_logic;
signal \N__2454\ : std_logic;
signal \N__2453\ : std_logic;
signal \N__2452\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2450\ : std_logic;
signal \N__2443\ : std_logic;
signal \N__2440\ : std_logic;
signal \N__2437\ : std_logic;
signal \N__2434\ : std_logic;
signal \N__2425\ : std_logic;
signal \N__2424\ : std_logic;
signal \N__2423\ : std_logic;
signal \N__2412\ : std_logic;
signal \N__2409\ : std_logic;
signal \N__2406\ : std_logic;
signal \N__2403\ : std_logic;
signal \N__2400\ : std_logic;
signal \N__2399\ : std_logic;
signal \N__2398\ : std_logic;
signal \N__2397\ : std_logic;
signal \N__2396\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2384\ : std_logic;
signal \N__2381\ : std_logic;
signal \N__2378\ : std_logic;
signal \N__2367\ : std_logic;
signal \N__2364\ : std_logic;
signal \N__2361\ : std_logic;
signal \N__2358\ : std_logic;
signal \N__2355\ : std_logic;
signal \N__2352\ : std_logic;
signal \N__2351\ : std_logic;
signal \N__2350\ : std_logic;
signal \N__2347\ : std_logic;
signal \N__2342\ : std_logic;
signal \N__2333\ : std_logic;
signal \N__2332\ : std_logic;
signal \N__2331\ : std_logic;
signal \N__2328\ : std_logic;
signal \N__2325\ : std_logic;
signal \N__2322\ : std_logic;
signal \N__2319\ : std_logic;
signal \N__2314\ : std_logic;
signal \N__2311\ : std_logic;
signal \N__2308\ : std_logic;
signal \N__2305\ : std_logic;
signal \N__2302\ : std_logic;
signal \N__2299\ : std_logic;
signal \N__2294\ : std_logic;
signal \N__2289\ : std_logic;
signal \N__2286\ : std_logic;
signal \N__2283\ : std_logic;
signal \N__2280\ : std_logic;
signal \N__2275\ : std_logic;
signal \N__2272\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2258\ : std_logic;
signal \N__2255\ : std_logic;
signal \N__2252\ : std_logic;
signal \N__2249\ : std_logic;
signal \N__2246\ : std_logic;
signal \N__2243\ : std_logic;
signal \N__2240\ : std_logic;
signal \N__2237\ : std_logic;
signal \N__2234\ : std_logic;
signal \N__2231\ : std_logic;
signal \N__2228\ : std_logic;
signal \N__2225\ : std_logic;
signal \N__2222\ : std_logic;
signal \N__2219\ : std_logic;
signal \N__2216\ : std_logic;
signal \N__2215\ : std_logic;
signal \N__2212\ : std_logic;
signal \N__2209\ : std_logic;
signal \N__2206\ : std_logic;
signal \N__2203\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \A_040_c_0\ : std_logic;
signal \A_AMIGA_c_0\ : std_logic;
signal \A_040_c_1\ : std_logic;
signal \RnW_c_i_0\ : std_logic;
signal \D_LL_AMIGA_in_3\ : std_logic;
signal \un1_D_LL_AMIGA_3\ : std_logic;
signal \A_AMIGA_c_1\ : std_logic;
signal \D_LL_AMIGA_in_7\ : std_logic;
signal \un1_D_LL_AMIGA_7\ : std_logic;
signal \D_LM_AMIGA_in_0\ : std_logic;
signal \un1_D_LM_AMIGA_0\ : std_logic;
signal \D_LM_AMIGA_in_6\ : std_logic;
signal \un1_D_LM_AMIGA_6\ : std_logic;
signal \D_LM_040_in_3\ : std_logic;
signal \D_UU_040_in_3\ : std_logic;
signal \un1_D_UU_040_3\ : std_logic;
signal \D_LM_040_in_2\ : std_logic;
signal \D_UU_040_in_2\ : std_logic;
signal \un1_D_UU_040_2\ : std_logic;
signal \D_LL_AMIGA_in_0\ : std_logic;
signal \un1_D_LL_AMIGA_0\ : std_logic;
signal \D_LL_AMIGA_in_4\ : std_logic;
signal \un1_D_LL_AMIGA_4\ : std_logic;
signal \D_LL_040_in_2\ : std_logic;
signal \D_UM_040_in_2\ : std_logic;
signal \un1_D_UM_040_2\ : std_logic;
signal \D_LM_AMIGA_in_2\ : std_logic;
signal \un1_D_LM_AMIGA_2\ : std_logic;
signal \D_LM_040_in_7\ : std_logic;
signal \D_UU_040_in_7\ : std_logic;
signal \un1_D_UU_040_7\ : std_logic;
signal \D_LL_AMIGA_in_5\ : std_logic;
signal \un1_D_LL_AMIGA_5\ : std_logic;
signal \D_LM_AMIGA_in_1\ : std_logic;
signal \un1_D_LM_AMIGA_1\ : std_logic;
signal \D_LM_AMIGA_in_3\ : std_logic;
signal \un1_D_LM_AMIGA_3\ : std_logic;
signal \D_UM_040_in_6\ : std_logic;
signal \D_LL_040_in_6\ : std_logic;
signal \un1_D_UM_040_6\ : std_logic;
signal \D_LM_AMIGA_in_5\ : std_logic;
signal \un1_D_LM_AMIGA_5\ : std_logic;
signal \D_UU_040_in_5\ : std_logic;
signal \D_LM_040_in_5\ : std_logic;
signal \un1_D_UU_040_5\ : std_logic;
signal \INVU111_CYCLE_SM.TA_EN_nessC_net\ : std_logic;
signal \INVU111_CYCLE_SM.TSnC_net\ : std_logic;
signal \D_UM_040_in_4\ : std_logic;
signal \D_LL_040_in_4\ : std_logic;
signal \un1_D_UM_040_4\ : std_logic;
signal \D_LL_AMIGA_in_1\ : std_logic;
signal \un1_D_LL_AMIGA_1\ : std_logic;
signal \U111_CYCLE_SM.A_OUTZ0\ : std_logic;
signal \INVU111_CYCLE_SM.A_OUTC_net\ : std_logic;
signal \U111_CYCLE_SM.un1_CYCLE_STATE_1_0\ : std_logic;
signal \U111_CYCLE_SM.un1_CYCLE_STATE_1_0_cascade_\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U111_CYCLE_SM.un1_CYCLE_STATE_1_0_0\ : std_logic;
signal \U111_CYCLE_SM.TA_ENZ0\ : std_logic;
signal \TAn_0_i\ : std_logic;
signal \D_LM_AMIGA_in_4\ : std_logic;
signal \un1_D_LM_AMIGA_4\ : std_logic;
signal \U111_CYCLE_SM.TS_EN10_cascade_\ : std_logic;
signal \U111_CYCLE_SM.TS_ENZ0\ : std_logic;
signal \U111_CYCLE_SM.LW_CYCLE_r_1_cascade_\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U111_CYCLE_SM.LW_CYCLE_STARTZ0\ : std_logic;
signal \INVU111_CYCLE_SM.TS_ENC_net\ : std_logic;
signal \INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\ : std_logic;
signal \D_UU_AMIGA_in_6\ : std_logic;
signal \un1_D_UU_AMIGA_6\ : std_logic;
signal \D_UU_040_in_0\ : std_logic;
signal \D_LM_040_in_0\ : std_logic;
signal \un1_D_UU_040_0\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\ : std_logic;
signal \D_UU_AMIGA_in_4\ : std_logic;
signal \un1_D_UU_AMIGA_4\ : std_logic;
signal \D_LL_040_in_0\ : std_logic;
signal \D_UM_040_in_0\ : std_logic;
signal \un1_D_UM_040_0\ : std_logic;
signal \GB_BUFFER_CLK40_THRU_CO\ : std_logic;
signal \un1_D_UM_AMIGA_0\ : std_logic;
signal \D_UM_AMIGA_in_0\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\ : std_logic;
signal \INVU111_CYCLE_SM.UM_LATCHED_nesr_0C_net\ : std_logic;
signal \INVU111_CYCLE_SM.CYCLE_STATE_1C_net\ : std_logic;
signal \CLK40\ : std_logic;
signal \TS_CPUn_c\ : std_logic;
signal \U111_CYCLE_SM.TS_EN_4\ : std_logic;
signal \TACKn_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0_cascade_\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa\ : std_logic;
signal \INVU111_CYCLE_SM.UU_LATCHED_nesr_0C_net\ : std_logic;
signal \D_LM_AMIGA_in_7\ : std_logic;
signal \un1_D_LM_AMIGA_7\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\ : std_logic;
signal \D_UM_AMIGA_in_4\ : std_logic;
signal \un1_D_UM_AMIGA_4\ : std_logic;
signal \D_LL_040_in_5\ : std_logic;
signal \D_UM_040_in_5\ : std_logic;
signal \un1_D_UM_040_5\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\ : std_logic;
signal \D_UU_AMIGA_in_0\ : std_logic;
signal \un1_D_UU_AMIGA_0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \D_LL_AMIGA_in_2\ : std_logic;
signal \un1_D_LL_AMIGA_2\ : std_logic;
signal \D_LL_AMIGA_in_6\ : std_logic;
signal \un1_D_LL_AMIGA_6\ : std_logic;
signal \un1_D_UM_AMIGA_2\ : std_logic;
signal \CLK80\ : std_logic;
signal \GB_BUFFER_CLK80_THRU_CO\ : std_logic;
signal \D_UM_AMIGA_in_2\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\ : std_logic;
signal \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net\ : std_logic;
signal \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\ : std_logic;
signal \INVU111_CYCLE_SM.UU_LATCHED_nesr_7C_net\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0\ : std_logic;
signal \D_UM_AMIGA_in_1\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\ : std_logic;
signal \un1_D_UM_AMIGA_1\ : std_logic;
signal \D_UM_AMIGA_in_3\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\ : std_logic;
signal \un1_D_UM_AMIGA_3\ : std_logic;
signal \D_LL_040_in_3\ : std_logic;
signal \D_UM_040_in_3\ : std_logic;
signal \un1_D_UM_040_3\ : std_logic;
signal \D_UM_AMIGA_in_7\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\ : std_logic;
signal \un1_D_UM_AMIGA_7\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\ : std_logic;
signal \D_UU_AMIGA_in_2\ : std_logic;
signal \un1_D_UU_AMIGA_2\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\ : std_logic;
signal \D_UU_AMIGA_in_5\ : std_logic;
signal \un1_D_UU_AMIGA_5\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\ : std_logic;
signal \D_UU_AMIGA_in_3\ : std_logic;
signal \un1_D_UU_AMIGA_3\ : std_logic;
signal \D_UU_040_in_6\ : std_logic;
signal \D_LM_040_in_6\ : std_logic;
signal \un1_D_UU_040_6\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\ : std_logic;
signal \D_UM_AMIGA_in_5\ : std_logic;
signal \un1_D_UM_AMIGA_5\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\ : std_logic;
signal \D_UU_AMIGA_in_7\ : std_logic;
signal \un1_D_UU_AMIGA_7\ : std_logic;
signal \D_UM_AMIGA_in_6\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\ : std_logic;
signal \un1_D_UM_AMIGA_6\ : std_logic;
signal \D_LL_040_in_1\ : std_logic;
signal \D_UM_040_in_1\ : std_logic;
signal \un1_D_UM_040_1\ : std_logic;
signal \U111_CYCLE_SM.LW_CYCLEZ0\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\ : std_logic;
signal \D_UU_AMIGA_in_1\ : std_logic;
signal \un1_D_UU_AMIGA_1\ : std_logic;
signal \D_LM_040_in_1\ : std_logic;
signal \D_UU_040_in_1\ : std_logic;
signal \un1_D_UU_040_1\ : std_logic;
signal \D_LL_040_in_7\ : std_logic;
signal \D_UM_040_in_7\ : std_logic;
signal \un1_D_UM_040_7\ : std_logic;
signal \D_LM_040_in_4\ : std_logic;
signal \D_UU_040_in_4\ : std_logic;
signal \U111_CYCLE_SM.FLIP\ : std_logic;
signal \un1_D_UU_040_4\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \PORTSIZE_c\ : std_logic;
signal \U111_CYCLE_SM.LW_TRANS_0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK40_IN_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \CPUBGn_wire\ : std_logic;
signal \A_040_wire\ : std_logic_vector(1 downto 0);
signal \A_AMIGA_wire\ : std_logic_vector(1 downto 0);
signal \CLK40B_wire\ : std_logic;
signal \TBI_CPUn_wire\ : std_logic;
signal \CLK40A_wire\ : std_logic;
signal \BUFDIR_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \TS_CPUn_wire\ : std_logic;
signal \CLKRAMA_wire\ : std_logic;
signal \TCI_CPUn_wire\ : std_logic;
signal \CLKRAMB_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \TAn_wire\ : std_logic;
signal \DMAn_wire\ : std_logic;
signal \CLK80_CPU_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \pll_pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK40_IN_wire\ <= CLK40_IN;
    \TACKn_wire\ <= TACKn;
    CPUBGn <= \CPUBGn_wire\;
    \A_040_wire\ <= A_040;
    A_AMIGA <= \A_AMIGA_wire\;
    CLK40B <= \CLK40B_wire\;
    TBI_CPUn <= \TBI_CPUn_wire\;
    CLK40A <= \CLK40A_wire\;
    BUFDIR <= \BUFDIR_wire\;
    \SIZ_wire\ <= SIZ;
    \TS_CPUn_wire\ <= TS_CPUn;
    CLKRAMA <= \CLKRAMA_wire\;
    TCI_CPUn <= \TCI_CPUn_wire\;
    CLKRAMB <= \CLKRAMB_wire\;
    BUFENn <= \BUFENn_wire\;
    \RnW_wire\ <= RnW;
    TAn <= \TAn_wire\;
    DMAn <= \DMAn_wire\;
    CLK80_CPU <= \CLK80_CPU_wire\;
    TSn <= \TSn_wire\;
    \PORTSIZE_wire\ <= PORTSIZE;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    \pll_pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll_pll\ : PLL40_2F
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            SCLK => '0',
            PLLOUTGLOBALA => \CLK80\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALB => \CLK40\,
            SDI => '0',
            PLLOUTCOREA => OPEN,
            BYPASS => '0',
            RESETB => \N__5041\,
            PLLOUTCOREB => OPEN,
            LOCK => OPEN,
            SDO => OPEN,
            EXTFEEDBACK => '0',
            DYNAMICDELAY => \pll_pll_DYNAMICDELAY_wire\,
            PLLIN => \N__7843\
        );

    \pll_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \VCCG0\,
            DIN => '0',
            DOUT => \N__7843\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \D_UM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7827\,
            DIN => \N__7826\,
            DOUT => \N__7825\,
            PACKAGEPIN => D_UM_040(3)
        );

    \D_UM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7827\,
            PADOUT => \N__7826\,
            PADIN => \N__7825\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4494\,
            DIN0 => \D_UM_040_in_3\,
            DOUT0 => \N__5804\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7818\,
            DIN => \N__7817\,
            DOUT => \N__7816\,
            PACKAGEPIN => D_LL_AMIGA(1)
        );

    \D_LL_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7818\,
            PADOUT => \N__7817\,
            PADIN => \N__7816\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2516\,
            DIN0 => \D_LL_AMIGA_in_1\,
            DOUT0 => \N__6725\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7809\,
            DIN => \N__7808\,
            DOUT => \N__7807\,
            PACKAGEPIN => D_UU_AMIGA(5)
        );

    \D_UU_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7809\,
            PADOUT => \N__7808\,
            PADIN => \N__7807\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2525\,
            DIN0 => \D_UU_AMIGA_in_5\,
            DOUT0 => \N__2999\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7800\,
            DIN => \N__7799\,
            DOUT => \N__7798\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7800\,
            PADOUT => \N__7799\,
            PADIN => \N__7798\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TACKn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7791\,
            DIN => \N__7790\,
            DOUT => \N__7789\,
            PACKAGEPIN => D_UU_040(6)
        );

    \D_UU_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7791\,
            PADOUT => \N__7790\,
            PADIN => \N__7789\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4550\,
            DIN0 => \D_UU_040_in_6\,
            DOUT0 => \N__3590\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CPUBGn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7782\,
            DIN => \N__7781\,
            DOUT => \N__7780\,
            PACKAGEPIN => \CPUBGn_wire\
        );

    \CPUBGn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7782\,
            PADOUT => \N__7781\,
            PADIN => \N__7780\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7773\,
            DIN => \N__7772\,
            DOUT => \N__7771\,
            PACKAGEPIN => D_LL_040(7)
        );

    \D_LL_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7773\,
            PADOUT => \N__7772\,
            PADIN => \N__7771\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4591\,
            DIN0 => \D_LL_040_in_7\,
            DOUT0 => \N__2969\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7764\,
            DIN => \N__7763\,
            DOUT => \N__7762\,
            PACKAGEPIN => D_LL_AMIGA(4)
        );

    \D_LL_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7764\,
            PADOUT => \N__7763\,
            PADIN => \N__7762\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2515\,
            DIN0 => \D_LL_AMIGA_in_4\,
            DOUT0 => \N__3548\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7755\,
            DIN => \N__7754\,
            DOUT => \N__7753\,
            PACKAGEPIN => D_UM_AMIGA(3)
        );

    \D_UM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7755\,
            PADOUT => \N__7754\,
            PADIN => \N__7753\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2502\,
            DIN0 => \D_UM_AMIGA_in_3\,
            DOUT0 => \N__5720\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7746\,
            DIN => \N__7745\,
            DOUT => \N__7744\,
            PACKAGEPIN => D_UU_040(3)
        );

    \D_UU_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7746\,
            PADOUT => \N__7745\,
            PADIN => \N__7744\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4545\,
            DIN0 => \D_UU_040_in_3\,
            DOUT0 => \N__5414\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7737\,
            DIN => \N__7736\,
            DOUT => \N__7735\,
            PACKAGEPIN => \A_040_wire\(1)
        );

    \A_040_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7737\,
            PADOUT => \N__7736\,
            PADIN => \N__7735\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7728\,
            DIN => \N__7727\,
            DOUT => \N__7726\,
            PACKAGEPIN => D_LM_AMIGA(3)
        );

    \D_LM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7728\,
            PADOUT => \N__7727\,
            PADIN => \N__7726\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2397\,
            DIN0 => \D_LM_AMIGA_in_3\,
            DOUT0 => \N__2885\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7719\,
            DIN => \N__7718\,
            DOUT => \N__7717\,
            PACKAGEPIN => D_LM_040(0)
        );

    \D_LM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7719\,
            PADOUT => \N__7718\,
            PADIN => \N__7717\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4592\,
            DIN0 => \D_LM_040_in_0\,
            DOUT0 => \N__2933\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7710\,
            DIN => \N__7709\,
            DOUT => \N__7708\,
            PACKAGEPIN => D_UM_AMIGA(6)
        );

    \D_UM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7710\,
            PADOUT => \N__7709\,
            PADIN => \N__7708\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2524\,
            DIN0 => \D_UM_AMIGA_in_6\,
            DOUT0 => \N__3113\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7701\,
            DIN => \N__7700\,
            DOUT => \N__7699\,
            PACKAGEPIN => D_LM_AMIGA(4)
        );

    \D_LM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7701\,
            PADOUT => \N__7700\,
            PADIN => \N__7699\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2450\,
            DIN0 => \D_LM_AMIGA_in_4\,
            DOUT0 => \N__6218\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7692\,
            DIN => \N__7691\,
            DOUT => \N__7690\,
            PACKAGEPIN => \A_AMIGA_wire\(1)
        );

    \A_AMIGA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7692\,
            PADOUT => \N__7691\,
            PADIN => \N__7690\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2215\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7683\,
            DIN => \N__7682\,
            DOUT => \N__7681\,
            PACKAGEPIN => D_LM_040(7)
        );

    \D_LM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7683\,
            PADOUT => \N__7682\,
            PADIN => \N__7681\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4413\,
            DIN0 => \D_LM_040_in_7\,
            DOUT0 => \N__4220\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7674\,
            DIN => \N__7673\,
            DOUT => \N__7672\,
            PACKAGEPIN => D_UM_040(4)
        );

    \D_UM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7674\,
            PADOUT => \N__7673\,
            PADIN => \N__7672\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4546\,
            DIN0 => \D_UM_040_in_4\,
            DOUT0 => \N__4145\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7665\,
            DIN => \N__7664\,
            DOUT => \N__7663\,
            PACKAGEPIN => \CLK40B_wire\
        );

    \CLK40B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7665\,
            PADOUT => \N__7664\,
            PADIN => \N__7663\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3841\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7656\,
            DIN => \N__7655\,
            DOUT => \N__7654\,
            PACKAGEPIN => D_UU_AMIGA(0)
        );

    \D_UU_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7656\,
            PADOUT => \N__7655\,
            PADIN => \N__7654\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2489\,
            DIN0 => \D_UU_AMIGA_in_0\,
            DOUT0 => \N__4001\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7647\,
            DIN => \N__7646\,
            DOUT => \N__7645\,
            PACKAGEPIN => \A_040_wire\(0)
        );

    \A_040_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7647\,
            PADOUT => \N__7646\,
            PADIN => \N__7645\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7638\,
            DIN => \N__7637\,
            DOUT => \N__7636\,
            PACKAGEPIN => D_LM_AMIGA(0)
        );

    \D_LM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7638\,
            PADOUT => \N__7637\,
            PADIN => \N__7636\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2351\,
            DIN0 => \D_LM_AMIGA_in_0\,
            DOUT0 => \N__4049\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7629\,
            DIN => \N__7628\,
            DOUT => \N__7627\,
            PACKAGEPIN => D_UM_040(1)
        );

    \D_UM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7629\,
            PADOUT => \N__7628\,
            PADIN => \N__7627\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4492\,
            DIN0 => \D_UM_040_in_1\,
            DOUT0 => \N__5153\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7620\,
            DIN => \N__7619\,
            DOUT => \N__7618\,
            PACKAGEPIN => \TBI_CPUn_wire\
        );

    \TBI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7620\,
            PADOUT => \N__7619\,
            PADIN => \N__7618\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7611\,
            DIN => \N__7610\,
            DOUT => \N__7609\,
            PACKAGEPIN => \CLK40A_wire\
        );

    \CLK40A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7611\,
            PADOUT => \N__7610\,
            PADIN => \N__7609\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3842\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7602\,
            DIN => \N__7601\,
            DOUT => \N__7600\,
            PACKAGEPIN => D_LM_040(3)
        );

    \D_LM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7602\,
            PADOUT => \N__7601\,
            PADIN => \N__7600\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4557\,
            DIN0 => \D_LM_040_in_3\,
            DOUT0 => \N__3188\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7593\,
            DIN => \N__7592\,
            DOUT => \N__7591\,
            PACKAGEPIN => D_LL_040(4)
        );

    \D_LL_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7593\,
            PADOUT => \N__7592\,
            PADIN => \N__7591\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4628\,
            DIN0 => \D_LL_040_in_4\,
            DOUT0 => \N__2663\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7584\,
            DIN => \N__7583\,
            DOUT => \N__7582\,
            PACKAGEPIN => D_LL_AMIGA(7)
        );

    \D_LL_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7584\,
            PADOUT => \N__7583\,
            PADIN => \N__7582\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2350\,
            DIN0 => \D_LL_AMIGA_in_7\,
            DOUT0 => \N__6305\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7575\,
            DIN => \N__7574\,
            DOUT => \N__7573\,
            PACKAGEPIN => D_UU_AMIGA(7)
        );

    \D_UU_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7575\,
            PADOUT => \N__7574\,
            PADIN => \N__7573\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2519\,
            DIN0 => \D_UU_AMIGA_in_7\,
            DOUT0 => \N__3293\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7566\,
            DIN => \N__7565\,
            DOUT => \N__7564\,
            PACKAGEPIN => \BUFDIR_wire\
        );

    \BUFDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7566\,
            PADOUT => \N__7565\,
            PADIN => \N__7564\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4631\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7557\,
            DIN => \N__7556\,
            DOUT => \N__7555\,
            PACKAGEPIN => D_LM_AMIGA(5)
        );

    \D_LM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7557\,
            PADOUT => \N__7556\,
            PADIN => \N__7555\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2452\,
            DIN0 => \D_LM_AMIGA_in_5\,
            DOUT0 => \N__3041\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7548\,
            DIN => \N__7547\,
            DOUT => \N__7546\,
            PACKAGEPIN => D_UU_040(4)
        );

    \D_UU_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7548\,
            PADOUT => \N__7547\,
            PADIN => \N__7546\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4588\,
            DIN0 => \D_UU_040_in_4\,
            DOUT0 => \N__3938\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7539\,
            DIN => \N__7538\,
            DOUT => \N__7537\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7539\,
            PADOUT => \N__7538\,
            PADIN => \N__7537\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7530\,
            DIN => \N__7529\,
            DOUT => \N__7528\,
            PACKAGEPIN => D_LM_040(6)
        );

    \D_LM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7530\,
            PADOUT => \N__7529\,
            PADIN => \N__7528\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4405\,
            DIN0 => \D_LM_040_in_6\,
            DOUT0 => \N__2900\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7521\,
            DIN => \N__7520\,
            DOUT => \N__7519\,
            PACKAGEPIN => D_UM_040(5)
        );

    \D_UM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7521\,
            PADOUT => \N__7520\,
            PADIN => \N__7519\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4547\,
            DIN0 => \D_UM_040_in_5\,
            DOUT0 => \N__6866\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TS_CPUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7512\,
            DIN => \N__7511\,
            DOUT => \N__7510\,
            PACKAGEPIN => \TS_CPUn_wire\
        );

    \TS_CPUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7512\,
            PADOUT => \N__7511\,
            PADIN => \N__7510\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TS_CPUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7503\,
            DIN => \N__7502\,
            DOUT => \N__7501\,
            PACKAGEPIN => D_LL_040(1)
        );

    \D_LL_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7503\,
            PADOUT => \N__7502\,
            PADIN => \N__7501\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4627\,
            DIN0 => \D_LL_040_in_1\,
            DOUT0 => \N__3473\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7494\,
            DIN => \N__7493\,
            DOUT => \N__7492\,
            PACKAGEPIN => D_LL_AMIGA(3)
        );

    \D_LL_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7494\,
            PADOUT => \N__7493\,
            PADIN => \N__7492\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2517\,
            DIN0 => \D_LL_AMIGA_in_3\,
            DOUT0 => \N__5782\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7485\,
            DIN => \N__7484\,
            DOUT => \N__7483\,
            PACKAGEPIN => D_UM_AMIGA(5)
        );

    \D_UM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7485\,
            PADOUT => \N__7484\,
            PADIN => \N__7483\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2396\,
            DIN0 => \D_UM_AMIGA_in_5\,
            DOUT0 => \N__5135\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7476\,
            DIN => \N__7475\,
            DOUT => \N__7474\,
            PACKAGEPIN => D_UU_040(1)
        );

    \D_UU_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7476\,
            PADOUT => \N__7475\,
            PADIN => \N__7474\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4495\,
            DIN0 => \D_UU_040_in_1\,
            DOUT0 => \N__6419\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7467\,
            DIN => \N__7466\,
            DOUT => \N__7465\,
            PACKAGEPIN => D_UU_AMIGA(3)
        );

    \D_UU_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7467\,
            PADOUT => \N__7466\,
            PADIN => \N__7465\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2521\,
            DIN0 => \D_UU_AMIGA_in_3\,
            DOUT0 => \N__2816\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7458\,
            DIN => \N__7457\,
            DOUT => \N__7456\,
            PACKAGEPIN => D_LM_AMIGA(1)
        );

    \D_LM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7458\,
            PADOUT => \N__7457\,
            PADIN => \N__7456\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2331\,
            DIN0 => \D_LM_AMIGA_in_1\,
            DOUT0 => \N__6398\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7449\,
            DIN => \N__7448\,
            DOUT => \N__7447\,
            PACKAGEPIN => D_LM_040(2)
        );

    \D_LM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7449\,
            PADOUT => \N__7448\,
            PADIN => \N__7447\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4590\,
            DIN0 => \D_LM_040_in_2\,
            DOUT0 => \N__3365\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7440\,
            DIN => \N__7439\,
            DOUT => \N__7438\,
            PACKAGEPIN => D_LL_040(5)
        );

    \D_LL_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7440\,
            PADOUT => \N__7439\,
            PADIN => \N__7438\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4593\,
            DIN0 => \D_LL_040_in_5\,
            DOUT0 => \N__3257\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7431\,
            DIN => \N__7430\,
            DOUT => \N__7429\,
            PACKAGEPIN => D_LL_AMIGA(6)
        );

    \D_LL_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7431\,
            PADOUT => \N__7430\,
            PADIN => \N__7429\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2423\,
            DIN0 => \D_LL_AMIGA_in_6\,
            DOUT0 => \N__3155\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7422\,
            DIN => \N__7421\,
            DOUT => \N__7420\,
            PACKAGEPIN => D_UU_AMIGA(6)
        );

    \D_UU_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7422\,
            PADOUT => \N__7421\,
            PADIN => \N__7420\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2520\,
            DIN0 => \D_UU_AMIGA_in_6\,
            DOUT0 => \N__5336\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7413\,
            DIN => \N__7412\,
            DOUT => \N__7411\,
            PACKAGEPIN => D_UM_AMIGA(1)
        );

    \D_UM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7413\,
            PADOUT => \N__7412\,
            PADIN => \N__7411\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2453\,
            DIN0 => \D_UM_AMIGA_in_1\,
            DOUT0 => \N__6662\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7404\,
            DIN => \N__7403\,
            DOUT => \N__7402\,
            PACKAGEPIN => D_UU_040(5)
        );

    \D_UU_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7404\,
            PADOUT => \N__7403\,
            PADIN => \N__7402\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4548\,
            DIN0 => \D_UU_040_in_5\,
            DOUT0 => \N__5486\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7395\,
            DIN => \N__7394\,
            DOUT => \N__7393\,
            PACKAGEPIN => \CLKRAMA_wire\
        );

    \CLKRAMA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7395\,
            PADOUT => \N__7394\,
            PADIN => \N__7393\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4889\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7386\,
            DIN => \N__7385\,
            DOUT => \N__7384\,
            PACKAGEPIN => D_UM_040(2)
        );

    \D_UM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7386\,
            PADOUT => \N__7385\,
            PADIN => \N__7384\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4473\,
            DIN0 => \D_UM_040_in_2\,
            DOUT0 => \N__4943\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7377\,
            DIN => \N__7376\,
            DOUT => \N__7375\,
            PACKAGEPIN => D_LL_040(2)
        );

    \D_LL_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7377\,
            PADOUT => \N__7376\,
            PADIN => \N__7375\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4611\,
            DIN0 => \D_LL_040_in_2\,
            DOUT0 => \N__5003\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7368\,
            DIN => \N__7367\,
            DOUT => \N__7366\,
            PACKAGEPIN => \TCI_CPUn_wire\
        );

    \TCI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7368\,
            PADOUT => \N__7367\,
            PADIN => \N__7366\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMB_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7359\,
            DIN => \N__7358\,
            DOUT => \N__7357\,
            PACKAGEPIN => \CLKRAMB_wire\
        );

    \CLKRAMB_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7359\,
            PADOUT => \N__7358\,
            PADIN => \N__7357\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4879\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7350\,
            DIN => \N__7349\,
            DOUT => \N__7348\,
            PACKAGEPIN => D_LL_AMIGA(2)
        );

    \D_LL_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7350\,
            PADOUT => \N__7349\,
            PADIN => \N__7348\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2518\,
            DIN0 => \D_LL_AMIGA_in_2\,
            DOUT0 => \N__2639\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7341\,
            DIN => \N__7340\,
            DOUT => \N__7339\,
            PACKAGEPIN => D_UM_AMIGA(4)
        );

    \D_UM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7341\,
            PADOUT => \N__7340\,
            PADIN => \N__7339\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2523\,
            DIN0 => \D_UM_AMIGA_in_4\,
            DOUT0 => \N__3512\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7332\,
            DIN => \N__7331\,
            DOUT => \N__7330\,
            PACKAGEPIN => D_UU_AMIGA(2)
        );

    \D_UU_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7332\,
            PADOUT => \N__7331\,
            PADIN => \N__7330\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2488\,
            DIN0 => \D_UU_AMIGA_in_2\,
            DOUT0 => \N__2735\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7323\,
            DIN => \N__7322\,
            DOUT => \N__7321\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7323\,
            PADOUT => \N__7322\,
            PADIN => \N__7321\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7314\,
            DIN => \N__7313\,
            DOUT => \N__7312\,
            PACKAGEPIN => D_LM_AMIGA(6)
        );

    \D_LM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7314\,
            PADOUT => \N__7313\,
            PADIN => \N__7312\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2500\,
            DIN0 => \D_LM_AMIGA_in_6\,
            DOUT0 => \N__5378\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7305\,
            DIN => \N__7304\,
            DOUT => \N__7303\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7305\,
            PADOUT => \N__7304\,
            PADIN => \N__7303\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7296\,
            DIN => \N__7295\,
            DOUT => \N__7294\,
            PACKAGEPIN => D_LM_040(5)
        );

    \D_LM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7296\,
            PADOUT => \N__7295\,
            PADIN => \N__7294\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4445\,
            DIN0 => \D_LM_040_in_5\,
            DOUT0 => \N__3083\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7287\,
            DIN => \N__7286\,
            DOUT => \N__7285\,
            PACKAGEPIN => D_UM_040(6)
        );

    \D_UM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7287\,
            PADOUT => \N__7286\,
            PADIN => \N__7285\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4406\,
            DIN0 => \D_UM_040_in_6\,
            DOUT0 => \N__6746\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TAn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7278\,
            DIN => \N__7277\,
            DOUT => \N__7276\,
            PACKAGEPIN => \TAn_wire\
        );

    \TAn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7278\,
            PADOUT => \N__7277\,
            PADIN => \N__7276\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3398\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMAn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7269\,
            DIN => \N__7268\,
            DOUT => \N__7267\,
            PACKAGEPIN => \DMAn_wire\
        );

    \DMAn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7269\,
            PADOUT => \N__7268\,
            PADIN => \N__7267\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5042\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7260\,
            DIN => \N__7259\,
            DOUT => \N__7258\,
            PACKAGEPIN => D_LL_040(6)
        );

    \D_LL_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7260\,
            PADOUT => \N__7259\,
            PADIN => \N__7258\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4594\,
            DIN0 => \D_LL_040_in_6\,
            DOUT0 => \N__4964\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7251\,
            DIN => \N__7250\,
            DOUT => \N__7249\,
            PACKAGEPIN => D_LL_AMIGA(5)
        );

    \D_LL_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7251\,
            PADOUT => \N__7250\,
            PADIN => \N__7249\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2424\,
            DIN0 => \D_LL_AMIGA_in_5\,
            DOUT0 => \N__4124\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7242\,
            DIN => \N__7241\,
            DOUT => \N__7240\,
            PACKAGEPIN => D_UM_AMIGA(0)
        );

    \D_UM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7242\,
            PADOUT => \N__7241\,
            PADIN => \N__7240\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2399\,
            DIN0 => \D_UM_AMIGA_in_0\,
            DOUT0 => \N__3863\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7233\,
            DIN => \N__7232\,
            DOUT => \N__7231\,
            PACKAGEPIN => D_UU_040(2)
        );

    \D_UU_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7233\,
            PADOUT => \N__7232\,
            PADIN => \N__7231\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4587\,
            DIN0 => \D_UU_040_in_2\,
            DOUT0 => \N__5567\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7224\,
            DIN => \N__7223\,
            DOUT => \N__7222\,
            PACKAGEPIN => D_LM_AMIGA(2)
        );

    \D_LM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7224\,
            PADOUT => \N__7223\,
            PADIN => \N__7222\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2398\,
            DIN0 => \D_LM_AMIGA_in_2\,
            DOUT0 => \N__2795\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK80_CPU_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7215\,
            DIN => \N__7214\,
            DOUT => \N__7213\,
            PACKAGEPIN => \CLK80_CPU_wire\
        );

    \CLK80_CPU_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7215\,
            PADOUT => \N__7214\,
            PADIN => \N__7213\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4878\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7206\,
            DIN => \N__7205\,
            DOUT => \N__7204\,
            PACKAGEPIN => D_LL_040(3)
        );

    \D_LL_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7206\,
            PADOUT => \N__7205\,
            PADIN => \N__7204\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4629\,
            DIN0 => \D_LL_040_in_3\,
            DOUT0 => \N__2243\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7197\,
            DIN => \N__7196\,
            DOUT => \N__7195\,
            PACKAGEPIN => D_LM_040(1)
        );

    \D_LM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7197\,
            PADOUT => \N__7196\,
            PADIN => \N__7195\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4589\,
            DIN0 => \D_LM_040_in_1\,
            DOUT0 => \N__3224\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7188\,
            DIN => \N__7187\,
            DOUT => \N__7186\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7188\,
            PADOUT => \N__7187\,
            PADIN => \N__7186\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3680\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7179\,
            DIN => \N__7178\,
            DOUT => \N__7177\,
            PACKAGEPIN => D_UM_AMIGA(7)
        );

    \D_UM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7179\,
            PADOUT => \N__7178\,
            PADIN => \N__7177\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2522\,
            DIN0 => \D_UM_AMIGA_in_7\,
            DOUT0 => \N__6233\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7170\,
            DIN => \N__7169\,
            DOUT => \N__7168\,
            PACKAGEPIN => D_LM_AMIGA(7)
        );

    \D_LM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7170\,
            PADOUT => \N__7169\,
            PADIN => \N__7168\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2499\,
            DIN0 => \D_LM_AMIGA_in_7\,
            DOUT0 => \N__3350\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7161\,
            DIN => \N__7160\,
            DOUT => \N__7159\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7161\,
            PADOUT => \N__7160\,
            PADIN => \N__7159\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \PORTSIZE_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7152\,
            DIN => \N__7151\,
            DOUT => \N__7150\,
            PACKAGEPIN => \A_AMIGA_wire\(0)
        );

    \A_AMIGA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7152\,
            PADOUT => \N__7151\,
            PADIN => \N__7150\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2552\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7143\,
            DIN => \N__7142\,
            DOUT => \N__7141\,
            PACKAGEPIN => D_LM_040(4)
        );

    \D_LM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7143\,
            PADOUT => \N__7142\,
            PADIN => \N__7141\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4519\,
            DIN0 => \D_LM_040_in_4\,
            DOUT0 => \N__3722\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7134\,
            DIN => \N__7133\,
            DOUT => \N__7132\,
            PACKAGEPIN => D_UM_040(7)
        );

    \D_UM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7134\,
            PADOUT => \N__7133\,
            PADIN => \N__7132\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4493\,
            DIN0 => \D_UM_040_in_7\,
            DOUT0 => \N__5639\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7125\,
            DIN => \N__7124\,
            DOUT => \N__7123\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7125\,
            PADOUT => \N__7124\,
            PADIN => \N__7123\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7116\,
            DIN => \N__7115\,
            DOUT => \N__7114\,
            PACKAGEPIN => D_UU_AMIGA(1)
        );

    \D_UU_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7116\,
            PADOUT => \N__7115\,
            PADIN => \N__7114\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2501\,
            DIN0 => \D_UU_AMIGA_in_1\,
            DOUT0 => \N__6329\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7107\,
            DIN => \N__7106\,
            DOUT => \N__7105\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7107\,
            PADOUT => \N__7106\,
            PADIN => \N__7105\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3840\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7098\,
            DIN => \N__7097\,
            DOUT => \N__7096\,
            PACKAGEPIN => D_UM_040(0)
        );

    \D_UM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7098\,
            PADOUT => \N__7097\,
            PADIN => \N__7096\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4444\,
            DIN0 => \D_UM_040_in_0\,
            DOUT0 => \N__3806\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7089\,
            DIN => \N__7088\,
            DOUT => \N__7087\,
            PACKAGEPIN => D_LL_AMIGA(0)
        );

    \D_LL_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7089\,
            PADOUT => \N__7088\,
            PADIN => \N__7087\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2332\,
            DIN0 => \D_LL_AMIGA_in_0\,
            DOUT0 => \N__3920\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7080\,
            DIN => \N__7079\,
            DOUT => \N__7078\,
            PACKAGEPIN => D_UU_AMIGA(4)
        );

    \D_UU_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7080\,
            PADOUT => \N__7079\,
            PADIN => \N__7078\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2487\,
            DIN0 => \D_UU_AMIGA_in_4\,
            DOUT0 => \N__5882\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7071\,
            DIN => \N__7070\,
            DOUT => \N__7069\,
            PACKAGEPIN => D_UU_040(7)
        );

    \D_UU_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7071\,
            PADOUT => \N__7070\,
            PADIN => \N__7069\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4549\,
            DIN0 => \D_UU_040_in_7\,
            DOUT0 => \N__6803\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7062\,
            DIN => \N__7061\,
            DOUT => \N__7060\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7062\,
            PADOUT => \N__7061\,
            PADIN => \N__7060\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7053\,
            DIN => \N__7052\,
            DOUT => \N__7051\,
            PACKAGEPIN => D_LL_040(0)
        );

    \D_LL_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7053\,
            PADOUT => \N__7052\,
            PADIN => \N__7051\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4630\,
            DIN0 => \D_LL_040_in_0\,
            DOUT0 => \N__2699\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7044\,
            DIN => \N__7043\,
            DOUT => \N__7042\,
            PACKAGEPIN => D_UM_AMIGA(2)
        );

    \D_UM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7044\,
            PADOUT => \N__7043\,
            PADIN => \N__7042\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2451\,
            DIN0 => \D_UM_AMIGA_in_2\,
            DOUT0 => \N__2585\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7035\,
            DIN => \N__7034\,
            DOUT => \N__7033\,
            PACKAGEPIN => D_UU_040(0)
        );

    \D_UU_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7035\,
            PADOUT => \N__7034\,
            PADIN => \N__7033\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4482\,
            DIN0 => \D_UU_040_in_0\,
            DOUT0 => \N__5057\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1799\ : InMux
    port map (
            O => \N__7016\,
            I => \N__7013\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__7013\,
            I => \N__7010\
        );

    \I__1797\ : Span4Mux_v
    port map (
            O => \N__7010\,
            I => \N__7007\
        );

    \I__1796\ : Span4Mux_v
    port map (
            O => \N__7007\,
            I => \N__7004\
        );

    \I__1795\ : Sp12to4
    port map (
            O => \N__7004\,
            I => \N__7001\
        );

    \I__1794\ : Span12Mux_h
    port map (
            O => \N__7001\,
            I => \N__6998\
        );

    \I__1793\ : Odrv12
    port map (
            O => \N__6998\,
            I => \SIZ_c_1\
        );

    \I__1792\ : InMux
    port map (
            O => \N__6995\,
            I => \N__6992\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__6992\,
            I => \N__6989\
        );

    \I__1790\ : Span4Mux_v
    port map (
            O => \N__6989\,
            I => \N__6986\
        );

    \I__1789\ : Span4Mux_h
    port map (
            O => \N__6986\,
            I => \N__6983\
        );

    \I__1788\ : Sp12to4
    port map (
            O => \N__6983\,
            I => \N__6980\
        );

    \I__1787\ : Odrv12
    port map (
            O => \N__6980\,
            I => \SIZ_c_0\
        );

    \I__1786\ : InMux
    port map (
            O => \N__6977\,
            I => \N__6974\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__6974\,
            I => \N__6970\
        );

    \I__1784\ : InMux
    port map (
            O => \N__6973\,
            I => \N__6967\
        );

    \I__1783\ : Span4Mux_v
    port map (
            O => \N__6970\,
            I => \N__6964\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__6967\,
            I => \N__6961\
        );

    \I__1781\ : Sp12to4
    port map (
            O => \N__6964\,
            I => \N__6958\
        );

    \I__1780\ : Span12Mux_v
    port map (
            O => \N__6961\,
            I => \N__6955\
        );

    \I__1779\ : Span12Mux_h
    port map (
            O => \N__6958\,
            I => \N__6952\
        );

    \I__1778\ : Span12Mux_h
    port map (
            O => \N__6955\,
            I => \N__6949\
        );

    \I__1777\ : Span12Mux_v
    port map (
            O => \N__6952\,
            I => \N__6946\
        );

    \I__1776\ : Odrv12
    port map (
            O => \N__6949\,
            I => \PORTSIZE_c\
        );

    \I__1775\ : Odrv12
    port map (
            O => \N__6946\,
            I => \PORTSIZE_c\
        );

    \I__1774\ : InMux
    port map (
            O => \N__6941\,
            I => \N__6937\
        );

    \I__1773\ : InMux
    port map (
            O => \N__6940\,
            I => \N__6934\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__6937\,
            I => \N__6931\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__6934\,
            I => \N__6928\
        );

    \I__1770\ : Span4Mux_v
    port map (
            O => \N__6931\,
            I => \N__6925\
        );

    \I__1769\ : Span12Mux_v
    port map (
            O => \N__6928\,
            I => \N__6922\
        );

    \I__1768\ : Span4Mux_h
    port map (
            O => \N__6925\,
            I => \N__6919\
        );

    \I__1767\ : Odrv12
    port map (
            O => \N__6922\,
            I => \U111_CYCLE_SM.LW_TRANS_0\
        );

    \I__1766\ : Odrv4
    port map (
            O => \N__6919\,
            I => \U111_CYCLE_SM.LW_TRANS_0\
        );

    \I__1765\ : InMux
    port map (
            O => \N__6914\,
            I => \N__6911\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__6911\,
            I => \N__6907\
        );

    \I__1763\ : InMux
    port map (
            O => \N__6910\,
            I => \N__6903\
        );

    \I__1762\ : Span4Mux_v
    port map (
            O => \N__6907\,
            I => \N__6900\
        );

    \I__1761\ : InMux
    port map (
            O => \N__6906\,
            I => \N__6897\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__6903\,
            I => \N__6894\
        );

    \I__1759\ : Sp12to4
    port map (
            O => \N__6900\,
            I => \N__6891\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__6897\,
            I => \N__6888\
        );

    \I__1757\ : Span12Mux_v
    port map (
            O => \N__6894\,
            I => \N__6885\
        );

    \I__1756\ : Span12Mux_h
    port map (
            O => \N__6891\,
            I => \N__6882\
        );

    \I__1755\ : Span12Mux_s7_v
    port map (
            O => \N__6888\,
            I => \N__6879\
        );

    \I__1754\ : Span12Mux_h
    port map (
            O => \N__6885\,
            I => \N__6876\
        );

    \I__1753\ : Span12Mux_v
    port map (
            O => \N__6882\,
            I => \N__6871\
        );

    \I__1752\ : Span12Mux_h
    port map (
            O => \N__6879\,
            I => \N__6871\
        );

    \I__1751\ : Odrv12
    port map (
            O => \N__6876\,
            I => \D_UM_AMIGA_in_5\
        );

    \I__1750\ : Odrv12
    port map (
            O => \N__6871\,
            I => \D_UM_AMIGA_in_5\
        );

    \I__1749\ : IoInMux
    port map (
            O => \N__6866\,
            I => \N__6863\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__6863\,
            I => \N__6860\
        );

    \I__1747\ : Span4Mux_s0_v
    port map (
            O => \N__6860\,
            I => \N__6857\
        );

    \I__1746\ : Sp12to4
    port map (
            O => \N__6857\,
            I => \N__6854\
        );

    \I__1745\ : Span12Mux_h
    port map (
            O => \N__6854\,
            I => \N__6851\
        );

    \I__1744\ : Odrv12
    port map (
            O => \N__6851\,
            I => \un1_D_UM_AMIGA_5\
        );

    \I__1743\ : InMux
    port map (
            O => \N__6848\,
            I => \N__6845\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__6845\,
            I => \N__6842\
        );

    \I__1741\ : Odrv12
    port map (
            O => \N__6842\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\
        );

    \I__1740\ : InMux
    port map (
            O => \N__6839\,
            I => \N__6836\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__6836\,
            I => \N__6832\
        );

    \I__1738\ : InMux
    port map (
            O => \N__6835\,
            I => \N__6829\
        );

    \I__1737\ : Span4Mux_v
    port map (
            O => \N__6832\,
            I => \N__6823\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__6829\,
            I => \N__6823\
        );

    \I__1735\ : InMux
    port map (
            O => \N__6828\,
            I => \N__6820\
        );

    \I__1734\ : Span4Mux_v
    port map (
            O => \N__6823\,
            I => \N__6815\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__6820\,
            I => \N__6815\
        );

    \I__1732\ : Span4Mux_v
    port map (
            O => \N__6815\,
            I => \N__6812\
        );

    \I__1731\ : Sp12to4
    port map (
            O => \N__6812\,
            I => \N__6809\
        );

    \I__1730\ : Span12Mux_h
    port map (
            O => \N__6809\,
            I => \N__6806\
        );

    \I__1729\ : Odrv12
    port map (
            O => \N__6806\,
            I => \D_UU_AMIGA_in_7\
        );

    \I__1728\ : IoInMux
    port map (
            O => \N__6803\,
            I => \N__6800\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__6800\,
            I => \N__6797\
        );

    \I__1726\ : Span12Mux_s11_v
    port map (
            O => \N__6797\,
            I => \N__6794\
        );

    \I__1725\ : Span12Mux_h
    port map (
            O => \N__6794\,
            I => \N__6791\
        );

    \I__1724\ : Odrv12
    port map (
            O => \N__6791\,
            I => \un1_D_UU_AMIGA_7\
        );

    \I__1723\ : InMux
    port map (
            O => \N__6788\,
            I => \N__6785\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__6785\,
            I => \N__6782\
        );

    \I__1721\ : Span4Mux_v
    port map (
            O => \N__6782\,
            I => \N__6779\
        );

    \I__1720\ : Span4Mux_v
    port map (
            O => \N__6779\,
            I => \N__6774\
        );

    \I__1719\ : InMux
    port map (
            O => \N__6778\,
            I => \N__6771\
        );

    \I__1718\ : InMux
    port map (
            O => \N__6777\,
            I => \N__6768\
        );

    \I__1717\ : Sp12to4
    port map (
            O => \N__6774\,
            I => \N__6761\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__6771\,
            I => \N__6761\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__6768\,
            I => \N__6761\
        );

    \I__1714\ : Span12Mux_h
    port map (
            O => \N__6761\,
            I => \N__6758\
        );

    \I__1713\ : Span12Mux_v
    port map (
            O => \N__6758\,
            I => \N__6755\
        );

    \I__1712\ : Odrv12
    port map (
            O => \N__6755\,
            I => \D_UM_AMIGA_in_6\
        );

    \I__1711\ : InMux
    port map (
            O => \N__6752\,
            I => \N__6749\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__6749\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\
        );

    \I__1709\ : IoInMux
    port map (
            O => \N__6746\,
            I => \N__6743\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__6743\,
            I => \N__6740\
        );

    \I__1707\ : IoSpan4Mux
    port map (
            O => \N__6740\,
            I => \N__6737\
        );

    \I__1706\ : Span4Mux_s3_h
    port map (
            O => \N__6737\,
            I => \N__6734\
        );

    \I__1705\ : Span4Mux_h
    port map (
            O => \N__6734\,
            I => \N__6731\
        );

    \I__1704\ : Span4Mux_h
    port map (
            O => \N__6731\,
            I => \N__6728\
        );

    \I__1703\ : Odrv4
    port map (
            O => \N__6728\,
            I => \un1_D_UM_AMIGA_6\
        );

    \I__1702\ : IoInMux
    port map (
            O => \N__6725\,
            I => \N__6721\
        );

    \I__1701\ : InMux
    port map (
            O => \N__6724\,
            I => \N__6718\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__6721\,
            I => \N__6715\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__6718\,
            I => \N__6712\
        );

    \I__1698\ : Span4Mux_s3_h
    port map (
            O => \N__6715\,
            I => \N__6709\
        );

    \I__1697\ : Span4Mux_v
    port map (
            O => \N__6712\,
            I => \N__6706\
        );

    \I__1696\ : Sp12to4
    port map (
            O => \N__6709\,
            I => \N__6703\
        );

    \I__1695\ : Span4Mux_v
    port map (
            O => \N__6706\,
            I => \N__6700\
        );

    \I__1694\ : Span12Mux_v
    port map (
            O => \N__6703\,
            I => \N__6697\
        );

    \I__1693\ : Sp12to4
    port map (
            O => \N__6700\,
            I => \N__6694\
        );

    \I__1692\ : Span12Mux_h
    port map (
            O => \N__6697\,
            I => \N__6691\
        );

    \I__1691\ : Span12Mux_h
    port map (
            O => \N__6694\,
            I => \N__6688\
        );

    \I__1690\ : Span12Mux_h
    port map (
            O => \N__6691\,
            I => \N__6685\
        );

    \I__1689\ : Span12Mux_v
    port map (
            O => \N__6688\,
            I => \N__6682\
        );

    \I__1688\ : Odrv12
    port map (
            O => \N__6685\,
            I => \D_LL_040_in_1\
        );

    \I__1687\ : Odrv12
    port map (
            O => \N__6682\,
            I => \D_LL_040_in_1\
        );

    \I__1686\ : InMux
    port map (
            O => \N__6677\,
            I => \N__6674\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__6674\,
            I => \N__6671\
        );

    \I__1684\ : Span12Mux_v
    port map (
            O => \N__6671\,
            I => \N__6668\
        );

    \I__1683\ : Span12Mux_h
    port map (
            O => \N__6668\,
            I => \N__6665\
        );

    \I__1682\ : Odrv12
    port map (
            O => \N__6665\,
            I => \D_UM_040_in_1\
        );

    \I__1681\ : IoInMux
    port map (
            O => \N__6662\,
            I => \N__6659\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__6659\,
            I => \N__6656\
        );

    \I__1679\ : IoSpan4Mux
    port map (
            O => \N__6656\,
            I => \N__6653\
        );

    \I__1678\ : Span4Mux_s3_h
    port map (
            O => \N__6653\,
            I => \N__6650\
        );

    \I__1677\ : Span4Mux_h
    port map (
            O => \N__6650\,
            I => \N__6647\
        );

    \I__1676\ : Span4Mux_h
    port map (
            O => \N__6647\,
            I => \N__6644\
        );

    \I__1675\ : Span4Mux_h
    port map (
            O => \N__6644\,
            I => \N__6641\
        );

    \I__1674\ : Odrv4
    port map (
            O => \N__6641\,
            I => \un1_D_UM_040_1\
        );

    \I__1673\ : InMux
    port map (
            O => \N__6638\,
            I => \N__6633\
        );

    \I__1672\ : InMux
    port map (
            O => \N__6637\,
            I => \N__6621\
        );

    \I__1671\ : InMux
    port map (
            O => \N__6636\,
            I => \N__6621\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__6633\,
            I => \N__6617\
        );

    \I__1669\ : InMux
    port map (
            O => \N__6632\,
            I => \N__6606\
        );

    \I__1668\ : InMux
    port map (
            O => \N__6631\,
            I => \N__6606\
        );

    \I__1667\ : InMux
    port map (
            O => \N__6630\,
            I => \N__6606\
        );

    \I__1666\ : InMux
    port map (
            O => \N__6629\,
            I => \N__6603\
        );

    \I__1665\ : InMux
    port map (
            O => \N__6628\,
            I => \N__6598\
        );

    \I__1664\ : InMux
    port map (
            O => \N__6627\,
            I => \N__6598\
        );

    \I__1663\ : InMux
    port map (
            O => \N__6626\,
            I => \N__6595\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__6621\,
            I => \N__6589\
        );

    \I__1661\ : InMux
    port map (
            O => \N__6620\,
            I => \N__6586\
        );

    \I__1660\ : Span4Mux_h
    port map (
            O => \N__6617\,
            I => \N__6583\
        );

    \I__1659\ : InMux
    port map (
            O => \N__6616\,
            I => \N__6578\
        );

    \I__1658\ : InMux
    port map (
            O => \N__6615\,
            I => \N__6578\
        );

    \I__1657\ : InMux
    port map (
            O => \N__6614\,
            I => \N__6575\
        );

    \I__1656\ : InMux
    port map (
            O => \N__6613\,
            I => \N__6572\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__6606\,
            I => \N__6563\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__6603\,
            I => \N__6563\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__6598\,
            I => \N__6563\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__6595\,
            I => \N__6563\
        );

    \I__1651\ : InMux
    port map (
            O => \N__6594\,
            I => \N__6560\
        );

    \I__1650\ : InMux
    port map (
            O => \N__6593\,
            I => \N__6557\
        );

    \I__1649\ : InMux
    port map (
            O => \N__6592\,
            I => \N__6554\
        );

    \I__1648\ : Span12Mux_h
    port map (
            O => \N__6589\,
            I => \N__6550\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__6586\,
            I => \N__6547\
        );

    \I__1646\ : Span4Mux_v
    port map (
            O => \N__6583\,
            I => \N__6544\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__6578\,
            I => \N__6541\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__6575\,
            I => \N__6538\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__6572\,
            I => \N__6535\
        );

    \I__1642\ : Span4Mux_v
    port map (
            O => \N__6563\,
            I => \N__6526\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__6560\,
            I => \N__6526\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__6557\,
            I => \N__6526\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__6554\,
            I => \N__6526\
        );

    \I__1638\ : InMux
    port map (
            O => \N__6553\,
            I => \N__6523\
        );

    \I__1637\ : Span12Mux_v
    port map (
            O => \N__6550\,
            I => \N__6518\
        );

    \I__1636\ : Span12Mux_h
    port map (
            O => \N__6547\,
            I => \N__6515\
        );

    \I__1635\ : Span4Mux_v
    port map (
            O => \N__6544\,
            I => \N__6508\
        );

    \I__1634\ : Span4Mux_v
    port map (
            O => \N__6541\,
            I => \N__6508\
        );

    \I__1633\ : Span4Mux_h
    port map (
            O => \N__6538\,
            I => \N__6508\
        );

    \I__1632\ : Span4Mux_v
    port map (
            O => \N__6535\,
            I => \N__6503\
        );

    \I__1631\ : Span4Mux_v
    port map (
            O => \N__6526\,
            I => \N__6503\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__6523\,
            I => \N__6500\
        );

    \I__1629\ : InMux
    port map (
            O => \N__6522\,
            I => \N__6497\
        );

    \I__1628\ : InMux
    port map (
            O => \N__6521\,
            I => \N__6494\
        );

    \I__1627\ : Odrv12
    port map (
            O => \N__6518\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1626\ : Odrv12
    port map (
            O => \N__6515\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1625\ : Odrv4
    port map (
            O => \N__6508\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1624\ : Odrv4
    port map (
            O => \N__6503\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1623\ : Odrv4
    port map (
            O => \N__6500\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__6497\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__6494\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1620\ : InMux
    port map (
            O => \N__6479\,
            I => \N__6476\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__6476\,
            I => \N__6473\
        );

    \I__1618\ : Span4Mux_v
    port map (
            O => \N__6473\,
            I => \N__6470\
        );

    \I__1617\ : Odrv4
    port map (
            O => \N__6470\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\
        );

    \I__1616\ : InMux
    port map (
            O => \N__6467\,
            I => \N__6463\
        );

    \I__1615\ : InMux
    port map (
            O => \N__6466\,
            I => \N__6460\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__6463\,
            I => \N__6456\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__6460\,
            I => \N__6453\
        );

    \I__1612\ : InMux
    port map (
            O => \N__6459\,
            I => \N__6450\
        );

    \I__1611\ : Span4Mux_v
    port map (
            O => \N__6456\,
            I => \N__6447\
        );

    \I__1610\ : Span4Mux_v
    port map (
            O => \N__6453\,
            I => \N__6444\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__6450\,
            I => \N__6441\
        );

    \I__1608\ : Span4Mux_h
    port map (
            O => \N__6447\,
            I => \N__6436\
        );

    \I__1607\ : Span4Mux_v
    port map (
            O => \N__6444\,
            I => \N__6436\
        );

    \I__1606\ : Span4Mux_v
    port map (
            O => \N__6441\,
            I => \N__6433\
        );

    \I__1605\ : Span4Mux_v
    port map (
            O => \N__6436\,
            I => \N__6430\
        );

    \I__1604\ : Sp12to4
    port map (
            O => \N__6433\,
            I => \N__6427\
        );

    \I__1603\ : Sp12to4
    port map (
            O => \N__6430\,
            I => \N__6422\
        );

    \I__1602\ : Span12Mux_h
    port map (
            O => \N__6427\,
            I => \N__6422\
        );

    \I__1601\ : Odrv12
    port map (
            O => \N__6422\,
            I => \D_UU_AMIGA_in_1\
        );

    \I__1600\ : IoInMux
    port map (
            O => \N__6419\,
            I => \N__6416\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__6416\,
            I => \N__6413\
        );

    \I__1598\ : IoSpan4Mux
    port map (
            O => \N__6413\,
            I => \N__6410\
        );

    \I__1597\ : Span4Mux_s3_h
    port map (
            O => \N__6410\,
            I => \N__6407\
        );

    \I__1596\ : Sp12to4
    port map (
            O => \N__6407\,
            I => \N__6404\
        );

    \I__1595\ : Span12Mux_h
    port map (
            O => \N__6404\,
            I => \N__6401\
        );

    \I__1594\ : Odrv12
    port map (
            O => \N__6401\,
            I => \un1_D_UU_AMIGA_1\
        );

    \I__1593\ : IoInMux
    port map (
            O => \N__6398\,
            I => \N__6394\
        );

    \I__1592\ : InMux
    port map (
            O => \N__6397\,
            I => \N__6391\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__6394\,
            I => \N__6388\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__6391\,
            I => \N__6385\
        );

    \I__1589\ : Span4Mux_s3_h
    port map (
            O => \N__6388\,
            I => \N__6382\
        );

    \I__1588\ : Span4Mux_h
    port map (
            O => \N__6385\,
            I => \N__6379\
        );

    \I__1587\ : Sp12to4
    port map (
            O => \N__6382\,
            I => \N__6376\
        );

    \I__1586\ : Sp12to4
    port map (
            O => \N__6379\,
            I => \N__6373\
        );

    \I__1585\ : Span12Mux_v
    port map (
            O => \N__6376\,
            I => \N__6370\
        );

    \I__1584\ : Span12Mux_v
    port map (
            O => \N__6373\,
            I => \N__6367\
        );

    \I__1583\ : Span12Mux_h
    port map (
            O => \N__6370\,
            I => \N__6364\
        );

    \I__1582\ : Span12Mux_v
    port map (
            O => \N__6367\,
            I => \N__6361\
        );

    \I__1581\ : Span12Mux_h
    port map (
            O => \N__6364\,
            I => \N__6358\
        );

    \I__1580\ : Span12Mux_h
    port map (
            O => \N__6361\,
            I => \N__6355\
        );

    \I__1579\ : Odrv12
    port map (
            O => \N__6358\,
            I => \D_LM_040_in_1\
        );

    \I__1578\ : Odrv12
    port map (
            O => \N__6355\,
            I => \D_LM_040_in_1\
        );

    \I__1577\ : InMux
    port map (
            O => \N__6350\,
            I => \N__6347\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__6347\,
            I => \N__6344\
        );

    \I__1575\ : Span4Mux_v
    port map (
            O => \N__6344\,
            I => \N__6341\
        );

    \I__1574\ : Span4Mux_v
    port map (
            O => \N__6341\,
            I => \N__6338\
        );

    \I__1573\ : Sp12to4
    port map (
            O => \N__6338\,
            I => \N__6335\
        );

    \I__1572\ : Span12Mux_h
    port map (
            O => \N__6335\,
            I => \N__6332\
        );

    \I__1571\ : Odrv12
    port map (
            O => \N__6332\,
            I => \D_UU_040_in_1\
        );

    \I__1570\ : IoInMux
    port map (
            O => \N__6329\,
            I => \N__6326\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__6326\,
            I => \N__6323\
        );

    \I__1568\ : IoSpan4Mux
    port map (
            O => \N__6323\,
            I => \N__6320\
        );

    \I__1567\ : Span4Mux_s3_h
    port map (
            O => \N__6320\,
            I => \N__6317\
        );

    \I__1566\ : Span4Mux_h
    port map (
            O => \N__6317\,
            I => \N__6314\
        );

    \I__1565\ : Span4Mux_h
    port map (
            O => \N__6314\,
            I => \N__6311\
        );

    \I__1564\ : Span4Mux_h
    port map (
            O => \N__6311\,
            I => \N__6308\
        );

    \I__1563\ : Odrv4
    port map (
            O => \N__6308\,
            I => \un1_D_UU_040_1\
        );

    \I__1562\ : IoInMux
    port map (
            O => \N__6305\,
            I => \N__6302\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__6302\,
            I => \N__6298\
        );

    \I__1560\ : InMux
    port map (
            O => \N__6301\,
            I => \N__6295\
        );

    \I__1559\ : IoSpan4Mux
    port map (
            O => \N__6298\,
            I => \N__6292\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__6295\,
            I => \N__6289\
        );

    \I__1557\ : Span4Mux_s3_h
    port map (
            O => \N__6292\,
            I => \N__6286\
        );

    \I__1556\ : Span4Mux_h
    port map (
            O => \N__6289\,
            I => \N__6283\
        );

    \I__1555\ : Sp12to4
    port map (
            O => \N__6286\,
            I => \N__6280\
        );

    \I__1554\ : Sp12to4
    port map (
            O => \N__6283\,
            I => \N__6277\
        );

    \I__1553\ : Span12Mux_v
    port map (
            O => \N__6280\,
            I => \N__6274\
        );

    \I__1552\ : Span12Mux_v
    port map (
            O => \N__6277\,
            I => \N__6271\
        );

    \I__1551\ : Span12Mux_h
    port map (
            O => \N__6274\,
            I => \N__6268\
        );

    \I__1550\ : Span12Mux_v
    port map (
            O => \N__6271\,
            I => \N__6265\
        );

    \I__1549\ : Span12Mux_h
    port map (
            O => \N__6268\,
            I => \N__6262\
        );

    \I__1548\ : Span12Mux_h
    port map (
            O => \N__6265\,
            I => \N__6259\
        );

    \I__1547\ : Odrv12
    port map (
            O => \N__6262\,
            I => \D_LL_040_in_7\
        );

    \I__1546\ : Odrv12
    port map (
            O => \N__6259\,
            I => \D_LL_040_in_7\
        );

    \I__1545\ : InMux
    port map (
            O => \N__6254\,
            I => \N__6251\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__6251\,
            I => \N__6248\
        );

    \I__1543\ : Span4Mux_v
    port map (
            O => \N__6248\,
            I => \N__6245\
        );

    \I__1542\ : Span4Mux_v
    port map (
            O => \N__6245\,
            I => \N__6242\
        );

    \I__1541\ : Sp12to4
    port map (
            O => \N__6242\,
            I => \N__6239\
        );

    \I__1540\ : Span12Mux_h
    port map (
            O => \N__6239\,
            I => \N__6236\
        );

    \I__1539\ : Odrv12
    port map (
            O => \N__6236\,
            I => \D_UM_040_in_7\
        );

    \I__1538\ : IoInMux
    port map (
            O => \N__6233\,
            I => \N__6230\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__6230\,
            I => \N__6227\
        );

    \I__1536\ : Span12Mux_s5_h
    port map (
            O => \N__6227\,
            I => \N__6224\
        );

    \I__1535\ : Span12Mux_h
    port map (
            O => \N__6224\,
            I => \N__6221\
        );

    \I__1534\ : Odrv12
    port map (
            O => \N__6221\,
            I => \un1_D_UM_040_7\
        );

    \I__1533\ : IoInMux
    port map (
            O => \N__6218\,
            I => \N__6215\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__6215\,
            I => \N__6212\
        );

    \I__1531\ : Span4Mux_s1_h
    port map (
            O => \N__6212\,
            I => \N__6209\
        );

    \I__1530\ : Sp12to4
    port map (
            O => \N__6209\,
            I => \N__6205\
        );

    \I__1529\ : InMux
    port map (
            O => \N__6208\,
            I => \N__6202\
        );

    \I__1528\ : Span12Mux_v
    port map (
            O => \N__6205\,
            I => \N__6199\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__6202\,
            I => \N__6196\
        );

    \I__1526\ : Span12Mux_h
    port map (
            O => \N__6199\,
            I => \N__6193\
        );

    \I__1525\ : Span12Mux_v
    port map (
            O => \N__6196\,
            I => \N__6190\
        );

    \I__1524\ : Span12Mux_h
    port map (
            O => \N__6193\,
            I => \N__6187\
        );

    \I__1523\ : Span12Mux_h
    port map (
            O => \N__6190\,
            I => \N__6184\
        );

    \I__1522\ : Odrv12
    port map (
            O => \N__6187\,
            I => \D_LM_040_in_4\
        );

    \I__1521\ : Odrv12
    port map (
            O => \N__6184\,
            I => \D_LM_040_in_4\
        );

    \I__1520\ : InMux
    port map (
            O => \N__6179\,
            I => \N__6176\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__6176\,
            I => \N__6173\
        );

    \I__1518\ : Span4Mux_h
    port map (
            O => \N__6173\,
            I => \N__6170\
        );

    \I__1517\ : Span4Mux_v
    port map (
            O => \N__6170\,
            I => \N__6167\
        );

    \I__1516\ : Span4Mux_h
    port map (
            O => \N__6167\,
            I => \N__6164\
        );

    \I__1515\ : Odrv4
    port map (
            O => \N__6164\,
            I => \D_UU_040_in_4\
        );

    \I__1514\ : InMux
    port map (
            O => \N__6161\,
            I => \N__6153\
        );

    \I__1513\ : InMux
    port map (
            O => \N__6160\,
            I => \N__6150\
        );

    \I__1512\ : InMux
    port map (
            O => \N__6159\,
            I => \N__6147\
        );

    \I__1511\ : InMux
    port map (
            O => \N__6158\,
            I => \N__6144\
        );

    \I__1510\ : InMux
    port map (
            O => \N__6157\,
            I => \N__6140\
        );

    \I__1509\ : InMux
    port map (
            O => \N__6156\,
            I => \N__6135\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__6153\,
            I => \N__6125\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__6150\,
            I => \N__6125\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__6147\,
            I => \N__6125\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__6144\,
            I => \N__6125\
        );

    \I__1504\ : InMux
    port map (
            O => \N__6143\,
            I => \N__6122\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__6140\,
            I => \N__6118\
        );

    \I__1502\ : InMux
    port map (
            O => \N__6139\,
            I => \N__6115\
        );

    \I__1501\ : InMux
    port map (
            O => \N__6138\,
            I => \N__6112\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__6135\,
            I => \N__6107\
        );

    \I__1499\ : InMux
    port map (
            O => \N__6134\,
            I => \N__6104\
        );

    \I__1498\ : Span4Mux_v
    port map (
            O => \N__6125\,
            I => \N__6099\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__6122\,
            I => \N__6099\
        );

    \I__1496\ : InMux
    port map (
            O => \N__6121\,
            I => \N__6093\
        );

    \I__1495\ : Span4Mux_h
    port map (
            O => \N__6118\,
            I => \N__6085\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__6115\,
            I => \N__6085\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__6112\,
            I => \N__6085\
        );

    \I__1492\ : InMux
    port map (
            O => \N__6111\,
            I => \N__6082\
        );

    \I__1491\ : InMux
    port map (
            O => \N__6110\,
            I => \N__6073\
        );

    \I__1490\ : Span4Mux_h
    port map (
            O => \N__6107\,
            I => \N__6068\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__6104\,
            I => \N__6068\
        );

    \I__1488\ : Span4Mux_v
    port map (
            O => \N__6099\,
            I => \N__6064\
        );

    \I__1487\ : InMux
    port map (
            O => \N__6098\,
            I => \N__6061\
        );

    \I__1486\ : InMux
    port map (
            O => \N__6097\,
            I => \N__6058\
        );

    \I__1485\ : InMux
    port map (
            O => \N__6096\,
            I => \N__6055\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__6093\,
            I => \N__6050\
        );

    \I__1483\ : InMux
    port map (
            O => \N__6092\,
            I => \N__6047\
        );

    \I__1482\ : Span4Mux_v
    port map (
            O => \N__6085\,
            I => \N__6044\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__6082\,
            I => \N__6041\
        );

    \I__1480\ : InMux
    port map (
            O => \N__6081\,
            I => \N__6038\
        );

    \I__1479\ : InMux
    port map (
            O => \N__6080\,
            I => \N__6035\
        );

    \I__1478\ : InMux
    port map (
            O => \N__6079\,
            I => \N__6032\
        );

    \I__1477\ : InMux
    port map (
            O => \N__6078\,
            I => \N__6029\
        );

    \I__1476\ : InMux
    port map (
            O => \N__6077\,
            I => \N__6026\
        );

    \I__1475\ : InMux
    port map (
            O => \N__6076\,
            I => \N__6022\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__6073\,
            I => \N__6019\
        );

    \I__1473\ : Span4Mux_v
    port map (
            O => \N__6068\,
            I => \N__6016\
        );

    \I__1472\ : InMux
    port map (
            O => \N__6067\,
            I => \N__6013\
        );

    \I__1471\ : Sp12to4
    port map (
            O => \N__6064\,
            I => \N__6008\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__6061\,
            I => \N__6008\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__6058\,
            I => \N__6003\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__6055\,
            I => \N__6003\
        );

    \I__1467\ : InMux
    port map (
            O => \N__6054\,
            I => \N__6000\
        );

    \I__1466\ : InMux
    port map (
            O => \N__6053\,
            I => \N__5997\
        );

    \I__1465\ : Span4Mux_v
    port map (
            O => \N__6050\,
            I => \N__5992\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__6047\,
            I => \N__5992\
        );

    \I__1463\ : Span4Mux_v
    port map (
            O => \N__6044\,
            I => \N__5977\
        );

    \I__1462\ : Span4Mux_v
    port map (
            O => \N__6041\,
            I => \N__5977\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__6038\,
            I => \N__5977\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__6035\,
            I => \N__5977\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__6032\,
            I => \N__5977\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__6029\,
            I => \N__5977\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__6026\,
            I => \N__5977\
        );

    \I__1456\ : InMux
    port map (
            O => \N__6025\,
            I => \N__5974\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__6022\,
            I => \N__5970\
        );

    \I__1454\ : Span12Mux_s10_v
    port map (
            O => \N__6019\,
            I => \N__5960\
        );

    \I__1453\ : Sp12to4
    port map (
            O => \N__6016\,
            I => \N__5960\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__6013\,
            I => \N__5960\
        );

    \I__1451\ : Span12Mux_h
    port map (
            O => \N__6008\,
            I => \N__5953\
        );

    \I__1450\ : Span12Mux_s10_v
    port map (
            O => \N__6003\,
            I => \N__5953\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__6000\,
            I => \N__5953\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__5997\,
            I => \N__5950\
        );

    \I__1447\ : Span4Mux_v
    port map (
            O => \N__5992\,
            I => \N__5947\
        );

    \I__1446\ : Span4Mux_v
    port map (
            O => \N__5977\,
            I => \N__5942\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__5974\,
            I => \N__5942\
        );

    \I__1444\ : InMux
    port map (
            O => \N__5973\,
            I => \N__5939\
        );

    \I__1443\ : Span4Mux_h
    port map (
            O => \N__5970\,
            I => \N__5936\
        );

    \I__1442\ : InMux
    port map (
            O => \N__5969\,
            I => \N__5931\
        );

    \I__1441\ : InMux
    port map (
            O => \N__5968\,
            I => \N__5931\
        );

    \I__1440\ : InMux
    port map (
            O => \N__5967\,
            I => \N__5927\
        );

    \I__1439\ : Span12Mux_v
    port map (
            O => \N__5960\,
            I => \N__5924\
        );

    \I__1438\ : Span12Mux_v
    port map (
            O => \N__5953\,
            I => \N__5921\
        );

    \I__1437\ : Span4Mux_v
    port map (
            O => \N__5950\,
            I => \N__5918\
        );

    \I__1436\ : Span4Mux_h
    port map (
            O => \N__5947\,
            I => \N__5913\
        );

    \I__1435\ : Span4Mux_v
    port map (
            O => \N__5942\,
            I => \N__5913\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__5939\,
            I => \N__5910\
        );

    \I__1433\ : Span4Mux_h
    port map (
            O => \N__5936\,
            I => \N__5905\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__5931\,
            I => \N__5905\
        );

    \I__1431\ : InMux
    port map (
            O => \N__5930\,
            I => \N__5902\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__5927\,
            I => \N__5899\
        );

    \I__1429\ : Odrv12
    port map (
            O => \N__5924\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__1428\ : Odrv12
    port map (
            O => \N__5921\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__1427\ : Odrv4
    port map (
            O => \N__5918\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__1426\ : Odrv4
    port map (
            O => \N__5913\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__1425\ : Odrv4
    port map (
            O => \N__5910\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__1424\ : Odrv4
    port map (
            O => \N__5905\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__5902\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__1422\ : Odrv4
    port map (
            O => \N__5899\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__1421\ : IoInMux
    port map (
            O => \N__5882\,
            I => \N__5879\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__5879\,
            I => \N__5876\
        );

    \I__1419\ : IoSpan4Mux
    port map (
            O => \N__5876\,
            I => \N__5873\
        );

    \I__1418\ : IoSpan4Mux
    port map (
            O => \N__5873\,
            I => \N__5870\
        );

    \I__1417\ : Sp12to4
    port map (
            O => \N__5870\,
            I => \N__5867\
        );

    \I__1416\ : Span12Mux_s6_v
    port map (
            O => \N__5867\,
            I => \N__5864\
        );

    \I__1415\ : Odrv12
    port map (
            O => \N__5864\,
            I => \un1_D_UU_040_4\
        );

    \I__1414\ : InMux
    port map (
            O => \N__5861\,
            I => \N__5858\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__5858\,
            I => \N__5854\
        );

    \I__1412\ : InMux
    port map (
            O => \N__5857\,
            I => \N__5851\
        );

    \I__1411\ : Span4Mux_v
    port map (
            O => \N__5854\,
            I => \N__5847\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__5851\,
            I => \N__5844\
        );

    \I__1409\ : InMux
    port map (
            O => \N__5850\,
            I => \N__5841\
        );

    \I__1408\ : Span4Mux_v
    port map (
            O => \N__5847\,
            I => \N__5838\
        );

    \I__1407\ : Span4Mux_v
    port map (
            O => \N__5844\,
            I => \N__5833\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__5841\,
            I => \N__5833\
        );

    \I__1405\ : Sp12to4
    port map (
            O => \N__5838\,
            I => \N__5830\
        );

    \I__1404\ : Sp12to4
    port map (
            O => \N__5833\,
            I => \N__5827\
        );

    \I__1403\ : Span12Mux_h
    port map (
            O => \N__5830\,
            I => \N__5824\
        );

    \I__1402\ : Span12Mux_v
    port map (
            O => \N__5827\,
            I => \N__5821\
        );

    \I__1401\ : Span12Mux_v
    port map (
            O => \N__5824\,
            I => \N__5816\
        );

    \I__1400\ : Span12Mux_h
    port map (
            O => \N__5821\,
            I => \N__5816\
        );

    \I__1399\ : Odrv12
    port map (
            O => \N__5816\,
            I => \D_UM_AMIGA_in_3\
        );

    \I__1398\ : InMux
    port map (
            O => \N__5813\,
            I => \N__5810\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__5810\,
            I => \N__5807\
        );

    \I__1396\ : Odrv12
    port map (
            O => \N__5807\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\
        );

    \I__1395\ : IoInMux
    port map (
            O => \N__5804\,
            I => \N__5801\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__5801\,
            I => \N__5798\
        );

    \I__1393\ : IoSpan4Mux
    port map (
            O => \N__5798\,
            I => \N__5795\
        );

    \I__1392\ : Span4Mux_s1_h
    port map (
            O => \N__5795\,
            I => \N__5792\
        );

    \I__1391\ : Sp12to4
    port map (
            O => \N__5792\,
            I => \N__5789\
        );

    \I__1390\ : Span12Mux_h
    port map (
            O => \N__5789\,
            I => \N__5786\
        );

    \I__1389\ : Odrv12
    port map (
            O => \N__5786\,
            I => \un1_D_UM_AMIGA_3\
        );

    \I__1388\ : InMux
    port map (
            O => \N__5783\,
            I => \N__5779\
        );

    \I__1387\ : IoInMux
    port map (
            O => \N__5782\,
            I => \N__5776\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__5779\,
            I => \N__5773\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__5776\,
            I => \N__5770\
        );

    \I__1384\ : Span4Mux_v
    port map (
            O => \N__5773\,
            I => \N__5767\
        );

    \I__1383\ : Span4Mux_s3_h
    port map (
            O => \N__5770\,
            I => \N__5764\
        );

    \I__1382\ : Sp12to4
    port map (
            O => \N__5767\,
            I => \N__5761\
        );

    \I__1381\ : Sp12to4
    port map (
            O => \N__5764\,
            I => \N__5758\
        );

    \I__1380\ : Span12Mux_h
    port map (
            O => \N__5761\,
            I => \N__5755\
        );

    \I__1379\ : Span12Mux_v
    port map (
            O => \N__5758\,
            I => \N__5752\
        );

    \I__1378\ : Span12Mux_v
    port map (
            O => \N__5755\,
            I => \N__5749\
        );

    \I__1377\ : Span12Mux_h
    port map (
            O => \N__5752\,
            I => \N__5746\
        );

    \I__1376\ : Span12Mux_v
    port map (
            O => \N__5749\,
            I => \N__5741\
        );

    \I__1375\ : Span12Mux_h
    port map (
            O => \N__5746\,
            I => \N__5741\
        );

    \I__1374\ : Odrv12
    port map (
            O => \N__5741\,
            I => \D_LL_040_in_3\
        );

    \I__1373\ : InMux
    port map (
            O => \N__5738\,
            I => \N__5735\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__5735\,
            I => \N__5732\
        );

    \I__1371\ : Sp12to4
    port map (
            O => \N__5732\,
            I => \N__5729\
        );

    \I__1370\ : Span12Mux_v
    port map (
            O => \N__5729\,
            I => \N__5726\
        );

    \I__1369\ : Span12Mux_h
    port map (
            O => \N__5726\,
            I => \N__5723\
        );

    \I__1368\ : Odrv12
    port map (
            O => \N__5723\,
            I => \D_UM_040_in_3\
        );

    \I__1367\ : IoInMux
    port map (
            O => \N__5720\,
            I => \N__5717\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__5717\,
            I => \N__5714\
        );

    \I__1365\ : IoSpan4Mux
    port map (
            O => \N__5714\,
            I => \N__5711\
        );

    \I__1364\ : Span4Mux_s3_h
    port map (
            O => \N__5711\,
            I => \N__5708\
        );

    \I__1363\ : Sp12to4
    port map (
            O => \N__5708\,
            I => \N__5705\
        );

    \I__1362\ : Span12Mux_h
    port map (
            O => \N__5705\,
            I => \N__5702\
        );

    \I__1361\ : Odrv12
    port map (
            O => \N__5702\,
            I => \un1_D_UM_040_3\
        );

    \I__1360\ : InMux
    port map (
            O => \N__5699\,
            I => \N__5696\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__5696\,
            I => \N__5691\
        );

    \I__1358\ : InMux
    port map (
            O => \N__5695\,
            I => \N__5688\
        );

    \I__1357\ : InMux
    port map (
            O => \N__5694\,
            I => \N__5685\
        );

    \I__1356\ : Span4Mux_h
    port map (
            O => \N__5691\,
            I => \N__5682\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__5688\,
            I => \N__5679\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__5685\,
            I => \N__5676\
        );

    \I__1353\ : Span4Mux_v
    port map (
            O => \N__5682\,
            I => \N__5671\
        );

    \I__1352\ : Span4Mux_h
    port map (
            O => \N__5679\,
            I => \N__5671\
        );

    \I__1351\ : Sp12to4
    port map (
            O => \N__5676\,
            I => \N__5668\
        );

    \I__1350\ : Span4Mux_v
    port map (
            O => \N__5671\,
            I => \N__5665\
        );

    \I__1349\ : Span12Mux_v
    port map (
            O => \N__5668\,
            I => \N__5662\
        );

    \I__1348\ : Sp12to4
    port map (
            O => \N__5665\,
            I => \N__5659\
        );

    \I__1347\ : Span12Mux_v
    port map (
            O => \N__5662\,
            I => \N__5656\
        );

    \I__1346\ : Span12Mux_h
    port map (
            O => \N__5659\,
            I => \N__5653\
        );

    \I__1345\ : Odrv12
    port map (
            O => \N__5656\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__1344\ : Odrv12
    port map (
            O => \N__5653\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__1343\ : InMux
    port map (
            O => \N__5648\,
            I => \N__5645\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__5645\,
            I => \N__5642\
        );

    \I__1341\ : Odrv12
    port map (
            O => \N__5642\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\
        );

    \I__1340\ : IoInMux
    port map (
            O => \N__5639\,
            I => \N__5636\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__5636\,
            I => \N__5633\
        );

    \I__1338\ : Span4Mux_s3_h
    port map (
            O => \N__5633\,
            I => \N__5630\
        );

    \I__1337\ : Sp12to4
    port map (
            O => \N__5630\,
            I => \N__5627\
        );

    \I__1336\ : Span12Mux_v
    port map (
            O => \N__5627\,
            I => \N__5624\
        );

    \I__1335\ : Span12Mux_h
    port map (
            O => \N__5624\,
            I => \N__5621\
        );

    \I__1334\ : Odrv12
    port map (
            O => \N__5621\,
            I => \un1_D_UM_AMIGA_7\
        );

    \I__1333\ : InMux
    port map (
            O => \N__5618\,
            I => \N__5615\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__5615\,
            I => \N__5612\
        );

    \I__1331\ : Odrv12
    port map (
            O => \N__5612\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\
        );

    \I__1330\ : InMux
    port map (
            O => \N__5609\,
            I => \N__5605\
        );

    \I__1329\ : InMux
    port map (
            O => \N__5608\,
            I => \N__5602\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__5605\,
            I => \N__5599\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__5602\,
            I => \N__5596\
        );

    \I__1326\ : Span4Mux_v
    port map (
            O => \N__5599\,
            I => \N__5593\
        );

    \I__1325\ : Span4Mux_v
    port map (
            O => \N__5596\,
            I => \N__5590\
        );

    \I__1324\ : Span4Mux_v
    port map (
            O => \N__5593\,
            I => \N__5586\
        );

    \I__1323\ : Span4Mux_v
    port map (
            O => \N__5590\,
            I => \N__5583\
        );

    \I__1322\ : InMux
    port map (
            O => \N__5589\,
            I => \N__5580\
        );

    \I__1321\ : Sp12to4
    port map (
            O => \N__5586\,
            I => \N__5573\
        );

    \I__1320\ : Sp12to4
    port map (
            O => \N__5583\,
            I => \N__5573\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__5580\,
            I => \N__5573\
        );

    \I__1318\ : Span12Mux_h
    port map (
            O => \N__5573\,
            I => \N__5570\
        );

    \I__1317\ : Odrv12
    port map (
            O => \N__5570\,
            I => \D_UU_AMIGA_in_2\
        );

    \I__1316\ : IoInMux
    port map (
            O => \N__5567\,
            I => \N__5564\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__5564\,
            I => \N__5561\
        );

    \I__1314\ : IoSpan4Mux
    port map (
            O => \N__5561\,
            I => \N__5558\
        );

    \I__1313\ : IoSpan4Mux
    port map (
            O => \N__5558\,
            I => \N__5555\
        );

    \I__1312\ : Span4Mux_s3_v
    port map (
            O => \N__5555\,
            I => \N__5552\
        );

    \I__1311\ : Span4Mux_v
    port map (
            O => \N__5552\,
            I => \N__5549\
        );

    \I__1310\ : Odrv4
    port map (
            O => \N__5549\,
            I => \un1_D_UU_AMIGA_2\
        );

    \I__1309\ : InMux
    port map (
            O => \N__5546\,
            I => \N__5543\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__5543\,
            I => \N__5540\
        );

    \I__1307\ : Span4Mux_v
    port map (
            O => \N__5540\,
            I => \N__5537\
        );

    \I__1306\ : Odrv4
    port map (
            O => \N__5537\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\
        );

    \I__1305\ : InMux
    port map (
            O => \N__5534\,
            I => \N__5530\
        );

    \I__1304\ : InMux
    port map (
            O => \N__5533\,
            I => \N__5526\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__5530\,
            I => \N__5523\
        );

    \I__1302\ : InMux
    port map (
            O => \N__5529\,
            I => \N__5520\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__5526\,
            I => \N__5517\
        );

    \I__1300\ : Span4Mux_h
    port map (
            O => \N__5523\,
            I => \N__5512\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__5520\,
            I => \N__5512\
        );

    \I__1298\ : Span4Mux_v
    port map (
            O => \N__5517\,
            I => \N__5509\
        );

    \I__1297\ : Span4Mux_h
    port map (
            O => \N__5512\,
            I => \N__5506\
        );

    \I__1296\ : Span4Mux_v
    port map (
            O => \N__5509\,
            I => \N__5503\
        );

    \I__1295\ : Sp12to4
    port map (
            O => \N__5506\,
            I => \N__5500\
        );

    \I__1294\ : Sp12to4
    port map (
            O => \N__5503\,
            I => \N__5497\
        );

    \I__1293\ : Span12Mux_v
    port map (
            O => \N__5500\,
            I => \N__5494\
        );

    \I__1292\ : Span12Mux_h
    port map (
            O => \N__5497\,
            I => \N__5491\
        );

    \I__1291\ : Odrv12
    port map (
            O => \N__5494\,
            I => \D_UU_AMIGA_in_5\
        );

    \I__1290\ : Odrv12
    port map (
            O => \N__5491\,
            I => \D_UU_AMIGA_in_5\
        );

    \I__1289\ : IoInMux
    port map (
            O => \N__5486\,
            I => \N__5483\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__5483\,
            I => \N__5480\
        );

    \I__1287\ : Span4Mux_s3_v
    port map (
            O => \N__5480\,
            I => \N__5477\
        );

    \I__1286\ : Span4Mux_v
    port map (
            O => \N__5477\,
            I => \N__5474\
        );

    \I__1285\ : Sp12to4
    port map (
            O => \N__5474\,
            I => \N__5471\
        );

    \I__1284\ : Odrv12
    port map (
            O => \N__5471\,
            I => \un1_D_UU_AMIGA_5\
        );

    \I__1283\ : InMux
    port map (
            O => \N__5468\,
            I => \N__5465\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__5465\,
            I => \N__5462\
        );

    \I__1281\ : Odrv12
    port map (
            O => \N__5462\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\
        );

    \I__1280\ : InMux
    port map (
            O => \N__5459\,
            I => \N__5455\
        );

    \I__1279\ : InMux
    port map (
            O => \N__5458\,
            I => \N__5452\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__5455\,
            I => \N__5448\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__5452\,
            I => \N__5445\
        );

    \I__1276\ : InMux
    port map (
            O => \N__5451\,
            I => \N__5442\
        );

    \I__1275\ : Span4Mux_v
    port map (
            O => \N__5448\,
            I => \N__5439\
        );

    \I__1274\ : Span4Mux_v
    port map (
            O => \N__5445\,
            I => \N__5434\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__5442\,
            I => \N__5434\
        );

    \I__1272\ : Span4Mux_v
    port map (
            O => \N__5439\,
            I => \N__5431\
        );

    \I__1271\ : Span4Mux_v
    port map (
            O => \N__5434\,
            I => \N__5428\
        );

    \I__1270\ : Span4Mux_v
    port map (
            O => \N__5431\,
            I => \N__5423\
        );

    \I__1269\ : Span4Mux_h
    port map (
            O => \N__5428\,
            I => \N__5423\
        );

    \I__1268\ : Sp12to4
    port map (
            O => \N__5423\,
            I => \N__5420\
        );

    \I__1267\ : Span12Mux_h
    port map (
            O => \N__5420\,
            I => \N__5417\
        );

    \I__1266\ : Odrv12
    port map (
            O => \N__5417\,
            I => \D_UU_AMIGA_in_3\
        );

    \I__1265\ : IoInMux
    port map (
            O => \N__5414\,
            I => \N__5411\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__5411\,
            I => \N__5408\
        );

    \I__1263\ : IoSpan4Mux
    port map (
            O => \N__5408\,
            I => \N__5405\
        );

    \I__1262\ : IoSpan4Mux
    port map (
            O => \N__5405\,
            I => \N__5402\
        );

    \I__1261\ : Sp12to4
    port map (
            O => \N__5402\,
            I => \N__5399\
        );

    \I__1260\ : Span12Mux_s7_h
    port map (
            O => \N__5399\,
            I => \N__5396\
        );

    \I__1259\ : Odrv12
    port map (
            O => \N__5396\,
            I => \un1_D_UU_AMIGA_3\
        );

    \I__1258\ : InMux
    port map (
            O => \N__5393\,
            I => \N__5390\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__5390\,
            I => \N__5387\
        );

    \I__1256\ : Span12Mux_v
    port map (
            O => \N__5387\,
            I => \N__5384\
        );

    \I__1255\ : Span12Mux_h
    port map (
            O => \N__5384\,
            I => \N__5381\
        );

    \I__1254\ : Odrv12
    port map (
            O => \N__5381\,
            I => \D_UU_040_in_6\
        );

    \I__1253\ : IoInMux
    port map (
            O => \N__5378\,
            I => \N__5375\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__5375\,
            I => \N__5372\
        );

    \I__1251\ : Span4Mux_s2_h
    port map (
            O => \N__5372\,
            I => \N__5368\
        );

    \I__1250\ : InMux
    port map (
            O => \N__5371\,
            I => \N__5365\
        );

    \I__1249\ : Span4Mux_v
    port map (
            O => \N__5368\,
            I => \N__5362\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__5365\,
            I => \N__5359\
        );

    \I__1247\ : Sp12to4
    port map (
            O => \N__5362\,
            I => \N__5356\
        );

    \I__1246\ : Sp12to4
    port map (
            O => \N__5359\,
            I => \N__5353\
        );

    \I__1245\ : Span12Mux_h
    port map (
            O => \N__5356\,
            I => \N__5350\
        );

    \I__1244\ : Span12Mux_s11_v
    port map (
            O => \N__5353\,
            I => \N__5347\
        );

    \I__1243\ : Span12Mux_h
    port map (
            O => \N__5350\,
            I => \N__5344\
        );

    \I__1242\ : Span12Mux_h
    port map (
            O => \N__5347\,
            I => \N__5341\
        );

    \I__1241\ : Odrv12
    port map (
            O => \N__5344\,
            I => \D_LM_040_in_6\
        );

    \I__1240\ : Odrv12
    port map (
            O => \N__5341\,
            I => \D_LM_040_in_6\
        );

    \I__1239\ : IoInMux
    port map (
            O => \N__5336\,
            I => \N__5333\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__5333\,
            I => \N__5330\
        );

    \I__1237\ : Span4Mux_s2_v
    port map (
            O => \N__5330\,
            I => \N__5327\
        );

    \I__1236\ : Span4Mux_v
    port map (
            O => \N__5327\,
            I => \N__5324\
        );

    \I__1235\ : Sp12to4
    port map (
            O => \N__5324\,
            I => \N__5321\
        );

    \I__1234\ : Span12Mux_s11_h
    port map (
            O => \N__5321\,
            I => \N__5318\
        );

    \I__1233\ : Odrv12
    port map (
            O => \N__5318\,
            I => \un1_D_UU_040_6\
        );

    \I__1232\ : InMux
    port map (
            O => \N__5315\,
            I => \N__5312\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__5312\,
            I => \N__5309\
        );

    \I__1230\ : Span4Mux_v
    port map (
            O => \N__5309\,
            I => \N__5306\
        );

    \I__1229\ : Odrv4
    port map (
            O => \N__5306\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\
        );

    \I__1228\ : CEMux
    port map (
            O => \N__5303\,
            I => \N__5295\
        );

    \I__1227\ : CEMux
    port map (
            O => \N__5302\,
            I => \N__5292\
        );

    \I__1226\ : CEMux
    port map (
            O => \N__5301\,
            I => \N__5289\
        );

    \I__1225\ : CEMux
    port map (
            O => \N__5300\,
            I => \N__5286\
        );

    \I__1224\ : CEMux
    port map (
            O => \N__5299\,
            I => \N__5283\
        );

    \I__1223\ : CEMux
    port map (
            O => \N__5298\,
            I => \N__5280\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__5295\,
            I => \N__5275\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__5292\,
            I => \N__5275\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__5289\,
            I => \N__5272\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__5286\,
            I => \N__5265\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__5283\,
            I => \N__5265\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__5280\,
            I => \N__5265\
        );

    \I__1216\ : Odrv4
    port map (
            O => \N__5275\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\
        );

    \I__1215\ : Odrv4
    port map (
            O => \N__5272\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\
        );

    \I__1214\ : Odrv4
    port map (
            O => \N__5265\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\
        );

    \I__1213\ : SRMux
    port map (
            O => \N__5258\,
            I => \N__5255\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__5255\,
            I => \N__5248\
        );

    \I__1211\ : SRMux
    port map (
            O => \N__5254\,
            I => \N__5245\
        );

    \I__1210\ : SRMux
    port map (
            O => \N__5253\,
            I => \N__5242\
        );

    \I__1209\ : SRMux
    port map (
            O => \N__5252\,
            I => \N__5239\
        );

    \I__1208\ : SRMux
    port map (
            O => \N__5251\,
            I => \N__5235\
        );

    \I__1207\ : Span4Mux_h
    port map (
            O => \N__5248\,
            I => \N__5230\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__5245\,
            I => \N__5230\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__5242\,
            I => \N__5227\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__5239\,
            I => \N__5224\
        );

    \I__1203\ : SRMux
    port map (
            O => \N__5238\,
            I => \N__5221\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__5235\,
            I => \N__5218\
        );

    \I__1201\ : Span4Mux_h
    port map (
            O => \N__5230\,
            I => \N__5213\
        );

    \I__1200\ : Span4Mux_h
    port map (
            O => \N__5227\,
            I => \N__5213\
        );

    \I__1199\ : Span4Mux_v
    port map (
            O => \N__5224\,
            I => \N__5206\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__5221\,
            I => \N__5206\
        );

    \I__1197\ : Span4Mux_h
    port map (
            O => \N__5218\,
            I => \N__5206\
        );

    \I__1196\ : Odrv4
    port map (
            O => \N__5213\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0\
        );

    \I__1195\ : Odrv4
    port map (
            O => \N__5206\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0\
        );

    \I__1194\ : InMux
    port map (
            O => \N__5201\,
            I => \N__5198\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__5198\,
            I => \N__5193\
        );

    \I__1192\ : InMux
    port map (
            O => \N__5197\,
            I => \N__5190\
        );

    \I__1191\ : InMux
    port map (
            O => \N__5196\,
            I => \N__5187\
        );

    \I__1190\ : Span4Mux_v
    port map (
            O => \N__5193\,
            I => \N__5184\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5190\,
            I => \N__5179\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__5187\,
            I => \N__5179\
        );

    \I__1187\ : Sp12to4
    port map (
            O => \N__5184\,
            I => \N__5176\
        );

    \I__1186\ : Span4Mux_v
    port map (
            O => \N__5179\,
            I => \N__5173\
        );

    \I__1185\ : Span12Mux_h
    port map (
            O => \N__5176\,
            I => \N__5170\
        );

    \I__1184\ : Sp12to4
    port map (
            O => \N__5173\,
            I => \N__5167\
        );

    \I__1183\ : Span12Mux_v
    port map (
            O => \N__5170\,
            I => \N__5162\
        );

    \I__1182\ : Span12Mux_h
    port map (
            O => \N__5167\,
            I => \N__5162\
        );

    \I__1181\ : Odrv12
    port map (
            O => \N__5162\,
            I => \D_UM_AMIGA_in_1\
        );

    \I__1180\ : InMux
    port map (
            O => \N__5159\,
            I => \N__5156\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__5156\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\
        );

    \I__1178\ : IoInMux
    port map (
            O => \N__5153\,
            I => \N__5150\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__5150\,
            I => \N__5147\
        );

    \I__1176\ : Span4Mux_s3_h
    port map (
            O => \N__5147\,
            I => \N__5144\
        );

    \I__1175\ : Sp12to4
    port map (
            O => \N__5144\,
            I => \N__5141\
        );

    \I__1174\ : Span12Mux_s11_v
    port map (
            O => \N__5141\,
            I => \N__5138\
        );

    \I__1173\ : Odrv12
    port map (
            O => \N__5138\,
            I => \un1_D_UM_AMIGA_1\
        );

    \I__1172\ : IoInMux
    port map (
            O => \N__5135\,
            I => \N__5132\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__5132\,
            I => \N__5129\
        );

    \I__1170\ : Span4Mux_s2_v
    port map (
            O => \N__5129\,
            I => \N__5126\
        );

    \I__1169\ : Span4Mux_v
    port map (
            O => \N__5126\,
            I => \N__5123\
        );

    \I__1168\ : Sp12to4
    port map (
            O => \N__5123\,
            I => \N__5120\
        );

    \I__1167\ : Span12Mux_s11_h
    port map (
            O => \N__5120\,
            I => \N__5117\
        );

    \I__1166\ : Odrv12
    port map (
            O => \N__5117\,
            I => \un1_D_UM_040_5\
        );

    \I__1165\ : InMux
    port map (
            O => \N__5114\,
            I => \N__5111\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__5111\,
            I => \N__5108\
        );

    \I__1163\ : Span4Mux_v
    port map (
            O => \N__5108\,
            I => \N__5105\
        );

    \I__1162\ : Odrv4
    port map (
            O => \N__5105\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\
        );

    \I__1161\ : InMux
    port map (
            O => \N__5102\,
            I => \N__5099\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__5099\,
            I => \N__5096\
        );

    \I__1159\ : Span4Mux_v
    port map (
            O => \N__5096\,
            I => \N__5091\
        );

    \I__1158\ : InMux
    port map (
            O => \N__5095\,
            I => \N__5088\
        );

    \I__1157\ : InMux
    port map (
            O => \N__5094\,
            I => \N__5085\
        );

    \I__1156\ : Span4Mux_v
    port map (
            O => \N__5091\,
            I => \N__5082\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__5088\,
            I => \N__5079\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__5085\,
            I => \N__5076\
        );

    \I__1153\ : Span4Mux_v
    port map (
            O => \N__5082\,
            I => \N__5073\
        );

    \I__1152\ : Span4Mux_v
    port map (
            O => \N__5079\,
            I => \N__5068\
        );

    \I__1151\ : Span4Mux_v
    port map (
            O => \N__5076\,
            I => \N__5068\
        );

    \I__1150\ : Sp12to4
    port map (
            O => \N__5073\,
            I => \N__5063\
        );

    \I__1149\ : Sp12to4
    port map (
            O => \N__5068\,
            I => \N__5063\
        );

    \I__1148\ : Span12Mux_h
    port map (
            O => \N__5063\,
            I => \N__5060\
        );

    \I__1147\ : Odrv12
    port map (
            O => \N__5060\,
            I => \D_UU_AMIGA_in_0\
        );

    \I__1146\ : IoInMux
    port map (
            O => \N__5057\,
            I => \N__5054\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__5054\,
            I => \N__5051\
        );

    \I__1144\ : Span12Mux_s8_v
    port map (
            O => \N__5051\,
            I => \N__5048\
        );

    \I__1143\ : Span12Mux_h
    port map (
            O => \N__5048\,
            I => \N__5045\
        );

    \I__1142\ : Odrv12
    port map (
            O => \N__5045\,
            I => \un1_D_UU_AMIGA_0\
        );

    \I__1141\ : IoInMux
    port map (
            O => \N__5042\,
            I => \N__5038\
        );

    \I__1140\ : IoInMux
    port map (
            O => \N__5041\,
            I => \N__5035\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__5038\,
            I => \N__5032\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__5035\,
            I => \N__5029\
        );

    \I__1137\ : Span12Mux_s6_v
    port map (
            O => \N__5032\,
            I => \N__5024\
        );

    \I__1136\ : Span12Mux_s6_v
    port map (
            O => \N__5029\,
            I => \N__5024\
        );

    \I__1135\ : Odrv12
    port map (
            O => \N__5024\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1134\ : InMux
    port map (
            O => \N__5021\,
            I => \N__5018\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__5018\,
            I => \N__5015\
        );

    \I__1132\ : Span4Mux_v
    port map (
            O => \N__5015\,
            I => \N__5012\
        );

    \I__1131\ : Sp12to4
    port map (
            O => \N__5012\,
            I => \N__5009\
        );

    \I__1130\ : Span12Mux_h
    port map (
            O => \N__5009\,
            I => \N__5006\
        );

    \I__1129\ : Odrv12
    port map (
            O => \N__5006\,
            I => \D_LL_AMIGA_in_2\
        );

    \I__1128\ : IoInMux
    port map (
            O => \N__5003\,
            I => \N__5000\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__5000\,
            I => \N__4997\
        );

    \I__1126\ : IoSpan4Mux
    port map (
            O => \N__4997\,
            I => \N__4994\
        );

    \I__1125\ : Span4Mux_s1_h
    port map (
            O => \N__4994\,
            I => \N__4991\
        );

    \I__1124\ : Sp12to4
    port map (
            O => \N__4991\,
            I => \N__4988\
        );

    \I__1123\ : Span12Mux_h
    port map (
            O => \N__4988\,
            I => \N__4985\
        );

    \I__1122\ : Odrv12
    port map (
            O => \N__4985\,
            I => \un1_D_LL_AMIGA_2\
        );

    \I__1121\ : InMux
    port map (
            O => \N__4982\,
            I => \N__4979\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__4979\,
            I => \N__4976\
        );

    \I__1119\ : Span4Mux_v
    port map (
            O => \N__4976\,
            I => \N__4973\
        );

    \I__1118\ : Sp12to4
    port map (
            O => \N__4973\,
            I => \N__4970\
        );

    \I__1117\ : Span12Mux_h
    port map (
            O => \N__4970\,
            I => \N__4967\
        );

    \I__1116\ : Odrv12
    port map (
            O => \N__4967\,
            I => \D_LL_AMIGA_in_6\
        );

    \I__1115\ : IoInMux
    port map (
            O => \N__4964\,
            I => \N__4961\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__4961\,
            I => \N__4958\
        );

    \I__1113\ : Span4Mux_s3_h
    port map (
            O => \N__4958\,
            I => \N__4955\
        );

    \I__1112\ : Sp12to4
    port map (
            O => \N__4955\,
            I => \N__4952\
        );

    \I__1111\ : Span12Mux_s9_v
    port map (
            O => \N__4952\,
            I => \N__4949\
        );

    \I__1110\ : Span12Mux_h
    port map (
            O => \N__4949\,
            I => \N__4946\
        );

    \I__1109\ : Odrv12
    port map (
            O => \N__4946\,
            I => \un1_D_LL_AMIGA_6\
        );

    \I__1108\ : IoInMux
    port map (
            O => \N__4943\,
            I => \N__4940\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__4940\,
            I => \N__4937\
        );

    \I__1106\ : Span12Mux_s7_h
    port map (
            O => \N__4937\,
            I => \N__4934\
        );

    \I__1105\ : Odrv12
    port map (
            O => \N__4934\,
            I => \un1_D_UM_AMIGA_2\
        );

    \I__1104\ : InMux
    port map (
            O => \N__4931\,
            I => \N__4928\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__4928\,
            I => \N__4924\
        );

    \I__1102\ : ClkMux
    port map (
            O => \N__4927\,
            I => \N__4892\
        );

    \I__1101\ : Glb2LocalMux
    port map (
            O => \N__4924\,
            I => \N__4892\
        );

    \I__1100\ : ClkMux
    port map (
            O => \N__4923\,
            I => \N__4892\
        );

    \I__1099\ : ClkMux
    port map (
            O => \N__4922\,
            I => \N__4892\
        );

    \I__1098\ : ClkMux
    port map (
            O => \N__4921\,
            I => \N__4892\
        );

    \I__1097\ : ClkMux
    port map (
            O => \N__4920\,
            I => \N__4892\
        );

    \I__1096\ : ClkMux
    port map (
            O => \N__4919\,
            I => \N__4892\
        );

    \I__1095\ : ClkMux
    port map (
            O => \N__4918\,
            I => \N__4892\
        );

    \I__1094\ : ClkMux
    port map (
            O => \N__4917\,
            I => \N__4892\
        );

    \I__1093\ : ClkMux
    port map (
            O => \N__4916\,
            I => \N__4892\
        );

    \I__1092\ : ClkMux
    port map (
            O => \N__4915\,
            I => \N__4892\
        );

    \I__1091\ : GlobalMux
    port map (
            O => \N__4892\,
            I => \CLK80\
        );

    \I__1090\ : IoInMux
    port map (
            O => \N__4889\,
            I => \N__4886\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__4886\,
            I => \N__4883\
        );

    \I__1088\ : IoSpan4Mux
    port map (
            O => \N__4883\,
            I => \N__4880\
        );

    \I__1087\ : IoSpan4Mux
    port map (
            O => \N__4880\,
            I => \N__4875\
        );

    \I__1086\ : IoInMux
    port map (
            O => \N__4879\,
            I => \N__4872\
        );

    \I__1085\ : IoInMux
    port map (
            O => \N__4878\,
            I => \N__4869\
        );

    \I__1084\ : Sp12to4
    port map (
            O => \N__4875\,
            I => \N__4864\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__4872\,
            I => \N__4864\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__4869\,
            I => \N__4861\
        );

    \I__1081\ : Span12Mux_s7_v
    port map (
            O => \N__4864\,
            I => \N__4858\
        );

    \I__1080\ : Span12Mux_s10_h
    port map (
            O => \N__4861\,
            I => \N__4855\
        );

    \I__1079\ : Odrv12
    port map (
            O => \N__4858\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__1078\ : Odrv12
    port map (
            O => \N__4855\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__1077\ : InMux
    port map (
            O => \N__4850\,
            I => \N__4846\
        );

    \I__1076\ : InMux
    port map (
            O => \N__4849\,
            I => \N__4842\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__4846\,
            I => \N__4839\
        );

    \I__1074\ : InMux
    port map (
            O => \N__4845\,
            I => \N__4836\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__4842\,
            I => \N__4833\
        );

    \I__1072\ : Span4Mux_h
    port map (
            O => \N__4839\,
            I => \N__4828\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__4836\,
            I => \N__4828\
        );

    \I__1070\ : Sp12to4
    port map (
            O => \N__4833\,
            I => \N__4825\
        );

    \I__1069\ : Span4Mux_v
    port map (
            O => \N__4828\,
            I => \N__4822\
        );

    \I__1068\ : Span12Mux_v
    port map (
            O => \N__4825\,
            I => \N__4817\
        );

    \I__1067\ : Sp12to4
    port map (
            O => \N__4822\,
            I => \N__4817\
        );

    \I__1066\ : Span12Mux_h
    port map (
            O => \N__4817\,
            I => \N__4814\
        );

    \I__1065\ : Odrv12
    port map (
            O => \N__4814\,
            I => \D_UM_AMIGA_in_2\
        );

    \I__1064\ : InMux
    port map (
            O => \N__4811\,
            I => \N__4808\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__4808\,
            I => \N__4805\
        );

    \I__1062\ : Odrv4
    port map (
            O => \N__4805\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\
        );

    \I__1061\ : InMux
    port map (
            O => \N__4802\,
            I => \N__4798\
        );

    \I__1060\ : InMux
    port map (
            O => \N__4801\,
            I => \N__4795\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__4798\,
            I => \N__4792\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__4795\,
            I => \N__4788\
        );

    \I__1057\ : Glb2LocalMux
    port map (
            O => \N__4792\,
            I => \N__4781\
        );

    \I__1056\ : ClkMux
    port map (
            O => \N__4791\,
            I => \N__4781\
        );

    \I__1055\ : Glb2LocalMux
    port map (
            O => \N__4788\,
            I => \N__4781\
        );

    \I__1054\ : GlobalMux
    port map (
            O => \N__4781\,
            I => \CLK40\
        );

    \I__1053\ : CascadeMux
    port map (
            O => \N__4778\,
            I => \N__4775\
        );

    \I__1052\ : InMux
    port map (
            O => \N__4775\,
            I => \N__4772\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__4772\,
            I => \N__4769\
        );

    \I__1050\ : Span12Mux_h
    port map (
            O => \N__4769\,
            I => \N__4766\
        );

    \I__1049\ : Span12Mux_v
    port map (
            O => \N__4766\,
            I => \N__4763\
        );

    \I__1048\ : Odrv12
    port map (
            O => \N__4763\,
            I => \TS_CPUn_c\
        );

    \I__1047\ : InMux
    port map (
            O => \N__4760\,
            I => \N__4757\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__4757\,
            I => \U111_CYCLE_SM.TS_EN_4\
        );

    \I__1045\ : InMux
    port map (
            O => \N__4754\,
            I => \N__4745\
        );

    \I__1044\ : InMux
    port map (
            O => \N__4753\,
            I => \N__4745\
        );

    \I__1043\ : InMux
    port map (
            O => \N__4752\,
            I => \N__4745\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__4745\,
            I => \N__4741\
        );

    \I__1041\ : CascadeMux
    port map (
            O => \N__4744\,
            I => \N__4738\
        );

    \I__1040\ : Sp12to4
    port map (
            O => \N__4741\,
            I => \N__4734\
        );

    \I__1039\ : InMux
    port map (
            O => \N__4738\,
            I => \N__4731\
        );

    \I__1038\ : InMux
    port map (
            O => \N__4737\,
            I => \N__4728\
        );

    \I__1037\ : Span12Mux_h
    port map (
            O => \N__4734\,
            I => \N__4721\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__4731\,
            I => \N__4721\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__4728\,
            I => \N__4721\
        );

    \I__1034\ : Span12Mux_v
    port map (
            O => \N__4721\,
            I => \N__4718\
        );

    \I__1033\ : Odrv12
    port map (
            O => \N__4718\,
            I => \TACKn_c\
        );

    \I__1032\ : InMux
    port map (
            O => \N__4715\,
            I => \N__4709\
        );

    \I__1031\ : InMux
    port map (
            O => \N__4714\,
            I => \N__4702\
        );

    \I__1030\ : InMux
    port map (
            O => \N__4713\,
            I => \N__4702\
        );

    \I__1029\ : InMux
    port map (
            O => \N__4712\,
            I => \N__4702\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__4709\,
            I => \N__4699\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__4702\,
            I => \N__4688\
        );

    \I__1026\ : Span4Mux_v
    port map (
            O => \N__4699\,
            I => \N__4688\
        );

    \I__1025\ : InMux
    port map (
            O => \N__4698\,
            I => \N__4683\
        );

    \I__1024\ : InMux
    port map (
            O => \N__4697\,
            I => \N__4683\
        );

    \I__1023\ : InMux
    port map (
            O => \N__4696\,
            I => \N__4678\
        );

    \I__1022\ : InMux
    port map (
            O => \N__4695\,
            I => \N__4678\
        );

    \I__1021\ : InMux
    port map (
            O => \N__4694\,
            I => \N__4673\
        );

    \I__1020\ : InMux
    port map (
            O => \N__4693\,
            I => \N__4673\
        );

    \I__1019\ : Odrv4
    port map (
            O => \N__4688\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__4683\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__4678\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__4673\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1015\ : CascadeMux
    port map (
            O => \N__4664\,
            I => \N__4658\
        );

    \I__1014\ : InMux
    port map (
            O => \N__4663\,
            I => \N__4650\
        );

    \I__1013\ : InMux
    port map (
            O => \N__4662\,
            I => \N__4650\
        );

    \I__1012\ : InMux
    port map (
            O => \N__4661\,
            I => \N__4647\
        );

    \I__1011\ : InMux
    port map (
            O => \N__4658\,
            I => \N__4638\
        );

    \I__1010\ : InMux
    port map (
            O => \N__4657\,
            I => \N__4638\
        );

    \I__1009\ : InMux
    port map (
            O => \N__4656\,
            I => \N__4638\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4655\,
            I => \N__4638\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__4650\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__4647\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__4638\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1004\ : IoInMux
    port map (
            O => \N__4631\,
            I => \N__4624\
        );

    \I__1003\ : IoInMux
    port map (
            O => \N__4630\,
            I => \N__4621\
        );

    \I__1002\ : IoInMux
    port map (
            O => \N__4629\,
            I => \N__4618\
        );

    \I__1001\ : IoInMux
    port map (
            O => \N__4628\,
            I => \N__4615\
        );

    \I__1000\ : IoInMux
    port map (
            O => \N__4627\,
            I => \N__4612\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__4624\,
            I => \N__4608\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__4621\,
            I => \N__4598\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__4618\,
            I => \N__4598\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__4615\,
            I => \N__4598\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__4612\,
            I => \N__4598\
        );

    \I__994\ : IoInMux
    port map (
            O => \N__4611\,
            I => \N__4595\
        );

    \I__993\ : Span4Mux_s3_v
    port map (
            O => \N__4608\,
            I => \N__4584\
        );

    \I__992\ : InMux
    port map (
            O => \N__4607\,
            I => \N__4581\
        );

    \I__991\ : IoSpan4Mux
    port map (
            O => \N__4598\,
            I => \N__4576\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__4595\,
            I => \N__4576\
        );

    \I__989\ : IoInMux
    port map (
            O => \N__4594\,
            I => \N__4573\
        );

    \I__988\ : IoInMux
    port map (
            O => \N__4593\,
            I => \N__4570\
        );

    \I__987\ : IoInMux
    port map (
            O => \N__4592\,
            I => \N__4567\
        );

    \I__986\ : IoInMux
    port map (
            O => \N__4591\,
            I => \N__4564\
        );

    \I__985\ : IoInMux
    port map (
            O => \N__4590\,
            I => \N__4561\
        );

    \I__984\ : IoInMux
    port map (
            O => \N__4589\,
            I => \N__4558\
        );

    \I__983\ : IoInMux
    port map (
            O => \N__4588\,
            I => \N__4554\
        );

    \I__982\ : IoInMux
    port map (
            O => \N__4587\,
            I => \N__4551\
        );

    \I__981\ : Span4Mux_h
    port map (
            O => \N__4584\,
            I => \N__4542\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__4581\,
            I => \N__4539\
        );

    \I__979\ : IoSpan4Mux
    port map (
            O => \N__4576\,
            I => \N__4523\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__4573\,
            I => \N__4523\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__4570\,
            I => \N__4523\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__4567\,
            I => \N__4523\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__4564\,
            I => \N__4523\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__4561\,
            I => \N__4523\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__4558\,
            I => \N__4523\
        );

    \I__972\ : IoInMux
    port map (
            O => \N__4557\,
            I => \N__4520\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__4554\,
            I => \N__4514\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__4551\,
            I => \N__4514\
        );

    \I__969\ : IoInMux
    port map (
            O => \N__4550\,
            I => \N__4511\
        );

    \I__968\ : IoInMux
    port map (
            O => \N__4549\,
            I => \N__4508\
        );

    \I__967\ : IoInMux
    port map (
            O => \N__4548\,
            I => \N__4505\
        );

    \I__966\ : IoInMux
    port map (
            O => \N__4547\,
            I => \N__4502\
        );

    \I__965\ : IoInMux
    port map (
            O => \N__4546\,
            I => \N__4499\
        );

    \I__964\ : IoInMux
    port map (
            O => \N__4545\,
            I => \N__4496\
        );

    \I__963\ : Span4Mux_v
    port map (
            O => \N__4542\,
            I => \N__4489\
        );

    \I__962\ : Span4Mux_v
    port map (
            O => \N__4539\,
            I => \N__4486\
        );

    \I__961\ : InMux
    port map (
            O => \N__4538\,
            I => \N__4483\
        );

    \I__960\ : IoSpan4Mux
    port map (
            O => \N__4523\,
            I => \N__4477\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4520\,
            I => \N__4477\
        );

    \I__958\ : IoInMux
    port map (
            O => \N__4519\,
            I => \N__4474\
        );

    \I__957\ : IoSpan4Mux
    port map (
            O => \N__4514\,
            I => \N__4458\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__4511\,
            I => \N__4458\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__4508\,
            I => \N__4458\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__4505\,
            I => \N__4458\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__4502\,
            I => \N__4458\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__4499\,
            I => \N__4458\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__4496\,
            I => \N__4458\
        );

    \I__950\ : IoInMux
    port map (
            O => \N__4495\,
            I => \N__4455\
        );

    \I__949\ : IoInMux
    port map (
            O => \N__4494\,
            I => \N__4452\
        );

    \I__948\ : IoInMux
    port map (
            O => \N__4493\,
            I => \N__4449\
        );

    \I__947\ : IoInMux
    port map (
            O => \N__4492\,
            I => \N__4446\
        );

    \I__946\ : Span4Mux_v
    port map (
            O => \N__4489\,
            I => \N__4439\
        );

    \I__945\ : Span4Mux_v
    port map (
            O => \N__4486\,
            I => \N__4439\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4483\,
            I => \N__4436\
        );

    \I__943\ : IoInMux
    port map (
            O => \N__4482\,
            I => \N__4433\
        );

    \I__942\ : IoSpan4Mux
    port map (
            O => \N__4477\,
            I => \N__4428\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__4474\,
            I => \N__4428\
        );

    \I__940\ : IoInMux
    port map (
            O => \N__4473\,
            I => \N__4425\
        );

    \I__939\ : IoSpan4Mux
    port map (
            O => \N__4458\,
            I => \N__4414\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4455\,
            I => \N__4414\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__4452\,
            I => \N__4414\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__4449\,
            I => \N__4414\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__4446\,
            I => \N__4414\
        );

    \I__934\ : IoInMux
    port map (
            O => \N__4445\,
            I => \N__4410\
        );

    \I__933\ : IoInMux
    port map (
            O => \N__4444\,
            I => \N__4407\
        );

    \I__932\ : Sp12to4
    port map (
            O => \N__4439\,
            I => \N__4402\
        );

    \I__931\ : Span12Mux_v
    port map (
            O => \N__4436\,
            I => \N__4399\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__4433\,
            I => \N__4396\
        );

    \I__929\ : IoSpan4Mux
    port map (
            O => \N__4428\,
            I => \N__4391\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__4425\,
            I => \N__4391\
        );

    \I__927\ : IoSpan4Mux
    port map (
            O => \N__4414\,
            I => \N__4388\
        );

    \I__926\ : IoInMux
    port map (
            O => \N__4413\,
            I => \N__4385\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__4410\,
            I => \N__4380\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__4407\,
            I => \N__4380\
        );

    \I__923\ : IoInMux
    port map (
            O => \N__4406\,
            I => \N__4377\
        );

    \I__922\ : IoInMux
    port map (
            O => \N__4405\,
            I => \N__4374\
        );

    \I__921\ : Span12Mux_h
    port map (
            O => \N__4402\,
            I => \N__4371\
        );

    \I__920\ : Span12Mux_h
    port map (
            O => \N__4399\,
            I => \N__4366\
        );

    \I__919\ : Span12Mux_s11_v
    port map (
            O => \N__4396\,
            I => \N__4366\
        );

    \I__918\ : IoSpan4Mux
    port map (
            O => \N__4391\,
            I => \N__4363\
        );

    \I__917\ : IoSpan4Mux
    port map (
            O => \N__4388\,
            I => \N__4358\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__4385\,
            I => \N__4358\
        );

    \I__915\ : IoSpan4Mux
    port map (
            O => \N__4380\,
            I => \N__4353\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__4377\,
            I => \N__4353\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__4374\,
            I => \N__4350\
        );

    \I__912\ : Odrv12
    port map (
            O => \N__4371\,
            I => \RnW_c\
        );

    \I__911\ : Odrv12
    port map (
            O => \N__4366\,
            I => \RnW_c\
        );

    \I__910\ : Odrv4
    port map (
            O => \N__4363\,
            I => \RnW_c\
        );

    \I__909\ : Odrv4
    port map (
            O => \N__4358\,
            I => \RnW_c\
        );

    \I__908\ : Odrv4
    port map (
            O => \N__4353\,
            I => \RnW_c\
        );

    \I__907\ : Odrv12
    port map (
            O => \N__4350\,
            I => \RnW_c\
        );

    \I__906\ : CascadeMux
    port map (
            O => \N__4337\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_\
        );

    \I__905\ : CascadeMux
    port map (
            O => \N__4334\,
            I => \N__4328\
        );

    \I__904\ : CascadeMux
    port map (
            O => \N__4333\,
            I => \N__4324\
        );

    \I__903\ : CascadeMux
    port map (
            O => \N__4332\,
            I => \N__4317\
        );

    \I__902\ : InMux
    port map (
            O => \N__4331\,
            I => \N__4314\
        );

    \I__901\ : InMux
    port map (
            O => \N__4328\,
            I => \N__4309\
        );

    \I__900\ : InMux
    port map (
            O => \N__4327\,
            I => \N__4309\
        );

    \I__899\ : InMux
    port map (
            O => \N__4324\,
            I => \N__4306\
        );

    \I__898\ : InMux
    port map (
            O => \N__4323\,
            I => \N__4301\
        );

    \I__897\ : InMux
    port map (
            O => \N__4322\,
            I => \N__4301\
        );

    \I__896\ : InMux
    port map (
            O => \N__4321\,
            I => \N__4294\
        );

    \I__895\ : InMux
    port map (
            O => \N__4320\,
            I => \N__4294\
        );

    \I__894\ : InMux
    port map (
            O => \N__4317\,
            I => \N__4294\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__4314\,
            I => \N__4291\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__4309\,
            I => \N__4284\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__4306\,
            I => \N__4284\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__4301\,
            I => \N__4284\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__4294\,
            I => \N__4281\
        );

    \I__888\ : Span4Mux_v
    port map (
            O => \N__4291\,
            I => \N__4276\
        );

    \I__887\ : Span4Mux_v
    port map (
            O => \N__4284\,
            I => \N__4276\
        );

    \I__886\ : Span4Mux_v
    port map (
            O => \N__4281\,
            I => \N__4273\
        );

    \I__885\ : Span4Mux_v
    port map (
            O => \N__4276\,
            I => \N__4270\
        );

    \I__884\ : Span4Mux_h
    port map (
            O => \N__4273\,
            I => \N__4267\
        );

    \I__883\ : Span4Mux_v
    port map (
            O => \N__4270\,
            I => \N__4264\
        );

    \I__882\ : Span4Mux_h
    port map (
            O => \N__4267\,
            I => \N__4261\
        );

    \I__881\ : Span4Mux_v
    port map (
            O => \N__4264\,
            I => \N__4258\
        );

    \I__880\ : Sp12to4
    port map (
            O => \N__4261\,
            I => \N__4255\
        );

    \I__879\ : Sp12to4
    port map (
            O => \N__4258\,
            I => \N__4252\
        );

    \I__878\ : Span12Mux_v
    port map (
            O => \N__4255\,
            I => \N__4247\
        );

    \I__877\ : Span12Mux_h
    port map (
            O => \N__4252\,
            I => \N__4247\
        );

    \I__876\ : Odrv12
    port map (
            O => \N__4247\,
            I => \RESETn_c\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__4244\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0_cascade_\
        );

    \I__874\ : InMux
    port map (
            O => \N__4241\,
            I => \N__4238\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__4238\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa\
        );

    \I__872\ : InMux
    port map (
            O => \N__4235\,
            I => \N__4232\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__4232\,
            I => \N__4229\
        );

    \I__870\ : Span12Mux_v
    port map (
            O => \N__4229\,
            I => \N__4226\
        );

    \I__869\ : Span12Mux_h
    port map (
            O => \N__4226\,
            I => \N__4223\
        );

    \I__868\ : Odrv12
    port map (
            O => \N__4223\,
            I => \D_LM_AMIGA_in_7\
        );

    \I__867\ : IoInMux
    port map (
            O => \N__4220\,
            I => \N__4217\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__4217\,
            I => \N__4214\
        );

    \I__865\ : IoSpan4Mux
    port map (
            O => \N__4214\,
            I => \N__4211\
        );

    \I__864\ : Span4Mux_s3_h
    port map (
            O => \N__4211\,
            I => \N__4208\
        );

    \I__863\ : Sp12to4
    port map (
            O => \N__4208\,
            I => \N__4205\
        );

    \I__862\ : Span12Mux_s11_h
    port map (
            O => \N__4205\,
            I => \N__4202\
        );

    \I__861\ : Odrv12
    port map (
            O => \N__4202\,
            I => \un1_D_LM_AMIGA_7\
        );

    \I__860\ : InMux
    port map (
            O => \N__4199\,
            I => \N__4196\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__4196\,
            I => \N__4193\
        );

    \I__858\ : Odrv4
    port map (
            O => \N__4193\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\
        );

    \I__857\ : InMux
    port map (
            O => \N__4190\,
            I => \N__4187\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__4187\,
            I => \N__4184\
        );

    \I__855\ : Span4Mux_v
    port map (
            O => \N__4184\,
            I => \N__4181\
        );

    \I__854\ : Span4Mux_v
    port map (
            O => \N__4181\,
            I => \N__4177\
        );

    \I__853\ : InMux
    port map (
            O => \N__4180\,
            I => \N__4174\
        );

    \I__852\ : Span4Mux_v
    port map (
            O => \N__4177\,
            I => \N__4168\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__4174\,
            I => \N__4168\
        );

    \I__850\ : InMux
    port map (
            O => \N__4173\,
            I => \N__4165\
        );

    \I__849\ : Span4Mux_h
    port map (
            O => \N__4168\,
            I => \N__4160\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__4165\,
            I => \N__4160\
        );

    \I__847\ : Span4Mux_v
    port map (
            O => \N__4160\,
            I => \N__4157\
        );

    \I__846\ : Span4Mux_v
    port map (
            O => \N__4157\,
            I => \N__4154\
        );

    \I__845\ : Sp12to4
    port map (
            O => \N__4154\,
            I => \N__4151\
        );

    \I__844\ : Span12Mux_h
    port map (
            O => \N__4151\,
            I => \N__4148\
        );

    \I__843\ : Odrv12
    port map (
            O => \N__4148\,
            I => \D_UM_AMIGA_in_4\
        );

    \I__842\ : IoInMux
    port map (
            O => \N__4145\,
            I => \N__4142\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__4142\,
            I => \N__4139\
        );

    \I__840\ : Span4Mux_s3_v
    port map (
            O => \N__4139\,
            I => \N__4136\
        );

    \I__839\ : Span4Mux_h
    port map (
            O => \N__4136\,
            I => \N__4133\
        );

    \I__838\ : Sp12to4
    port map (
            O => \N__4133\,
            I => \N__4130\
        );

    \I__837\ : Span12Mux_h
    port map (
            O => \N__4130\,
            I => \N__4127\
        );

    \I__836\ : Odrv12
    port map (
            O => \N__4127\,
            I => \un1_D_UM_AMIGA_4\
        );

    \I__835\ : IoInMux
    port map (
            O => \N__4124\,
            I => \N__4121\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__4121\,
            I => \N__4118\
        );

    \I__833\ : IoSpan4Mux
    port map (
            O => \N__4118\,
            I => \N__4115\
        );

    \I__832\ : Span4Mux_s3_h
    port map (
            O => \N__4115\,
            I => \N__4111\
        );

    \I__831\ : InMux
    port map (
            O => \N__4114\,
            I => \N__4108\
        );

    \I__830\ : Sp12to4
    port map (
            O => \N__4111\,
            I => \N__4105\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__4108\,
            I => \N__4102\
        );

    \I__828\ : Span12Mux_v
    port map (
            O => \N__4105\,
            I => \N__4099\
        );

    \I__827\ : Span12Mux_v
    port map (
            O => \N__4102\,
            I => \N__4096\
        );

    \I__826\ : Span12Mux_h
    port map (
            O => \N__4099\,
            I => \N__4091\
        );

    \I__825\ : Span12Mux_v
    port map (
            O => \N__4096\,
            I => \N__4091\
        );

    \I__824\ : Span12Mux_h
    port map (
            O => \N__4091\,
            I => \N__4088\
        );

    \I__823\ : Odrv12
    port map (
            O => \N__4088\,
            I => \D_LL_040_in_5\
        );

    \I__822\ : InMux
    port map (
            O => \N__4085\,
            I => \N__4082\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4082\,
            I => \N__4079\
        );

    \I__820\ : Span4Mux_v
    port map (
            O => \N__4079\,
            I => \N__4076\
        );

    \I__819\ : Sp12to4
    port map (
            O => \N__4076\,
            I => \N__4073\
        );

    \I__818\ : Span12Mux_h
    port map (
            O => \N__4073\,
            I => \N__4070\
        );

    \I__817\ : Odrv12
    port map (
            O => \N__4070\,
            I => \D_UM_040_in_5\
        );

    \I__816\ : InMux
    port map (
            O => \N__4067\,
            I => \N__4064\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__4064\,
            I => \N__4061\
        );

    \I__814\ : Sp12to4
    port map (
            O => \N__4061\,
            I => \N__4058\
        );

    \I__813\ : Span12Mux_v
    port map (
            O => \N__4058\,
            I => \N__4055\
        );

    \I__812\ : Span12Mux_h
    port map (
            O => \N__4055\,
            I => \N__4052\
        );

    \I__811\ : Odrv12
    port map (
            O => \N__4052\,
            I => \D_UU_040_in_0\
        );

    \I__810\ : IoInMux
    port map (
            O => \N__4049\,
            I => \N__4046\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__4046\,
            I => \N__4042\
        );

    \I__808\ : InMux
    port map (
            O => \N__4045\,
            I => \N__4039\
        );

    \I__807\ : IoSpan4Mux
    port map (
            O => \N__4042\,
            I => \N__4036\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__4039\,
            I => \N__4033\
        );

    \I__805\ : IoSpan4Mux
    port map (
            O => \N__4036\,
            I => \N__4030\
        );

    \I__804\ : Span4Mux_v
    port map (
            O => \N__4033\,
            I => \N__4027\
        );

    \I__803\ : Span4Mux_s2_h
    port map (
            O => \N__4030\,
            I => \N__4024\
        );

    \I__802\ : Sp12to4
    port map (
            O => \N__4027\,
            I => \N__4021\
        );

    \I__801\ : Sp12to4
    port map (
            O => \N__4024\,
            I => \N__4018\
        );

    \I__800\ : Span12Mux_h
    port map (
            O => \N__4021\,
            I => \N__4015\
        );

    \I__799\ : Span12Mux_h
    port map (
            O => \N__4018\,
            I => \N__4012\
        );

    \I__798\ : Span12Mux_v
    port map (
            O => \N__4015\,
            I => \N__4009\
        );

    \I__797\ : Span12Mux_h
    port map (
            O => \N__4012\,
            I => \N__4004\
        );

    \I__796\ : Span12Mux_v
    port map (
            O => \N__4009\,
            I => \N__4004\
        );

    \I__795\ : Odrv12
    port map (
            O => \N__4004\,
            I => \D_LM_040_in_0\
        );

    \I__794\ : IoInMux
    port map (
            O => \N__4001\,
            I => \N__3998\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__3998\,
            I => \N__3995\
        );

    \I__792\ : IoSpan4Mux
    port map (
            O => \N__3995\,
            I => \N__3992\
        );

    \I__791\ : Sp12to4
    port map (
            O => \N__3992\,
            I => \N__3989\
        );

    \I__790\ : Span12Mux_s6_v
    port map (
            O => \N__3989\,
            I => \N__3986\
        );

    \I__789\ : Odrv12
    port map (
            O => \N__3986\,
            I => \un1_D_UU_040_0\
        );

    \I__788\ : InMux
    port map (
            O => \N__3983\,
            I => \N__3980\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__3980\,
            I => \N__3977\
        );

    \I__786\ : Odrv12
    port map (
            O => \N__3977\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\
        );

    \I__785\ : InMux
    port map (
            O => \N__3974\,
            I => \N__3970\
        );

    \I__784\ : InMux
    port map (
            O => \N__3973\,
            I => \N__3967\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__3970\,
            I => \N__3962\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__3967\,
            I => \N__3962\
        );

    \I__781\ : Span4Mux_v
    port map (
            O => \N__3962\,
            I => \N__3958\
        );

    \I__780\ : InMux
    port map (
            O => \N__3961\,
            I => \N__3955\
        );

    \I__779\ : Span4Mux_v
    port map (
            O => \N__3958\,
            I => \N__3950\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__3955\,
            I => \N__3950\
        );

    \I__777\ : Span4Mux_v
    port map (
            O => \N__3950\,
            I => \N__3947\
        );

    \I__776\ : IoSpan4Mux
    port map (
            O => \N__3947\,
            I => \N__3944\
        );

    \I__775\ : IoSpan4Mux
    port map (
            O => \N__3944\,
            I => \N__3941\
        );

    \I__774\ : Odrv4
    port map (
            O => \N__3941\,
            I => \D_UU_AMIGA_in_4\
        );

    \I__773\ : IoInMux
    port map (
            O => \N__3938\,
            I => \N__3935\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__3935\,
            I => \N__3932\
        );

    \I__771\ : Span4Mux_s2_v
    port map (
            O => \N__3932\,
            I => \N__3929\
        );

    \I__770\ : Span4Mux_v
    port map (
            O => \N__3929\,
            I => \N__3926\
        );

    \I__769\ : Sp12to4
    port map (
            O => \N__3926\,
            I => \N__3923\
        );

    \I__768\ : Odrv12
    port map (
            O => \N__3923\,
            I => \un1_D_UU_AMIGA_4\
        );

    \I__767\ : IoInMux
    port map (
            O => \N__3920\,
            I => \N__3917\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__3917\,
            I => \N__3913\
        );

    \I__765\ : InMux
    port map (
            O => \N__3916\,
            I => \N__3910\
        );

    \I__764\ : IoSpan4Mux
    port map (
            O => \N__3913\,
            I => \N__3907\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__3910\,
            I => \N__3904\
        );

    \I__762\ : Span4Mux_s2_h
    port map (
            O => \N__3907\,
            I => \N__3901\
        );

    \I__761\ : Span4Mux_v
    port map (
            O => \N__3904\,
            I => \N__3898\
        );

    \I__760\ : Sp12to4
    port map (
            O => \N__3901\,
            I => \N__3895\
        );

    \I__759\ : Sp12to4
    port map (
            O => \N__3898\,
            I => \N__3892\
        );

    \I__758\ : Span12Mux_h
    port map (
            O => \N__3895\,
            I => \N__3889\
        );

    \I__757\ : Span12Mux_h
    port map (
            O => \N__3892\,
            I => \N__3886\
        );

    \I__756\ : Span12Mux_h
    port map (
            O => \N__3889\,
            I => \N__3883\
        );

    \I__755\ : Span12Mux_v
    port map (
            O => \N__3886\,
            I => \N__3880\
        );

    \I__754\ : Odrv12
    port map (
            O => \N__3883\,
            I => \D_LL_040_in_0\
        );

    \I__753\ : Odrv12
    port map (
            O => \N__3880\,
            I => \D_LL_040_in_0\
        );

    \I__752\ : InMux
    port map (
            O => \N__3875\,
            I => \N__3872\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__3872\,
            I => \N__3869\
        );

    \I__750\ : Span12Mux_h
    port map (
            O => \N__3869\,
            I => \N__3866\
        );

    \I__749\ : Odrv12
    port map (
            O => \N__3866\,
            I => \D_UM_040_in_0\
        );

    \I__748\ : IoInMux
    port map (
            O => \N__3863\,
            I => \N__3860\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__3860\,
            I => \N__3857\
        );

    \I__746\ : Span4Mux_s3_h
    port map (
            O => \N__3857\,
            I => \N__3854\
        );

    \I__745\ : Span4Mux_h
    port map (
            O => \N__3854\,
            I => \N__3851\
        );

    \I__744\ : Span4Mux_h
    port map (
            O => \N__3851\,
            I => \N__3848\
        );

    \I__743\ : Span4Mux_h
    port map (
            O => \N__3848\,
            I => \N__3845\
        );

    \I__742\ : Odrv4
    port map (
            O => \N__3845\,
            I => \un1_D_UM_040_0\
        );

    \I__741\ : IoInMux
    port map (
            O => \N__3842\,
            I => \N__3837\
        );

    \I__740\ : IoInMux
    port map (
            O => \N__3841\,
            I => \N__3834\
        );

    \I__739\ : IoInMux
    port map (
            O => \N__3840\,
            I => \N__3831\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__3837\,
            I => \N__3828\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__3834\,
            I => \N__3825\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__3831\,
            I => \N__3822\
        );

    \I__735\ : Span12Mux_s4_h
    port map (
            O => \N__3828\,
            I => \N__3819\
        );

    \I__734\ : Span12Mux_s7_v
    port map (
            O => \N__3825\,
            I => \N__3816\
        );

    \I__733\ : Span12Mux_s7_h
    port map (
            O => \N__3822\,
            I => \N__3813\
        );

    \I__732\ : Odrv12
    port map (
            O => \N__3819\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__731\ : Odrv12
    port map (
            O => \N__3816\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__730\ : Odrv12
    port map (
            O => \N__3813\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__729\ : IoInMux
    port map (
            O => \N__3806\,
            I => \N__3803\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__3803\,
            I => \N__3800\
        );

    \I__727\ : Span4Mux_s3_h
    port map (
            O => \N__3800\,
            I => \N__3797\
        );

    \I__726\ : Span4Mux_h
    port map (
            O => \N__3797\,
            I => \N__3794\
        );

    \I__725\ : Span4Mux_h
    port map (
            O => \N__3794\,
            I => \N__3791\
        );

    \I__724\ : Span4Mux_h
    port map (
            O => \N__3791\,
            I => \N__3788\
        );

    \I__723\ : Odrv4
    port map (
            O => \N__3788\,
            I => \un1_D_UM_AMIGA_0\
        );

    \I__722\ : InMux
    port map (
            O => \N__3785\,
            I => \N__3782\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__3782\,
            I => \N__3779\
        );

    \I__720\ : Span4Mux_v
    port map (
            O => \N__3779\,
            I => \N__3775\
        );

    \I__719\ : InMux
    port map (
            O => \N__3778\,
            I => \N__3772\
        );

    \I__718\ : Span4Mux_v
    port map (
            O => \N__3775\,
            I => \N__3769\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__3772\,
            I => \N__3766\
        );

    \I__716\ : Span4Mux_v
    port map (
            O => \N__3769\,
            I => \N__3760\
        );

    \I__715\ : Span4Mux_v
    port map (
            O => \N__3766\,
            I => \N__3760\
        );

    \I__714\ : InMux
    port map (
            O => \N__3765\,
            I => \N__3757\
        );

    \I__713\ : Sp12to4
    port map (
            O => \N__3760\,
            I => \N__3752\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__3757\,
            I => \N__3752\
        );

    \I__711\ : Span12Mux_h
    port map (
            O => \N__3752\,
            I => \N__3749\
        );

    \I__710\ : Odrv12
    port map (
            O => \N__3749\,
            I => \D_UM_AMIGA_in_0\
        );

    \I__709\ : InMux
    port map (
            O => \N__3746\,
            I => \N__3743\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__3743\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\
        );

    \I__707\ : InMux
    port map (
            O => \N__3740\,
            I => \N__3737\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__3737\,
            I => \N__3734\
        );

    \I__705\ : Span4Mux_v
    port map (
            O => \N__3734\,
            I => \N__3731\
        );

    \I__704\ : Sp12to4
    port map (
            O => \N__3731\,
            I => \N__3728\
        );

    \I__703\ : Span12Mux_h
    port map (
            O => \N__3728\,
            I => \N__3725\
        );

    \I__702\ : Odrv12
    port map (
            O => \N__3725\,
            I => \D_LM_AMIGA_in_4\
        );

    \I__701\ : IoInMux
    port map (
            O => \N__3722\,
            I => \N__3719\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__3719\,
            I => \N__3716\
        );

    \I__699\ : IoSpan4Mux
    port map (
            O => \N__3716\,
            I => \N__3713\
        );

    \I__698\ : IoSpan4Mux
    port map (
            O => \N__3713\,
            I => \N__3710\
        );

    \I__697\ : Span4Mux_s0_h
    port map (
            O => \N__3710\,
            I => \N__3707\
        );

    \I__696\ : Sp12to4
    port map (
            O => \N__3707\,
            I => \N__3704\
        );

    \I__695\ : Span12Mux_s9_h
    port map (
            O => \N__3704\,
            I => \N__3701\
        );

    \I__694\ : Odrv12
    port map (
            O => \N__3701\,
            I => \un1_D_LM_AMIGA_4\
        );

    \I__693\ : CascadeMux
    port map (
            O => \N__3698\,
            I => \U111_CYCLE_SM.TS_EN10_cascade_\
        );

    \I__692\ : InMux
    port map (
            O => \N__3695\,
            I => \N__3691\
        );

    \I__691\ : InMux
    port map (
            O => \N__3694\,
            I => \N__3688\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__3691\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__3688\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__688\ : CascadeMux
    port map (
            O => \N__3683\,
            I => \U111_CYCLE_SM.LW_CYCLE_r_1_cascade_\
        );

    \I__687\ : IoInMux
    port map (
            O => \N__3680\,
            I => \N__3677\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__3677\,
            I => \N__3674\
        );

    \I__685\ : IoSpan4Mux
    port map (
            O => \N__3674\,
            I => \N__3671\
        );

    \I__684\ : Span4Mux_s0_v
    port map (
            O => \N__3671\,
            I => \N__3668\
        );

    \I__683\ : Sp12to4
    port map (
            O => \N__3668\,
            I => \N__3665\
        );

    \I__682\ : Span12Mux_v
    port map (
            O => \N__3665\,
            I => \N__3661\
        );

    \I__681\ : InMux
    port map (
            O => \N__3664\,
            I => \N__3658\
        );

    \I__680\ : Odrv12
    port map (
            O => \N__3661\,
            I => \TSn_c\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__3658\,
            I => \TSn_c\
        );

    \I__678\ : CascadeMux
    port map (
            O => \N__3653\,
            I => \N__3649\
        );

    \I__677\ : InMux
    port map (
            O => \N__3652\,
            I => \N__3646\
        );

    \I__676\ : InMux
    port map (
            O => \N__3649\,
            I => \N__3643\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__3646\,
            I => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3643\,
            I => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\
        );

    \I__673\ : InMux
    port map (
            O => \N__3638\,
            I => \N__3635\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__3635\,
            I => \N__3632\
        );

    \I__671\ : Odrv12
    port map (
            O => \N__3632\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\
        );

    \I__670\ : InMux
    port map (
            O => \N__3629\,
            I => \N__3625\
        );

    \I__669\ : InMux
    port map (
            O => \N__3628\,
            I => \N__3622\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__3625\,
            I => \N__3618\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__3622\,
            I => \N__3615\
        );

    \I__666\ : InMux
    port map (
            O => \N__3621\,
            I => \N__3612\
        );

    \I__665\ : Span4Mux_v
    port map (
            O => \N__3618\,
            I => \N__3609\
        );

    \I__664\ : Span4Mux_v
    port map (
            O => \N__3615\,
            I => \N__3604\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__3612\,
            I => \N__3604\
        );

    \I__662\ : Span4Mux_v
    port map (
            O => \N__3609\,
            I => \N__3599\
        );

    \I__661\ : Span4Mux_v
    port map (
            O => \N__3604\,
            I => \N__3599\
        );

    \I__660\ : Sp12to4
    port map (
            O => \N__3599\,
            I => \N__3596\
        );

    \I__659\ : Span12Mux_h
    port map (
            O => \N__3596\,
            I => \N__3593\
        );

    \I__658\ : Odrv12
    port map (
            O => \N__3593\,
            I => \D_UU_AMIGA_in_6\
        );

    \I__657\ : IoInMux
    port map (
            O => \N__3590\,
            I => \N__3587\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__3587\,
            I => \N__3584\
        );

    \I__655\ : IoSpan4Mux
    port map (
            O => \N__3584\,
            I => \N__3581\
        );

    \I__654\ : IoSpan4Mux
    port map (
            O => \N__3581\,
            I => \N__3578\
        );

    \I__653\ : Sp12to4
    port map (
            O => \N__3578\,
            I => \N__3575\
        );

    \I__652\ : Span12Mux_s6_v
    port map (
            O => \N__3575\,
            I => \N__3572\
        );

    \I__651\ : Odrv12
    port map (
            O => \N__3572\,
            I => \un1_D_UU_AMIGA_6\
        );

    \I__650\ : InMux
    port map (
            O => \N__3569\,
            I => \N__3566\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__3566\,
            I => \N__3563\
        );

    \I__648\ : Span4Mux_v
    port map (
            O => \N__3563\,
            I => \N__3560\
        );

    \I__647\ : Span4Mux_h
    port map (
            O => \N__3560\,
            I => \N__3557\
        );

    \I__646\ : Sp12to4
    port map (
            O => \N__3557\,
            I => \N__3554\
        );

    \I__645\ : Span12Mux_h
    port map (
            O => \N__3554\,
            I => \N__3551\
        );

    \I__644\ : Odrv12
    port map (
            O => \N__3551\,
            I => \D_UM_040_in_4\
        );

    \I__643\ : IoInMux
    port map (
            O => \N__3548\,
            I => \N__3545\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__3545\,
            I => \N__3541\
        );

    \I__641\ : InMux
    port map (
            O => \N__3544\,
            I => \N__3538\
        );

    \I__640\ : Span4Mux_s2_h
    port map (
            O => \N__3541\,
            I => \N__3535\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__3538\,
            I => \N__3532\
        );

    \I__638\ : Span4Mux_v
    port map (
            O => \N__3535\,
            I => \N__3529\
        );

    \I__637\ : Span12Mux_v
    port map (
            O => \N__3532\,
            I => \N__3526\
        );

    \I__636\ : Sp12to4
    port map (
            O => \N__3529\,
            I => \N__3523\
        );

    \I__635\ : Span12Mux_v
    port map (
            O => \N__3526\,
            I => \N__3518\
        );

    \I__634\ : Span12Mux_h
    port map (
            O => \N__3523\,
            I => \N__3518\
        );

    \I__633\ : Span12Mux_h
    port map (
            O => \N__3518\,
            I => \N__3515\
        );

    \I__632\ : Odrv12
    port map (
            O => \N__3515\,
            I => \D_LL_040_in_4\
        );

    \I__631\ : IoInMux
    port map (
            O => \N__3512\,
            I => \N__3509\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__3509\,
            I => \N__3506\
        );

    \I__629\ : Span4Mux_s1_h
    port map (
            O => \N__3506\,
            I => \N__3503\
        );

    \I__628\ : Span4Mux_h
    port map (
            O => \N__3503\,
            I => \N__3500\
        );

    \I__627\ : Span4Mux_h
    port map (
            O => \N__3500\,
            I => \N__3497\
        );

    \I__626\ : Span4Mux_h
    port map (
            O => \N__3497\,
            I => \N__3494\
        );

    \I__625\ : Odrv4
    port map (
            O => \N__3494\,
            I => \un1_D_UM_040_4\
        );

    \I__624\ : InMux
    port map (
            O => \N__3491\,
            I => \N__3488\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3488\,
            I => \N__3485\
        );

    \I__622\ : Span4Mux_v
    port map (
            O => \N__3485\,
            I => \N__3482\
        );

    \I__621\ : Sp12to4
    port map (
            O => \N__3482\,
            I => \N__3479\
        );

    \I__620\ : Span12Mux_h
    port map (
            O => \N__3479\,
            I => \N__3476\
        );

    \I__619\ : Odrv12
    port map (
            O => \N__3476\,
            I => \D_LL_AMIGA_in_1\
        );

    \I__618\ : IoInMux
    port map (
            O => \N__3473\,
            I => \N__3470\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__3470\,
            I => \N__3467\
        );

    \I__616\ : IoSpan4Mux
    port map (
            O => \N__3467\,
            I => \N__3464\
        );

    \I__615\ : Span4Mux_s3_h
    port map (
            O => \N__3464\,
            I => \N__3461\
        );

    \I__614\ : Sp12to4
    port map (
            O => \N__3461\,
            I => \N__3458\
        );

    \I__613\ : Span12Mux_h
    port map (
            O => \N__3458\,
            I => \N__3455\
        );

    \I__612\ : Odrv12
    port map (
            O => \N__3455\,
            I => \un1_D_LL_AMIGA_1\
        );

    \I__611\ : InMux
    port map (
            O => \N__3452\,
            I => \N__3449\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__3449\,
            I => \N__3446\
        );

    \I__609\ : Span12Mux_h
    port map (
            O => \N__3446\,
            I => \N__3442\
        );

    \I__608\ : InMux
    port map (
            O => \N__3445\,
            I => \N__3439\
        );

    \I__607\ : Odrv12
    port map (
            O => \N__3442\,
            I => \U111_CYCLE_SM.A_OUTZ0\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__3439\,
            I => \U111_CYCLE_SM.A_OUTZ0\
        );

    \I__605\ : InMux
    port map (
            O => \N__3434\,
            I => \N__3431\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__3431\,
            I => \U111_CYCLE_SM.un1_CYCLE_STATE_1_0\
        );

    \I__603\ : CascadeMux
    port map (
            O => \N__3428\,
            I => \U111_CYCLE_SM.un1_CYCLE_STATE_1_0_cascade_\
        );

    \I__602\ : InMux
    port map (
            O => \N__3425\,
            I => \N__3421\
        );

    \I__601\ : SRMux
    port map (
            O => \N__3424\,
            I => \N__3418\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__3421\,
            I => \RESETn_c_i\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__3418\,
            I => \RESETn_c_i\
        );

    \I__598\ : CEMux
    port map (
            O => \N__3413\,
            I => \N__3410\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__3410\,
            I => \N__3407\
        );

    \I__596\ : Odrv12
    port map (
            O => \N__3407\,
            I => \U111_CYCLE_SM.un1_CYCLE_STATE_1_0_0\
        );

    \I__595\ : InMux
    port map (
            O => \N__3404\,
            I => \N__3401\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__3401\,
            I => \U111_CYCLE_SM.TA_ENZ0\
        );

    \I__593\ : IoInMux
    port map (
            O => \N__3398\,
            I => \N__3395\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__3395\,
            I => \N__3392\
        );

    \I__591\ : Span4Mux_s2_v
    port map (
            O => \N__3392\,
            I => \N__3389\
        );

    \I__590\ : Sp12to4
    port map (
            O => \N__3389\,
            I => \N__3386\
        );

    \I__589\ : Span12Mux_h
    port map (
            O => \N__3386\,
            I => \N__3383\
        );

    \I__588\ : Span12Mux_v
    port map (
            O => \N__3383\,
            I => \N__3380\
        );

    \I__587\ : Odrv12
    port map (
            O => \N__3380\,
            I => \TAn_0_i\
        );

    \I__586\ : InMux
    port map (
            O => \N__3377\,
            I => \N__3374\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__3374\,
            I => \N__3371\
        );

    \I__584\ : Span12Mux_h
    port map (
            O => \N__3371\,
            I => \N__3368\
        );

    \I__583\ : Odrv12
    port map (
            O => \N__3368\,
            I => \D_LM_AMIGA_in_2\
        );

    \I__582\ : IoInMux
    port map (
            O => \N__3365\,
            I => \N__3362\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__3362\,
            I => \N__3359\
        );

    \I__580\ : Span12Mux_s8_h
    port map (
            O => \N__3359\,
            I => \N__3356\
        );

    \I__579\ : Span12Mux_h
    port map (
            O => \N__3356\,
            I => \N__3353\
        );

    \I__578\ : Odrv12
    port map (
            O => \N__3353\,
            I => \un1_D_LM_AMIGA_2\
        );

    \I__577\ : IoInMux
    port map (
            O => \N__3350\,
            I => \N__3347\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__3347\,
            I => \N__3344\
        );

    \I__575\ : IoSpan4Mux
    port map (
            O => \N__3344\,
            I => \N__3340\
        );

    \I__574\ : InMux
    port map (
            O => \N__3343\,
            I => \N__3337\
        );

    \I__573\ : Span4Mux_s2_h
    port map (
            O => \N__3340\,
            I => \N__3334\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__3337\,
            I => \N__3331\
        );

    \I__571\ : Sp12to4
    port map (
            O => \N__3334\,
            I => \N__3328\
        );

    \I__570\ : Span4Mux_v
    port map (
            O => \N__3331\,
            I => \N__3325\
        );

    \I__569\ : Span12Mux_h
    port map (
            O => \N__3328\,
            I => \N__3320\
        );

    \I__568\ : Sp12to4
    port map (
            O => \N__3325\,
            I => \N__3320\
        );

    \I__567\ : Span12Mux_h
    port map (
            O => \N__3320\,
            I => \N__3317\
        );

    \I__566\ : Odrv12
    port map (
            O => \N__3317\,
            I => \D_LM_040_in_7\
        );

    \I__565\ : InMux
    port map (
            O => \N__3314\,
            I => \N__3311\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__3311\,
            I => \N__3308\
        );

    \I__563\ : Span4Mux_v
    port map (
            O => \N__3308\,
            I => \N__3305\
        );

    \I__562\ : Span4Mux_h
    port map (
            O => \N__3305\,
            I => \N__3302\
        );

    \I__561\ : Sp12to4
    port map (
            O => \N__3302\,
            I => \N__3299\
        );

    \I__560\ : Span12Mux_h
    port map (
            O => \N__3299\,
            I => \N__3296\
        );

    \I__559\ : Odrv12
    port map (
            O => \N__3296\,
            I => \D_UU_040_in_7\
        );

    \I__558\ : IoInMux
    port map (
            O => \N__3293\,
            I => \N__3290\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__3290\,
            I => \N__3287\
        );

    \I__556\ : Span4Mux_s3_v
    port map (
            O => \N__3287\,
            I => \N__3284\
        );

    \I__555\ : Span4Mux_h
    port map (
            O => \N__3284\,
            I => \N__3281\
        );

    \I__554\ : Span4Mux_h
    port map (
            O => \N__3281\,
            I => \N__3278\
        );

    \I__553\ : Odrv4
    port map (
            O => \N__3278\,
            I => \un1_D_UU_040_7\
        );

    \I__552\ : InMux
    port map (
            O => \N__3275\,
            I => \N__3272\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3272\,
            I => \N__3269\
        );

    \I__550\ : Span4Mux_v
    port map (
            O => \N__3269\,
            I => \N__3266\
        );

    \I__549\ : Sp12to4
    port map (
            O => \N__3266\,
            I => \N__3263\
        );

    \I__548\ : Span12Mux_h
    port map (
            O => \N__3263\,
            I => \N__3260\
        );

    \I__547\ : Odrv12
    port map (
            O => \N__3260\,
            I => \D_LL_AMIGA_in_5\
        );

    \I__546\ : IoInMux
    port map (
            O => \N__3257\,
            I => \N__3254\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__3254\,
            I => \N__3251\
        );

    \I__544\ : IoSpan4Mux
    port map (
            O => \N__3251\,
            I => \N__3248\
        );

    \I__543\ : Sp12to4
    port map (
            O => \N__3248\,
            I => \N__3245\
        );

    \I__542\ : Span12Mux_s7_h
    port map (
            O => \N__3245\,
            I => \N__3242\
        );

    \I__541\ : Span12Mux_h
    port map (
            O => \N__3242\,
            I => \N__3239\
        );

    \I__540\ : Odrv12
    port map (
            O => \N__3239\,
            I => \un1_D_LL_AMIGA_5\
        );

    \I__539\ : InMux
    port map (
            O => \N__3236\,
            I => \N__3233\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3233\,
            I => \N__3230\
        );

    \I__537\ : Span12Mux_h
    port map (
            O => \N__3230\,
            I => \N__3227\
        );

    \I__536\ : Odrv12
    port map (
            O => \N__3227\,
            I => \D_LM_AMIGA_in_1\
        );

    \I__535\ : IoInMux
    port map (
            O => \N__3224\,
            I => \N__3221\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__3221\,
            I => \N__3218\
        );

    \I__533\ : Span4Mux_s2_h
    port map (
            O => \N__3218\,
            I => \N__3215\
        );

    \I__532\ : Span4Mux_v
    port map (
            O => \N__3215\,
            I => \N__3212\
        );

    \I__531\ : Span4Mux_h
    port map (
            O => \N__3212\,
            I => \N__3209\
        );

    \I__530\ : Sp12to4
    port map (
            O => \N__3209\,
            I => \N__3206\
        );

    \I__529\ : Span12Mux_h
    port map (
            O => \N__3206\,
            I => \N__3203\
        );

    \I__528\ : Odrv12
    port map (
            O => \N__3203\,
            I => \un1_D_LM_AMIGA_1\
        );

    \I__527\ : InMux
    port map (
            O => \N__3200\,
            I => \N__3197\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__3197\,
            I => \N__3194\
        );

    \I__525\ : Span12Mux_h
    port map (
            O => \N__3194\,
            I => \N__3191\
        );

    \I__524\ : Odrv12
    port map (
            O => \N__3191\,
            I => \D_LM_AMIGA_in_3\
        );

    \I__523\ : IoInMux
    port map (
            O => \N__3188\,
            I => \N__3185\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__3185\,
            I => \N__3182\
        );

    \I__521\ : Span12Mux_s7_h
    port map (
            O => \N__3182\,
            I => \N__3179\
        );

    \I__520\ : Span12Mux_h
    port map (
            O => \N__3179\,
            I => \N__3176\
        );

    \I__519\ : Odrv12
    port map (
            O => \N__3176\,
            I => \un1_D_LM_AMIGA_3\
        );

    \I__518\ : InMux
    port map (
            O => \N__3173\,
            I => \N__3170\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3170\,
            I => \N__3167\
        );

    \I__516\ : Span4Mux_v
    port map (
            O => \N__3167\,
            I => \N__3164\
        );

    \I__515\ : Sp12to4
    port map (
            O => \N__3164\,
            I => \N__3161\
        );

    \I__514\ : Span12Mux_h
    port map (
            O => \N__3161\,
            I => \N__3158\
        );

    \I__513\ : Odrv12
    port map (
            O => \N__3158\,
            I => \D_UM_040_in_6\
        );

    \I__512\ : IoInMux
    port map (
            O => \N__3155\,
            I => \N__3152\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__3152\,
            I => \N__3149\
        );

    \I__510\ : IoSpan4Mux
    port map (
            O => \N__3149\,
            I => \N__3145\
        );

    \I__509\ : InMux
    port map (
            O => \N__3148\,
            I => \N__3142\
        );

    \I__508\ : IoSpan4Mux
    port map (
            O => \N__3145\,
            I => \N__3139\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__3142\,
            I => \N__3136\
        );

    \I__506\ : Span4Mux_s2_h
    port map (
            O => \N__3139\,
            I => \N__3133\
        );

    \I__505\ : Span4Mux_v
    port map (
            O => \N__3136\,
            I => \N__3130\
        );

    \I__504\ : Sp12to4
    port map (
            O => \N__3133\,
            I => \N__3127\
        );

    \I__503\ : Sp12to4
    port map (
            O => \N__3130\,
            I => \N__3124\
        );

    \I__502\ : Span12Mux_h
    port map (
            O => \N__3127\,
            I => \N__3119\
        );

    \I__501\ : Span12Mux_v
    port map (
            O => \N__3124\,
            I => \N__3119\
        );

    \I__500\ : Span12Mux_h
    port map (
            O => \N__3119\,
            I => \N__3116\
        );

    \I__499\ : Odrv12
    port map (
            O => \N__3116\,
            I => \D_LL_040_in_6\
        );

    \I__498\ : IoInMux
    port map (
            O => \N__3113\,
            I => \N__3110\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3110\,
            I => \N__3107\
        );

    \I__496\ : Span12Mux_s10_h
    port map (
            O => \N__3107\,
            I => \N__3104\
        );

    \I__495\ : Span12Mux_v
    port map (
            O => \N__3104\,
            I => \N__3101\
        );

    \I__494\ : Odrv12
    port map (
            O => \N__3101\,
            I => \un1_D_UM_040_6\
        );

    \I__493\ : InMux
    port map (
            O => \N__3098\,
            I => \N__3095\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__3095\,
            I => \N__3092\
        );

    \I__491\ : Span4Mux_v
    port map (
            O => \N__3092\,
            I => \N__3089\
        );

    \I__490\ : Sp12to4
    port map (
            O => \N__3089\,
            I => \N__3086\
        );

    \I__489\ : Odrv12
    port map (
            O => \N__3086\,
            I => \D_LM_AMIGA_in_5\
        );

    \I__488\ : IoInMux
    port map (
            O => \N__3083\,
            I => \N__3080\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__3080\,
            I => \N__3077\
        );

    \I__486\ : IoSpan4Mux
    port map (
            O => \N__3077\,
            I => \N__3074\
        );

    \I__485\ : Sp12to4
    port map (
            O => \N__3074\,
            I => \N__3071\
        );

    \I__484\ : Span12Mux_s7_h
    port map (
            O => \N__3071\,
            I => \N__3068\
        );

    \I__483\ : Span12Mux_h
    port map (
            O => \N__3068\,
            I => \N__3065\
        );

    \I__482\ : Odrv12
    port map (
            O => \N__3065\,
            I => \un1_D_LM_AMIGA_5\
        );

    \I__481\ : InMux
    port map (
            O => \N__3062\,
            I => \N__3059\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3059\,
            I => \N__3056\
        );

    \I__479\ : Span4Mux_v
    port map (
            O => \N__3056\,
            I => \N__3053\
        );

    \I__478\ : Span4Mux_h
    port map (
            O => \N__3053\,
            I => \N__3050\
        );

    \I__477\ : Sp12to4
    port map (
            O => \N__3050\,
            I => \N__3047\
        );

    \I__476\ : Span12Mux_h
    port map (
            O => \N__3047\,
            I => \N__3044\
        );

    \I__475\ : Odrv12
    port map (
            O => \N__3044\,
            I => \D_UU_040_in_5\
        );

    \I__474\ : IoInMux
    port map (
            O => \N__3041\,
            I => \N__3038\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__3038\,
            I => \N__3035\
        );

    \I__472\ : IoSpan4Mux
    port map (
            O => \N__3035\,
            I => \N__3032\
        );

    \I__471\ : IoSpan4Mux
    port map (
            O => \N__3032\,
            I => \N__3029\
        );

    \I__470\ : Span4Mux_s2_h
    port map (
            O => \N__3029\,
            I => \N__3025\
        );

    \I__469\ : InMux
    port map (
            O => \N__3028\,
            I => \N__3022\
        );

    \I__468\ : Sp12to4
    port map (
            O => \N__3025\,
            I => \N__3019\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__3022\,
            I => \N__3016\
        );

    \I__466\ : Span12Mux_h
    port map (
            O => \N__3019\,
            I => \N__3011\
        );

    \I__465\ : Sp12to4
    port map (
            O => \N__3016\,
            I => \N__3011\
        );

    \I__464\ : Span12Mux_v
    port map (
            O => \N__3011\,
            I => \N__3008\
        );

    \I__463\ : Span12Mux_h
    port map (
            O => \N__3008\,
            I => \N__3005\
        );

    \I__462\ : Span12Mux_v
    port map (
            O => \N__3005\,
            I => \N__3002\
        );

    \I__461\ : Odrv12
    port map (
            O => \N__3002\,
            I => \D_LM_040_in_5\
        );

    \I__460\ : IoInMux
    port map (
            O => \N__2999\,
            I => \N__2996\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__2996\,
            I => \N__2993\
        );

    \I__458\ : Span12Mux_s0_h
    port map (
            O => \N__2993\,
            I => \N__2990\
        );

    \I__457\ : Span12Mux_h
    port map (
            O => \N__2990\,
            I => \N__2987\
        );

    \I__456\ : Odrv12
    port map (
            O => \N__2987\,
            I => \un1_D_UU_040_5\
        );

    \I__455\ : InMux
    port map (
            O => \N__2984\,
            I => \N__2981\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__2981\,
            I => \N__2978\
        );

    \I__453\ : Span4Mux_v
    port map (
            O => \N__2978\,
            I => \N__2975\
        );

    \I__452\ : Sp12to4
    port map (
            O => \N__2975\,
            I => \N__2972\
        );

    \I__451\ : Odrv12
    port map (
            O => \N__2972\,
            I => \D_LL_AMIGA_in_7\
        );

    \I__450\ : IoInMux
    port map (
            O => \N__2969\,
            I => \N__2966\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__2966\,
            I => \N__2963\
        );

    \I__448\ : Span4Mux_s1_h
    port map (
            O => \N__2963\,
            I => \N__2960\
        );

    \I__447\ : Sp12to4
    port map (
            O => \N__2960\,
            I => \N__2957\
        );

    \I__446\ : Span12Mux_v
    port map (
            O => \N__2957\,
            I => \N__2954\
        );

    \I__445\ : Span12Mux_h
    port map (
            O => \N__2954\,
            I => \N__2951\
        );

    \I__444\ : Odrv12
    port map (
            O => \N__2951\,
            I => \un1_D_LL_AMIGA_7\
        );

    \I__443\ : InMux
    port map (
            O => \N__2948\,
            I => \N__2945\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__2945\,
            I => \N__2942\
        );

    \I__441\ : Span4Mux_v
    port map (
            O => \N__2942\,
            I => \N__2939\
        );

    \I__440\ : Sp12to4
    port map (
            O => \N__2939\,
            I => \N__2936\
        );

    \I__439\ : Odrv12
    port map (
            O => \N__2936\,
            I => \D_LM_AMIGA_in_0\
        );

    \I__438\ : IoInMux
    port map (
            O => \N__2933\,
            I => \N__2930\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__2930\,
            I => \N__2927\
        );

    \I__436\ : Span12Mux_s9_h
    port map (
            O => \N__2927\,
            I => \N__2924\
        );

    \I__435\ : Span12Mux_h
    port map (
            O => \N__2924\,
            I => \N__2921\
        );

    \I__434\ : Odrv12
    port map (
            O => \N__2921\,
            I => \un1_D_LM_AMIGA_0\
        );

    \I__433\ : InMux
    port map (
            O => \N__2918\,
            I => \N__2915\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__2915\,
            I => \N__2912\
        );

    \I__431\ : Span4Mux_h
    port map (
            O => \N__2912\,
            I => \N__2909\
        );

    \I__430\ : Span4Mux_v
    port map (
            O => \N__2909\,
            I => \N__2906\
        );

    \I__429\ : Span4Mux_h
    port map (
            O => \N__2906\,
            I => \N__2903\
        );

    \I__428\ : Odrv4
    port map (
            O => \N__2903\,
            I => \D_LM_AMIGA_in_6\
        );

    \I__427\ : IoInMux
    port map (
            O => \N__2900\,
            I => \N__2897\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__2897\,
            I => \N__2894\
        );

    \I__425\ : Span12Mux_s4_h
    port map (
            O => \N__2894\,
            I => \N__2891\
        );

    \I__424\ : Span12Mux_h
    port map (
            O => \N__2891\,
            I => \N__2888\
        );

    \I__423\ : Odrv12
    port map (
            O => \N__2888\,
            I => \un1_D_LM_AMIGA_6\
        );

    \I__422\ : IoInMux
    port map (
            O => \N__2885\,
            I => \N__2882\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__2882\,
            I => \N__2879\
        );

    \I__420\ : IoSpan4Mux
    port map (
            O => \N__2879\,
            I => \N__2875\
        );

    \I__419\ : InMux
    port map (
            O => \N__2878\,
            I => \N__2872\
        );

    \I__418\ : IoSpan4Mux
    port map (
            O => \N__2875\,
            I => \N__2869\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__2872\,
            I => \N__2866\
        );

    \I__416\ : Span4Mux_s2_h
    port map (
            O => \N__2869\,
            I => \N__2863\
        );

    \I__415\ : Span4Mux_v
    port map (
            O => \N__2866\,
            I => \N__2860\
        );

    \I__414\ : Sp12to4
    port map (
            O => \N__2863\,
            I => \N__2857\
        );

    \I__413\ : Sp12to4
    port map (
            O => \N__2860\,
            I => \N__2854\
        );

    \I__412\ : Span12Mux_h
    port map (
            O => \N__2857\,
            I => \N__2851\
        );

    \I__411\ : Span12Mux_h
    port map (
            O => \N__2854\,
            I => \N__2848\
        );

    \I__410\ : Span12Mux_h
    port map (
            O => \N__2851\,
            I => \N__2845\
        );

    \I__409\ : Span12Mux_v
    port map (
            O => \N__2848\,
            I => \N__2842\
        );

    \I__408\ : Odrv12
    port map (
            O => \N__2845\,
            I => \D_LM_040_in_3\
        );

    \I__407\ : Odrv12
    port map (
            O => \N__2842\,
            I => \D_LM_040_in_3\
        );

    \I__406\ : InMux
    port map (
            O => \N__2837\,
            I => \N__2834\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__2834\,
            I => \N__2831\
        );

    \I__404\ : Span4Mux_v
    port map (
            O => \N__2831\,
            I => \N__2828\
        );

    \I__403\ : Sp12to4
    port map (
            O => \N__2828\,
            I => \N__2825\
        );

    \I__402\ : Span12Mux_h
    port map (
            O => \N__2825\,
            I => \N__2822\
        );

    \I__401\ : Span12Mux_h
    port map (
            O => \N__2822\,
            I => \N__2819\
        );

    \I__400\ : Odrv12
    port map (
            O => \N__2819\,
            I => \D_UU_040_in_3\
        );

    \I__399\ : IoInMux
    port map (
            O => \N__2816\,
            I => \N__2813\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__2813\,
            I => \N__2810\
        );

    \I__397\ : IoSpan4Mux
    port map (
            O => \N__2810\,
            I => \N__2807\
        );

    \I__396\ : IoSpan4Mux
    port map (
            O => \N__2807\,
            I => \N__2804\
        );

    \I__395\ : Span4Mux_s2_v
    port map (
            O => \N__2804\,
            I => \N__2801\
        );

    \I__394\ : Span4Mux_v
    port map (
            O => \N__2801\,
            I => \N__2798\
        );

    \I__393\ : Odrv4
    port map (
            O => \N__2798\,
            I => \un1_D_UU_040_3\
        );

    \I__392\ : IoInMux
    port map (
            O => \N__2795\,
            I => \N__2791\
        );

    \I__391\ : InMux
    port map (
            O => \N__2794\,
            I => \N__2788\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__2791\,
            I => \N__2785\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__2788\,
            I => \N__2782\
        );

    \I__388\ : Span4Mux_s2_h
    port map (
            O => \N__2785\,
            I => \N__2779\
        );

    \I__387\ : Span4Mux_h
    port map (
            O => \N__2782\,
            I => \N__2776\
        );

    \I__386\ : Sp12to4
    port map (
            O => \N__2779\,
            I => \N__2773\
        );

    \I__385\ : Sp12to4
    port map (
            O => \N__2776\,
            I => \N__2770\
        );

    \I__384\ : Span12Mux_h
    port map (
            O => \N__2773\,
            I => \N__2765\
        );

    \I__383\ : Span12Mux_v
    port map (
            O => \N__2770\,
            I => \N__2765\
        );

    \I__382\ : Span12Mux_v
    port map (
            O => \N__2765\,
            I => \N__2762\
        );

    \I__381\ : Span12Mux_h
    port map (
            O => \N__2762\,
            I => \N__2759\
        );

    \I__380\ : Odrv12
    port map (
            O => \N__2759\,
            I => \D_LM_040_in_2\
        );

    \I__379\ : InMux
    port map (
            O => \N__2756\,
            I => \N__2753\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__2753\,
            I => \N__2750\
        );

    \I__377\ : Span4Mux_v
    port map (
            O => \N__2750\,
            I => \N__2747\
        );

    \I__376\ : Span4Mux_h
    port map (
            O => \N__2747\,
            I => \N__2744\
        );

    \I__375\ : Sp12to4
    port map (
            O => \N__2744\,
            I => \N__2741\
        );

    \I__374\ : Span12Mux_h
    port map (
            O => \N__2741\,
            I => \N__2738\
        );

    \I__373\ : Odrv12
    port map (
            O => \N__2738\,
            I => \D_UU_040_in_2\
        );

    \I__372\ : IoInMux
    port map (
            O => \N__2735\,
            I => \N__2732\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__2732\,
            I => \N__2729\
        );

    \I__370\ : IoSpan4Mux
    port map (
            O => \N__2729\,
            I => \N__2726\
        );

    \I__369\ : IoSpan4Mux
    port map (
            O => \N__2726\,
            I => \N__2723\
        );

    \I__368\ : Span4Mux_s3_v
    port map (
            O => \N__2723\,
            I => \N__2720\
        );

    \I__367\ : Odrv4
    port map (
            O => \N__2720\,
            I => \un1_D_UU_040_2\
        );

    \I__366\ : InMux
    port map (
            O => \N__2717\,
            I => \N__2714\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__2714\,
            I => \N__2711\
        );

    \I__364\ : Span4Mux_v
    port map (
            O => \N__2711\,
            I => \N__2708\
        );

    \I__363\ : Span4Mux_h
    port map (
            O => \N__2708\,
            I => \N__2705\
        );

    \I__362\ : Span4Mux_h
    port map (
            O => \N__2705\,
            I => \N__2702\
        );

    \I__361\ : Odrv4
    port map (
            O => \N__2702\,
            I => \D_LL_AMIGA_in_0\
        );

    \I__360\ : IoInMux
    port map (
            O => \N__2699\,
            I => \N__2696\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__2696\,
            I => \N__2693\
        );

    \I__358\ : Span4Mux_s0_h
    port map (
            O => \N__2693\,
            I => \N__2690\
        );

    \I__357\ : Sp12to4
    port map (
            O => \N__2690\,
            I => \N__2687\
        );

    \I__356\ : Span12Mux_s6_v
    port map (
            O => \N__2687\,
            I => \N__2684\
        );

    \I__355\ : Span12Mux_h
    port map (
            O => \N__2684\,
            I => \N__2681\
        );

    \I__354\ : Odrv12
    port map (
            O => \N__2681\,
            I => \un1_D_LL_AMIGA_0\
        );

    \I__353\ : InMux
    port map (
            O => \N__2678\,
            I => \N__2675\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__2675\,
            I => \N__2672\
        );

    \I__351\ : Span4Mux_v
    port map (
            O => \N__2672\,
            I => \N__2669\
        );

    \I__350\ : Sp12to4
    port map (
            O => \N__2669\,
            I => \N__2666\
        );

    \I__349\ : Odrv12
    port map (
            O => \N__2666\,
            I => \D_LL_AMIGA_in_4\
        );

    \I__348\ : IoInMux
    port map (
            O => \N__2663\,
            I => \N__2660\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__2660\,
            I => \N__2657\
        );

    \I__346\ : IoSpan4Mux
    port map (
            O => \N__2657\,
            I => \N__2654\
        );

    \I__345\ : Span4Mux_s1_h
    port map (
            O => \N__2654\,
            I => \N__2651\
        );

    \I__344\ : Span4Mux_v
    port map (
            O => \N__2651\,
            I => \N__2648\
        );

    \I__343\ : Sp12to4
    port map (
            O => \N__2648\,
            I => \N__2645\
        );

    \I__342\ : Span12Mux_s10_h
    port map (
            O => \N__2645\,
            I => \N__2642\
        );

    \I__341\ : Odrv12
    port map (
            O => \N__2642\,
            I => \un1_D_LL_AMIGA_4\
        );

    \I__340\ : IoInMux
    port map (
            O => \N__2639\,
            I => \N__2636\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__2636\,
            I => \N__2632\
        );

    \I__338\ : InMux
    port map (
            O => \N__2635\,
            I => \N__2629\
        );

    \I__337\ : IoSpan4Mux
    port map (
            O => \N__2632\,
            I => \N__2626\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2629\,
            I => \N__2623\
        );

    \I__335\ : Span4Mux_s2_h
    port map (
            O => \N__2626\,
            I => \N__2620\
        );

    \I__334\ : Span4Mux_v
    port map (
            O => \N__2623\,
            I => \N__2617\
        );

    \I__333\ : Sp12to4
    port map (
            O => \N__2620\,
            I => \N__2614\
        );

    \I__332\ : Sp12to4
    port map (
            O => \N__2617\,
            I => \N__2611\
        );

    \I__331\ : Span12Mux_h
    port map (
            O => \N__2614\,
            I => \N__2608\
        );

    \I__330\ : Span12Mux_h
    port map (
            O => \N__2611\,
            I => \N__2605\
        );

    \I__329\ : Span12Mux_h
    port map (
            O => \N__2608\,
            I => \N__2600\
        );

    \I__328\ : Span12Mux_v
    port map (
            O => \N__2605\,
            I => \N__2600\
        );

    \I__327\ : Odrv12
    port map (
            O => \N__2600\,
            I => \D_LL_040_in_2\
        );

    \I__326\ : InMux
    port map (
            O => \N__2597\,
            I => \N__2594\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__2594\,
            I => \N__2591\
        );

    \I__324\ : Span12Mux_h
    port map (
            O => \N__2591\,
            I => \N__2588\
        );

    \I__323\ : Odrv12
    port map (
            O => \N__2588\,
            I => \D_UM_040_in_2\
        );

    \I__322\ : IoInMux
    port map (
            O => \N__2585\,
            I => \N__2582\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__2582\,
            I => \N__2579\
        );

    \I__320\ : Span4Mux_s2_h
    port map (
            O => \N__2579\,
            I => \N__2576\
        );

    \I__319\ : Span4Mux_v
    port map (
            O => \N__2576\,
            I => \N__2573\
        );

    \I__318\ : Sp12to4
    port map (
            O => \N__2573\,
            I => \N__2570\
        );

    \I__317\ : Odrv12
    port map (
            O => \N__2570\,
            I => \un1_D_UM_040_2\
        );

    \I__316\ : InMux
    port map (
            O => \N__2567\,
            I => \N__2564\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__2564\,
            I => \N__2561\
        );

    \I__314\ : Span4Mux_h
    port map (
            O => \N__2561\,
            I => \N__2558\
        );

    \I__313\ : Span4Mux_v
    port map (
            O => \N__2558\,
            I => \N__2555\
        );

    \I__312\ : Odrv4
    port map (
            O => \N__2555\,
            I => \A_040_c_0\
        );

    \I__311\ : IoInMux
    port map (
            O => \N__2552\,
            I => \N__2549\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__2549\,
            I => \N__2546\
        );

    \I__309\ : Span4Mux_s2_v
    port map (
            O => \N__2546\,
            I => \N__2543\
        );

    \I__308\ : Span4Mux_v
    port map (
            O => \N__2543\,
            I => \N__2540\
        );

    \I__307\ : Odrv4
    port map (
            O => \N__2540\,
            I => \A_AMIGA_c_0\
        );

    \I__306\ : InMux
    port map (
            O => \N__2537\,
            I => \N__2534\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__2534\,
            I => \N__2531\
        );

    \I__304\ : Span12Mux_h
    port map (
            O => \N__2531\,
            I => \N__2528\
        );

    \I__303\ : Odrv12
    port map (
            O => \N__2528\,
            I => \A_040_c_1\
        );

    \I__302\ : IoInMux
    port map (
            O => \N__2525\,
            I => \N__2512\
        );

    \I__301\ : IoInMux
    port map (
            O => \N__2524\,
            I => \N__2509\
        );

    \I__300\ : IoInMux
    port map (
            O => \N__2523\,
            I => \N__2506\
        );

    \I__299\ : IoInMux
    port map (
            O => \N__2522\,
            I => \N__2503\
        );

    \I__298\ : IoInMux
    port map (
            O => \N__2521\,
            I => \N__2496\
        );

    \I__297\ : IoInMux
    port map (
            O => \N__2520\,
            I => \N__2493\
        );

    \I__296\ : IoInMux
    port map (
            O => \N__2519\,
            I => \N__2490\
        );

    \I__295\ : IoInMux
    port map (
            O => \N__2518\,
            I => \N__2484\
        );

    \I__294\ : IoInMux
    port map (
            O => \N__2517\,
            I => \N__2481\
        );

    \I__293\ : IoInMux
    port map (
            O => \N__2516\,
            I => \N__2478\
        );

    \I__292\ : IoInMux
    port map (
            O => \N__2515\,
            I => \N__2475\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__2512\,
            I => \N__2466\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__2509\,
            I => \N__2466\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__2506\,
            I => \N__2466\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__2503\,
            I => \N__2466\
        );

    \I__287\ : IoInMux
    port map (
            O => \N__2502\,
            I => \N__2463\
        );

    \I__286\ : IoInMux
    port map (
            O => \N__2501\,
            I => \N__2460\
        );

    \I__285\ : IoInMux
    port map (
            O => \N__2500\,
            I => \N__2457\
        );

    \I__284\ : IoInMux
    port map (
            O => \N__2499\,
            I => \N__2454\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__2496\,
            I => \N__2443\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__2493\,
            I => \N__2443\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__2490\,
            I => \N__2443\
        );

    \I__280\ : IoInMux
    port map (
            O => \N__2489\,
            I => \N__2440\
        );

    \I__279\ : IoInMux
    port map (
            O => \N__2488\,
            I => \N__2437\
        );

    \I__278\ : IoInMux
    port map (
            O => \N__2487\,
            I => \N__2434\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__2484\,
            I => \N__2425\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__2481\,
            I => \N__2425\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2478\,
            I => \N__2425\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__2475\,
            I => \N__2425\
        );

    \I__273\ : IoSpan4Mux
    port map (
            O => \N__2466\,
            I => \N__2412\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__2463\,
            I => \N__2412\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__2460\,
            I => \N__2412\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2457\,
            I => \N__2412\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__2454\,
            I => \N__2412\
        );

    \I__268\ : IoInMux
    port map (
            O => \N__2453\,
            I => \N__2409\
        );

    \I__267\ : IoInMux
    port map (
            O => \N__2452\,
            I => \N__2406\
        );

    \I__266\ : IoInMux
    port map (
            O => \N__2451\,
            I => \N__2403\
        );

    \I__265\ : IoInMux
    port map (
            O => \N__2450\,
            I => \N__2400\
        );

    \I__264\ : IoSpan4Mux
    port map (
            O => \N__2443\,
            I => \N__2387\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__2440\,
            I => \N__2387\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__2437\,
            I => \N__2387\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__2434\,
            I => \N__2387\
        );

    \I__260\ : IoSpan4Mux
    port map (
            O => \N__2425\,
            I => \N__2384\
        );

    \I__259\ : IoInMux
    port map (
            O => \N__2424\,
            I => \N__2381\
        );

    \I__258\ : IoInMux
    port map (
            O => \N__2423\,
            I => \N__2378\
        );

    \I__257\ : IoSpan4Mux
    port map (
            O => \N__2412\,
            I => \N__2367\
        );

    \I__256\ : LocalMux
    port map (
            O => \N__2409\,
            I => \N__2367\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__2406\,
            I => \N__2367\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__2403\,
            I => \N__2367\
        );

    \I__253\ : LocalMux
    port map (
            O => \N__2400\,
            I => \N__2367\
        );

    \I__252\ : IoInMux
    port map (
            O => \N__2399\,
            I => \N__2364\
        );

    \I__251\ : IoInMux
    port map (
            O => \N__2398\,
            I => \N__2361\
        );

    \I__250\ : IoInMux
    port map (
            O => \N__2397\,
            I => \N__2358\
        );

    \I__249\ : IoInMux
    port map (
            O => \N__2396\,
            I => \N__2355\
        );

    \I__248\ : IoSpan4Mux
    port map (
            O => \N__2387\,
            I => \N__2352\
        );

    \I__247\ : Span4Mux_s3_h
    port map (
            O => \N__2384\,
            I => \N__2347\
        );

    \I__246\ : LocalMux
    port map (
            O => \N__2381\,
            I => \N__2342\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__2378\,
            I => \N__2342\
        );

    \I__244\ : IoSpan4Mux
    port map (
            O => \N__2367\,
            I => \N__2333\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__2364\,
            I => \N__2333\
        );

    \I__242\ : LocalMux
    port map (
            O => \N__2361\,
            I => \N__2333\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__2358\,
            I => \N__2333\
        );

    \I__240\ : LocalMux
    port map (
            O => \N__2355\,
            I => \N__2328\
        );

    \I__239\ : Span4Mux_s3_v
    port map (
            O => \N__2352\,
            I => \N__2325\
        );

    \I__238\ : IoInMux
    port map (
            O => \N__2351\,
            I => \N__2322\
        );

    \I__237\ : IoInMux
    port map (
            O => \N__2350\,
            I => \N__2319\
        );

    \I__236\ : Span4Mux_v
    port map (
            O => \N__2347\,
            I => \N__2314\
        );

    \I__235\ : Span4Mux_s3_h
    port map (
            O => \N__2342\,
            I => \N__2314\
        );

    \I__234\ : IoSpan4Mux
    port map (
            O => \N__2333\,
            I => \N__2311\
        );

    \I__233\ : IoInMux
    port map (
            O => \N__2332\,
            I => \N__2308\
        );

    \I__232\ : IoInMux
    port map (
            O => \N__2331\,
            I => \N__2305\
        );

    \I__231\ : Span12Mux_s5_v
    port map (
            O => \N__2328\,
            I => \N__2302\
        );

    \I__230\ : Span4Mux_v
    port map (
            O => \N__2325\,
            I => \N__2299\
        );

    \I__229\ : LocalMux
    port map (
            O => \N__2322\,
            I => \N__2294\
        );

    \I__228\ : LocalMux
    port map (
            O => \N__2319\,
            I => \N__2294\
        );

    \I__227\ : Span4Mux_v
    port map (
            O => \N__2314\,
            I => \N__2289\
        );

    \I__226\ : Span4Mux_s3_h
    port map (
            O => \N__2311\,
            I => \N__2289\
        );

    \I__225\ : LocalMux
    port map (
            O => \N__2308\,
            I => \N__2286\
        );

    \I__224\ : LocalMux
    port map (
            O => \N__2305\,
            I => \N__2283\
        );

    \I__223\ : Span12Mux_v
    port map (
            O => \N__2302\,
            I => \N__2280\
        );

    \I__222\ : Sp12to4
    port map (
            O => \N__2299\,
            I => \N__2275\
        );

    \I__221\ : Span12Mux_s9_h
    port map (
            O => \N__2294\,
            I => \N__2275\
        );

    \I__220\ : Span4Mux_h
    port map (
            O => \N__2289\,
            I => \N__2272\
        );

    \I__219\ : Span12Mux_s9_h
    port map (
            O => \N__2286\,
            I => \N__2267\
        );

    \I__218\ : Span12Mux_s9_h
    port map (
            O => \N__2283\,
            I => \N__2267\
        );

    \I__217\ : Odrv12
    port map (
            O => \N__2280\,
            I => \RnW_c_i_0\
        );

    \I__216\ : Odrv12
    port map (
            O => \N__2275\,
            I => \RnW_c_i_0\
        );

    \I__215\ : Odrv4
    port map (
            O => \N__2272\,
            I => \RnW_c_i_0\
        );

    \I__214\ : Odrv12
    port map (
            O => \N__2267\,
            I => \RnW_c_i_0\
        );

    \I__213\ : InMux
    port map (
            O => \N__2258\,
            I => \N__2255\
        );

    \I__212\ : LocalMux
    port map (
            O => \N__2255\,
            I => \N__2252\
        );

    \I__211\ : Span4Mux_v
    port map (
            O => \N__2252\,
            I => \N__2249\
        );

    \I__210\ : Sp12to4
    port map (
            O => \N__2249\,
            I => \N__2246\
        );

    \I__209\ : Odrv12
    port map (
            O => \N__2246\,
            I => \D_LL_AMIGA_in_3\
        );

    \I__208\ : IoInMux
    port map (
            O => \N__2243\,
            I => \N__2240\
        );

    \I__207\ : LocalMux
    port map (
            O => \N__2240\,
            I => \N__2237\
        );

    \I__206\ : IoSpan4Mux
    port map (
            O => \N__2237\,
            I => \N__2234\
        );

    \I__205\ : IoSpan4Mux
    port map (
            O => \N__2234\,
            I => \N__2231\
        );

    \I__204\ : Span4Mux_s2_h
    port map (
            O => \N__2231\,
            I => \N__2228\
        );

    \I__203\ : Sp12to4
    port map (
            O => \N__2228\,
            I => \N__2225\
        );

    \I__202\ : Span12Mux_s9_h
    port map (
            O => \N__2225\,
            I => \N__2222\
        );

    \I__201\ : Odrv12
    port map (
            O => \N__2222\,
            I => \un1_D_LL_AMIGA_3\
        );

    \I__200\ : InMux
    port map (
            O => \N__2219\,
            I => \N__2216\
        );

    \I__199\ : LocalMux
    port map (
            O => \N__2216\,
            I => \N__2212\
        );

    \I__198\ : IoInMux
    port map (
            O => \N__2215\,
            I => \N__2209\
        );

    \I__197\ : Span4Mux_v
    port map (
            O => \N__2212\,
            I => \N__2206\
        );

    \I__196\ : LocalMux
    port map (
            O => \N__2209\,
            I => \N__2203\
        );

    \I__195\ : Odrv4
    port map (
            O => \N__2206\,
            I => \A_AMIGA_c_1\
        );

    \I__194\ : Odrv12
    port map (
            O => \N__2203\,
            I => \A_AMIGA_c_1\
        );

    \INVU111_CYCLE_SM.UU_LATCHED_nesr_7C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UU_LATCHED_nesr_7C_net\,
            I => \N__4918\
        );

    \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            I => \N__4921\
        );

    \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net\,
            I => \N__4923\
        );

    \INVU111_CYCLE_SM.UU_LATCHED_nesr_0C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UU_LATCHED_nesr_0C_net\,
            I => \N__4915\
        );

    \INVU111_CYCLE_SM.CYCLE_STATE_1C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.CYCLE_STATE_1C_net\,
            I => \N__4916\
        );

    \INVU111_CYCLE_SM.UM_LATCHED_nesr_0C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UM_LATCHED_nesr_0C_net\,
            I => \N__4919\
        );

    \INVU111_CYCLE_SM.UU_LATCHED_nesr_4C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net\,
            I => \N__4917\
        );

    \INVU111_CYCLE_SM.TS_ENC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.TS_ENC_net\,
            I => \N__4920\
        );

    \INVU111_CYCLE_SM.A_OUTC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.A_OUTC_net\,
            I => \N__4922\
        );

    \INVU111_CYCLE_SM.TSnC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.TSnC_net\,
            I => \N__4791\
        );

    \INVU111_CYCLE_SM.TA_EN_nessC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.TA_EN_nessC_net\,
            I => \N__4927\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6637\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2567\,
            lcout => \A_AMIGA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__3452\,
            in1 => \N__2537\,
            in2 => \_gnd_net_\,
            in3 => \N__6636\,
            lcout => \A_AMIGA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RnW_c_sbtinv_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4607\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RnW_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIGCUI2_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5861\,
            in1 => \N__5967\,
            in2 => \_gnd_net_\,
            in3 => \N__2258\,
            lcout => \un1_D_LL_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIM3VM1_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__2219\,
            in1 => \N__6940\,
            in2 => \_gnd_net_\,
            in3 => \N__6638\,
            lcout => \U111_CYCLE_SM.FLIP\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIOKUI2_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2984\,
            in1 => \N__5969\,
            in2 => \_gnd_net_\,
            in3 => \N__5694\,
            lcout => \un1_D_LL_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIJDJF2_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5102\,
            in1 => \N__5968\,
            in2 => \_gnd_net_\,
            in3 => \N__2948\,
            lcout => \un1_D_LM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIVPJF2_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__3629\,
            in1 => \N__6054\,
            in2 => \_gnd_net_\,
            in3 => \N__2918\,
            lcout => \un1_D_LM_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI3JQV1_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__2878\,
            in1 => \N__6097\,
            in2 => \_gnd_net_\,
            in3 => \N__2837\,
            lcout => \un1_D_UU_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI1HQV1_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__2794\,
            in1 => \N__6096\,
            in2 => \_gnd_net_\,
            in3 => \N__2756\,
            lcout => \un1_D_UU_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIA6UI2_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2717\,
            in1 => \N__5973\,
            in2 => \_gnd_net_\,
            in3 => \N__3785\,
            lcout => \un1_D_LL_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIIEUI2_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2678\,
            in1 => \N__5930\,
            in2 => \_gnd_net_\,
            in3 => \N__4190\,
            lcout => \un1_D_LL_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIOROB2_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__2635\,
            in1 => \N__6077\,
            in2 => \_gnd_net_\,
            in3 => \N__2597\,
            lcout => \un1_D_UM_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNINHJF2_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6079\,
            in1 => \N__5608\,
            in2 => \_gnd_net_\,
            in3 => \N__3377\,
            lcout => \un1_D_LM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIBRQV1_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__3343\,
            in1 => \N__6138\,
            in2 => \_gnd_net_\,
            in3 => \N__3314\,
            lcout => \un1_D_UU_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIKGUI2_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6914\,
            in1 => \N__6025\,
            in2 => \_gnd_net_\,
            in3 => \N__3275\,
            lcout => \un1_D_LL_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNILFJF2_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__3236\,
            in1 => \N__6078\,
            in2 => \_gnd_net_\,
            in3 => \N__6466\,
            lcout => \un1_D_LM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIPJJF2_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6080\,
            in1 => \N__5459\,
            in2 => \_gnd_net_\,
            in3 => \N__3200\,
            lcout => \un1_D_LM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI04PB2_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6081\,
            in1 => \N__3173\,
            in2 => \_gnd_net_\,
            in3 => \N__3148\,
            lcout => \un1_D_UM_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNITNJF2_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6111\,
            in1 => \N__5529\,
            in2 => \_gnd_net_\,
            in3 => \N__3098\,
            lcout => \un1_D_LM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI7NQV1_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6139\,
            in1 => \N__3062\,
            in2 => \_gnd_net_\,
            in3 => \N__3028\,
            lcout => \un1_D_UU_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_EN_ness_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4715\,
            lcout => \U111_CYCLE_SM.TA_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TA_EN_nessC_net\,
            ce => \N__3413\,
            sr => \N__3424\
        );

    \RESETn_ibuf_RNIM9SF_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4322\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TSn_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__4323\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3694\,
            lcout => \TSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TSnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNISVOB2_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6134\,
            in1 => \N__3569\,
            in2 => \_gnd_net_\,
            in3 => \N__3544\,
            lcout => \un1_D_UM_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIC8UI2_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5201\,
            in1 => \N__6053\,
            in2 => \_gnd_net_\,
            in3 => \N__3491\,
            lcout => \un1_D_LL_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A_OUT_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__3445\,
            in1 => \N__3434\,
            in2 => \N__4333\,
            in3 => \N__4696\,
            lcout => \U111_CYCLE_SM.A_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.A_OUTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_START_RNIIU7U_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__6521\,
            in1 => \N__4661\,
            in2 => \N__3653\,
            in3 => \N__4695\,
            lcout => \U111_CYCLE_SM.un1_CYCLE_STATE_1_0\,
            ltout => \U111_CYCLE_SM.un1_CYCLE_STATE_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_EN_ness_RNO_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3428\,
            in3 => \N__3425\,
            lcout => \U111_CYCLE_SM.un1_CYCLE_STATE_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_EN_ness_RNIPNOD_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__3404\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4737\,
            lcout => \TAn_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIRLJF2_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6067\,
            in1 => \N__3974\,
            in2 => \_gnd_net_\,
            in3 => \N__3740\,
            lcout => \un1_D_LM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4662\,
            in2 => \_gnd_net_\,
            in3 => \N__4712\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.TS_EN10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__4331\,
            in1 => \N__4760\,
            in2 => \N__3698\,
            in3 => \N__3695\,
            lcout => \U111_CYCLE_SM.TS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TS_ENC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000100010"
        )
    port map (
            in0 => \N__3652\,
            in1 => \N__4663\,
            in2 => \N__4744\,
            in3 => \N__4713\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.LW_CYCLE_r_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110001000000"
        )
    port map (
            in0 => \N__4714\,
            in1 => \N__4327\,
            in2 => \N__3683\,
            in3 => \N__6522\,
            lcout => \U111_CYCLE_SM.LW_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TS_ENC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_START_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__6977\,
            in1 => \N__6941\,
            in2 => \N__4334\,
            in3 => \N__3664\,
            lcout => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TS_ENC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__3973\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net\,
            ce => \N__5300\,
            sr => \N__5254\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3628\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net\,
            ce => \N__5300\,
            sr => \N__5254\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__3638\,
            in1 => \N__3621\,
            in2 => \_gnd_net_\,
            in3 => \N__6616\,
            lcout => \un1_D_UU_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNITCQV1_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__4067\,
            in1 => \N__6110\,
            in2 => \_gnd_net_\,
            in3 => \N__4045\,
            lcout => \un1_D_UU_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6615\,
            in1 => \N__3983\,
            in2 => \_gnd_net_\,
            in3 => \N__3961\,
            lcout => \un1_D_UU_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIKNOB2_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6121\,
            in1 => \N__3916\,
            in2 => \_gnd_net_\,
            in3 => \N__3875\,
            lcout => \un1_D_UM_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK40_THRU_LUT4_0_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4802\,
            lcout => \GB_BUFFER_CLK40_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6553\,
            in1 => \N__3746\,
            in2 => \_gnd_net_\,
            in3 => \N__3778\,
            lcout => \un1_D_UM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3765\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_0C_net\,
            ce => \N__5298\,
            sr => \N__5251\
        );

    \U111_CYCLE_SM.CYCLE_STATE_1_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001101000000000"
        )
    port map (
            in0 => \N__4694\,
            in1 => \N__4753\,
            in2 => \N__4664\,
            in3 => \N__4320\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.CYCLE_STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__4752\,
            in1 => \N__4657\,
            in2 => \N__4332\,
            in3 => \N__4698\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.CYCLE_STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_1_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000010"
        )
    port map (
            in0 => \N__4801\,
            in1 => \N__4656\,
            in2 => \N__4778\,
            in3 => \N__4697\,
            lcout => \U111_CYCLE_SM.TS_EN_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIFCLM_0_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__4754\,
            in1 => \N__4693\,
            in2 => \_gnd_net_\,
            in3 => \N__4655\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa\,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1_0_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011111111"
        )
    port map (
            in0 => \N__4538\,
            in1 => \_gnd_net_\,
            in2 => \N__4337\,
            in3 => \N__4321\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0\,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIGG4C2_0_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4244\,
            in3 => \N__4241\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5095\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_0C_net\,
            ce => \N__5299\,
            sr => \N__5253\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4180\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_0C_net\,
            ce => \N__5299\,
            sr => \N__5253\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI1SJF2_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6835\,
            in1 => \N__6098\,
            in2 => \_gnd_net_\,
            in3 => \N__4235\,
            lcout => \un1_D_LM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4199\,
            in1 => \N__4173\,
            in2 => \_gnd_net_\,
            in3 => \N__6593\,
            lcout => \un1_D_UM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIU1PB2_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4114\,
            in1 => \N__6157\,
            in2 => \_gnd_net_\,
            in3 => \N__4085\,
            lcout => \un1_D_UM_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5114\,
            in1 => \N__5094\,
            in2 => \_gnd_net_\,
            in3 => \N__6629\,
            lcout => \un1_D_UU_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIEAUI2_LC_13_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6076\,
            in1 => \N__4849\,
            in2 => \_gnd_net_\,
            in3 => \N__5021\,
            lcout => \un1_D_LL_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIMIUI2_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6788\,
            in1 => \N__6092\,
            in2 => \_gnd_net_\,
            in3 => \N__4982\,
            lcout => \un1_D_LL_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4850\,
            in1 => \N__4811\,
            in2 => \_gnd_net_\,
            in3 => \N__6613\,
            lcout => \un1_D_UM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK80_THRU_LUT4_0_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4931\,
            lcout => \GB_BUFFER_CLK80_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6777\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net\,
            ce => \N__5302\,
            sr => \N__5252\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4845\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net\,
            ce => \N__5302\,
            sr => \N__5252\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5857\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            ce => \N__5301\,
            sr => \N__5238\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5609\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            ce => \N__5301\,
            sr => \N__5238\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6839\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_7C_net\,
            ce => \N__5303\,
            sr => \N__5258\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6467\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_7C_net\,
            ce => \N__5303\,
            sr => \N__5258\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5458\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_7C_net\,
            ce => \N__5303\,
            sr => \N__5258\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5534\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_7C_net\,
            ce => \N__5303\,
            sr => \N__5258\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5699\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_7C_net\,
            ce => \N__5303\,
            sr => \N__5258\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5197\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_7C_net\,
            ce => \N__5303\,
            sr => \N__5258\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6910\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_7C_net\,
            ce => \N__5303\,
            sr => \N__5258\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5196\,
            in1 => \N__5159\,
            in2 => \_gnd_net_\,
            in3 => \N__6592\,
            lcout => \un1_D_UM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5850\,
            in1 => \N__5813\,
            in2 => \_gnd_net_\,
            in3 => \N__6594\,
            lcout => \un1_D_UM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIQTOB2_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5783\,
            in1 => \N__6158\,
            in2 => \_gnd_net_\,
            in3 => \N__5738\,
            lcout => \un1_D_UM_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5695\,
            in1 => \N__5648\,
            in2 => \_gnd_net_\,
            in3 => \N__6626\,
            lcout => \un1_D_UM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5618\,
            in1 => \N__5589\,
            in2 => \_gnd_net_\,
            in3 => \N__6627\,
            lcout => \un1_D_UU_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6628\,
            in1 => \N__5546\,
            in2 => \_gnd_net_\,
            in3 => \N__5533\,
            lcout => \un1_D_UU_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6631\,
            in1 => \N__5468\,
            in2 => \_gnd_net_\,
            in3 => \N__5451\,
            lcout => \un1_D_UU_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI9PQV1_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__5393\,
            in1 => \N__6156\,
            in2 => \_gnd_net_\,
            in3 => \N__5371\,
            lcout => \un1_D_UU_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6630\,
            in1 => \N__5315\,
            in2 => \_gnd_net_\,
            in3 => \N__6906\,
            lcout => \un1_D_UM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6848\,
            in1 => \N__6828\,
            in2 => \_gnd_net_\,
            in3 => \N__6632\,
            lcout => \un1_D_UU_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6778\,
            in1 => \N__6752\,
            in2 => \_gnd_net_\,
            in3 => \N__6614\,
            lcout => \un1_D_UM_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIMPOB2_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6724\,
            in1 => \N__6143\,
            in2 => \_gnd_net_\,
            in3 => \N__6677\,
            lcout => \un1_D_UM_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6620\,
            in1 => \N__6479\,
            in2 => \_gnd_net_\,
            in3 => \N__6459\,
            lcout => \un1_D_UU_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIVEQV1_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6397\,
            in1 => \N__6159\,
            in2 => \_gnd_net_\,
            in3 => \N__6350\,
            lcout => \un1_D_UU_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI26PB2_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6301\,
            in1 => \N__6160\,
            in2 => \_gnd_net_\,
            in3 => \N__6254\,
            lcout => \un1_D_UM_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI5LQV1_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6208\,
            in1 => \N__6179\,
            in2 => \_gnd_net_\,
            in3 => \N__6161\,
            lcout => \un1_D_UU_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_TRANS_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__7016\,
            in1 => \N__6995\,
            in2 => \_gnd_net_\,
            in3 => \N__6973\,
            lcout => \U111_CYCLE_SM.LW_TRANS_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Dec 21 2024 14:06:00

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U409_TOP" view "INTERFACE"

module U409_TOP (
    A,
    RnW,
    CIACS1n,
    TT1,
    TICK50,
    RAMSPACEn,
    TT0,
    TICK60,
    LBENn,
    CLKCIA,
    CIACS0n,
    CLK6,
    CLK40_IN,
    CLK28_IN,
    REGSPACEn,
    BUFENn,
    TSn,
    RESETn,
    OVL,
    TACKn,
    ROMENn,
    PORTSIZE);

    input [31:1] A;
    input RnW;
    output CIACS1n;
    input TT1;
    output TICK50;
    output RAMSPACEn;
    input TT0;
    output TICK60;
    input LBENn;
    output CLKCIA;
    output CIACS0n;
    input CLK6;
    input CLK40_IN;
    input CLK28_IN;
    output REGSPACEn;
    output BUFENn;
    input TSn;
    input RESETn;
    input OVL;
    inout TACKn;
    output ROMENn;
    output PORTSIZE;

    wire N__6079;
    wire N__6078;
    wire N__6077;
    wire N__6069;
    wire N__6068;
    wire N__6067;
    wire N__6058;
    wire N__6057;
    wire N__6056;
    wire N__6049;
    wire N__6048;
    wire N__6047;
    wire N__6040;
    wire N__6039;
    wire N__6038;
    wire N__6031;
    wire N__6030;
    wire N__6029;
    wire N__6022;
    wire N__6021;
    wire N__6020;
    wire N__6013;
    wire N__6012;
    wire N__6011;
    wire N__6004;
    wire N__6003;
    wire N__6002;
    wire N__5995;
    wire N__5994;
    wire N__5993;
    wire N__5986;
    wire N__5985;
    wire N__5984;
    wire N__5977;
    wire N__5976;
    wire N__5975;
    wire N__5968;
    wire N__5967;
    wire N__5966;
    wire N__5959;
    wire N__5958;
    wire N__5957;
    wire N__5950;
    wire N__5949;
    wire N__5948;
    wire N__5941;
    wire N__5940;
    wire N__5939;
    wire N__5932;
    wire N__5931;
    wire N__5930;
    wire N__5923;
    wire N__5922;
    wire N__5921;
    wire N__5914;
    wire N__5913;
    wire N__5912;
    wire N__5905;
    wire N__5904;
    wire N__5903;
    wire N__5896;
    wire N__5895;
    wire N__5894;
    wire N__5887;
    wire N__5886;
    wire N__5885;
    wire N__5878;
    wire N__5877;
    wire N__5876;
    wire N__5869;
    wire N__5868;
    wire N__5867;
    wire N__5860;
    wire N__5859;
    wire N__5858;
    wire N__5851;
    wire N__5850;
    wire N__5849;
    wire N__5842;
    wire N__5841;
    wire N__5840;
    wire N__5833;
    wire N__5832;
    wire N__5831;
    wire N__5824;
    wire N__5823;
    wire N__5822;
    wire N__5815;
    wire N__5814;
    wire N__5813;
    wire N__5806;
    wire N__5805;
    wire N__5804;
    wire N__5797;
    wire N__5796;
    wire N__5795;
    wire N__5788;
    wire N__5787;
    wire N__5786;
    wire N__5779;
    wire N__5778;
    wire N__5777;
    wire N__5770;
    wire N__5769;
    wire N__5768;
    wire N__5751;
    wire N__5750;
    wire N__5749;
    wire N__5746;
    wire N__5745;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5727;
    wire N__5724;
    wire N__5721;
    wire N__5718;
    wire N__5715;
    wire N__5712;
    wire N__5711;
    wire N__5710;
    wire N__5709;
    wire N__5708;
    wire N__5707;
    wire N__5706;
    wire N__5705;
    wire N__5702;
    wire N__5699;
    wire N__5696;
    wire N__5689;
    wire N__5682;
    wire N__5673;
    wire N__5672;
    wire N__5671;
    wire N__5670;
    wire N__5669;
    wire N__5668;
    wire N__5667;
    wire N__5664;
    wire N__5657;
    wire N__5650;
    wire N__5643;
    wire N__5642;
    wire N__5641;
    wire N__5640;
    wire N__5631;
    wire N__5628;
    wire N__5625;
    wire N__5622;
    wire N__5619;
    wire N__5616;
    wire N__5613;
    wire N__5610;
    wire N__5607;
    wire N__5604;
    wire N__5601;
    wire N__5598;
    wire N__5595;
    wire N__5592;
    wire N__5589;
    wire N__5586;
    wire N__5583;
    wire N__5580;
    wire N__5577;
    wire N__5576;
    wire N__5573;
    wire N__5570;
    wire N__5567;
    wire N__5564;
    wire N__5559;
    wire N__5556;
    wire N__5553;
    wire N__5550;
    wire N__5547;
    wire N__5544;
    wire N__5541;
    wire N__5538;
    wire N__5537;
    wire N__5534;
    wire N__5533;
    wire N__5530;
    wire N__5529;
    wire N__5526;
    wire N__5525;
    wire N__5524;
    wire N__5523;
    wire N__5522;
    wire N__5521;
    wire N__5520;
    wire N__5517;
    wire N__5516;
    wire N__5515;
    wire N__5514;
    wire N__5513;
    wire N__5512;
    wire N__5511;
    wire N__5508;
    wire N__5505;
    wire N__5504;
    wire N__5501;
    wire N__5492;
    wire N__5489;
    wire N__5486;
    wire N__5479;
    wire N__5476;
    wire N__5469;
    wire N__5468;
    wire N__5463;
    wire N__5460;
    wire N__5459;
    wire N__5444;
    wire N__5441;
    wire N__5436;
    wire N__5435;
    wire N__5432;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5397;
    wire N__5392;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5375;
    wire N__5372;
    wire N__5367;
    wire N__5366;
    wire N__5365;
    wire N__5362;
    wire N__5359;
    wire N__5356;
    wire N__5353;
    wire N__5350;
    wire N__5347;
    wire N__5344;
    wire N__5341;
    wire N__5338;
    wire N__5335;
    wire N__5332;
    wire N__5329;
    wire N__5322;
    wire N__5319;
    wire N__5318;
    wire N__5315;
    wire N__5312;
    wire N__5307;
    wire N__5306;
    wire N__5305;
    wire N__5304;
    wire N__5303;
    wire N__5302;
    wire N__5301;
    wire N__5300;
    wire N__5299;
    wire N__5280;
    wire N__5277;
    wire N__5274;
    wire N__5271;
    wire N__5268;
    wire N__5265;
    wire N__5262;
    wire N__5259;
    wire N__5258;
    wire N__5257;
    wire N__5256;
    wire N__5251;
    wire N__5246;
    wire N__5241;
    wire N__5240;
    wire N__5239;
    wire N__5238;
    wire N__5237;
    wire N__5236;
    wire N__5227;
    wire N__5222;
    wire N__5217;
    wire N__5216;
    wire N__5213;
    wire N__5212;
    wire N__5211;
    wire N__5208;
    wire N__5203;
    wire N__5200;
    wire N__5193;
    wire N__5190;
    wire N__5189;
    wire N__5186;
    wire N__5183;
    wire N__5178;
    wire N__5175;
    wire N__5174;
    wire N__5171;
    wire N__5168;
    wire N__5163;
    wire N__5160;
    wire N__5157;
    wire N__5154;
    wire N__5151;
    wire N__5150;
    wire N__5147;
    wire N__5144;
    wire N__5139;
    wire N__5136;
    wire N__5133;
    wire N__5132;
    wire N__5129;
    wire N__5126;
    wire N__5121;
    wire N__5118;
    wire N__5115;
    wire N__5112;
    wire N__5109;
    wire N__5108;
    wire N__5105;
    wire N__5102;
    wire N__5097;
    wire N__5094;
    wire N__5093;
    wire N__5090;
    wire N__5087;
    wire N__5082;
    wire N__5079;
    wire N__5076;
    wire N__5073;
    wire N__5072;
    wire N__5069;
    wire N__5066;
    wire N__5061;
    wire N__5058;
    wire N__5055;
    wire N__5052;
    wire N__5051;
    wire N__5048;
    wire N__5045;
    wire N__5040;
    wire N__5037;
    wire N__5034;
    wire N__5031;
    wire N__5028;
    wire N__5025;
    wire N__5024;
    wire N__5023;
    wire N__5022;
    wire N__5021;
    wire N__5014;
    wire N__5009;
    wire N__5004;
    wire N__5001;
    wire N__5000;
    wire N__4999;
    wire N__4998;
    wire N__4995;
    wire N__4990;
    wire N__4987;
    wire N__4984;
    wire N__4977;
    wire N__4974;
    wire N__4971;
    wire N__4968;
    wire N__4965;
    wire N__4962;
    wire N__4961;
    wire N__4958;
    wire N__4957;
    wire N__4952;
    wire N__4949;
    wire N__4944;
    wire N__4943;
    wire N__4942;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4930;
    wire N__4927;
    wire N__4920;
    wire N__4919;
    wire N__4916;
    wire N__4913;
    wire N__4908;
    wire N__4905;
    wire N__4904;
    wire N__4901;
    wire N__4898;
    wire N__4893;
    wire N__4890;
    wire N__4887;
    wire N__4884;
    wire N__4881;
    wire N__4880;
    wire N__4877;
    wire N__4874;
    wire N__4869;
    wire N__4866;
    wire N__4865;
    wire N__4862;
    wire N__4859;
    wire N__4854;
    wire N__4851;
    wire N__4848;
    wire N__4845;
    wire N__4844;
    wire N__4841;
    wire N__4838;
    wire N__4833;
    wire N__4830;
    wire N__4827;
    wire N__4824;
    wire N__4823;
    wire N__4820;
    wire N__4817;
    wire N__4812;
    wire N__4809;
    wire N__4808;
    wire N__4803;
    wire N__4800;
    wire N__4799;
    wire N__4798;
    wire N__4797;
    wire N__4796;
    wire N__4795;
    wire N__4794;
    wire N__4791;
    wire N__4788;
    wire N__4785;
    wire N__4782;
    wire N__4773;
    wire N__4764;
    wire N__4763;
    wire N__4762;
    wire N__4761;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4747;
    wire N__4740;
    wire N__4739;
    wire N__4738;
    wire N__4735;
    wire N__4730;
    wire N__4725;
    wire N__4722;
    wire N__4719;
    wire N__4716;
    wire N__4713;
    wire N__4712;
    wire N__4711;
    wire N__4710;
    wire N__4705;
    wire N__4702;
    wire N__4699;
    wire N__4692;
    wire N__4689;
    wire N__4688;
    wire N__4687;
    wire N__4684;
    wire N__4683;
    wire N__4680;
    wire N__4679;
    wire N__4676;
    wire N__4673;
    wire N__4670;
    wire N__4667;
    wire N__4662;
    wire N__4659;
    wire N__4656;
    wire N__4653;
    wire N__4652;
    wire N__4649;
    wire N__4644;
    wire N__4641;
    wire N__4638;
    wire N__4633;
    wire N__4630;
    wire N__4627;
    wire N__4624;
    wire N__4621;
    wire N__4618;
    wire N__4615;
    wire N__4612;
    wire N__4609;
    wire N__4606;
    wire N__4599;
    wire N__4598;
    wire N__4597;
    wire N__4594;
    wire N__4591;
    wire N__4588;
    wire N__4585;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4565;
    wire N__4560;
    wire N__4557;
    wire N__4554;
    wire N__4553;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4539;
    wire N__4538;
    wire N__4537;
    wire N__4532;
    wire N__4529;
    wire N__4524;
    wire N__4521;
    wire N__4518;
    wire N__4515;
    wire N__4514;
    wire N__4513;
    wire N__4512;
    wire N__4509;
    wire N__4506;
    wire N__4501;
    wire N__4494;
    wire N__4493;
    wire N__4492;
    wire N__4485;
    wire N__4482;
    wire N__4481;
    wire N__4480;
    wire N__4477;
    wire N__4476;
    wire N__4475;
    wire N__4472;
    wire N__4463;
    wire N__4458;
    wire N__4455;
    wire N__4454;
    wire N__4453;
    wire N__4452;
    wire N__4451;
    wire N__4450;
    wire N__4449;
    wire N__4448;
    wire N__4443;
    wire N__4436;
    wire N__4429;
    wire N__4422;
    wire N__4421;
    wire N__4420;
    wire N__4419;
    wire N__4418;
    wire N__4417;
    wire N__4416;
    wire N__4415;
    wire N__4410;
    wire N__4403;
    wire N__4396;
    wire N__4389;
    wire N__4388;
    wire N__4387;
    wire N__4384;
    wire N__4383;
    wire N__4382;
    wire N__4379;
    wire N__4378;
    wire N__4377;
    wire N__4376;
    wire N__4371;
    wire N__4364;
    wire N__4357;
    wire N__4350;
    wire N__4347;
    wire N__4344;
    wire N__4341;
    wire N__4338;
    wire N__4335;
    wire N__4334;
    wire N__4331;
    wire N__4328;
    wire N__4323;
    wire N__4320;
    wire N__4317;
    wire N__4316;
    wire N__4313;
    wire N__4312;
    wire N__4309;
    wire N__4308;
    wire N__4305;
    wire N__4300;
    wire N__4297;
    wire N__4292;
    wire N__4287;
    wire N__4284;
    wire N__4281;
    wire N__4278;
    wire N__4275;
    wire N__4272;
    wire N__4269;
    wire N__4266;
    wire N__4263;
    wire N__4260;
    wire N__4257;
    wire N__4256;
    wire N__4255;
    wire N__4252;
    wire N__4249;
    wire N__4246;
    wire N__4239;
    wire N__4238;
    wire N__4235;
    wire N__4232;
    wire N__4227;
    wire N__4224;
    wire N__4221;
    wire N__4218;
    wire N__4215;
    wire N__4212;
    wire N__4209;
    wire N__4206;
    wire N__4203;
    wire N__4200;
    wire N__4197;
    wire N__4194;
    wire N__4193;
    wire N__4190;
    wire N__4187;
    wire N__4182;
    wire N__4179;
    wire N__4176;
    wire N__4173;
    wire N__4170;
    wire N__4167;
    wire N__4166;
    wire N__4163;
    wire N__4160;
    wire N__4155;
    wire N__4154;
    wire N__4151;
    wire N__4148;
    wire N__4143;
    wire N__4142;
    wire N__4139;
    wire N__4136;
    wire N__4131;
    wire N__4128;
    wire N__4125;
    wire N__4124;
    wire N__4121;
    wire N__4118;
    wire N__4113;
    wire N__4112;
    wire N__4109;
    wire N__4106;
    wire N__4101;
    wire N__4100;
    wire N__4099;
    wire N__4096;
    wire N__4095;
    wire N__4092;
    wire N__4091;
    wire N__4090;
    wire N__4089;
    wire N__4084;
    wire N__4079;
    wire N__4072;
    wire N__4065;
    wire N__4064;
    wire N__4063;
    wire N__4062;
    wire N__4059;
    wire N__4058;
    wire N__4057;
    wire N__4056;
    wire N__4055;
    wire N__4050;
    wire N__4043;
    wire N__4036;
    wire N__4029;
    wire N__4028;
    wire N__4027;
    wire N__4026;
    wire N__4019;
    wire N__4016;
    wire N__4015;
    wire N__4014;
    wire N__4013;
    wire N__4010;
    wire N__4007;
    wire N__4004;
    wire N__4001;
    wire N__3998;
    wire N__3995;
    wire N__3984;
    wire N__3981;
    wire N__3978;
    wire N__3975;
    wire N__3972;
    wire N__3969;
    wire N__3968;
    wire N__3967;
    wire N__3964;
    wire N__3961;
    wire N__3960;
    wire N__3957;
    wire N__3950;
    wire N__3945;
    wire N__3944;
    wire N__3939;
    wire N__3936;
    wire N__3935;
    wire N__3934;
    wire N__3931;
    wire N__3928;
    wire N__3925;
    wire N__3918;
    wire N__3917;
    wire N__3914;
    wire N__3913;
    wire N__3912;
    wire N__3909;
    wire N__3904;
    wire N__3901;
    wire N__3898;
    wire N__3891;
    wire N__3888;
    wire N__3887;
    wire N__3884;
    wire N__3881;
    wire N__3876;
    wire N__3873;
    wire N__3870;
    wire N__3869;
    wire N__3866;
    wire N__3863;
    wire N__3860;
    wire N__3855;
    wire N__3852;
    wire N__3849;
    wire N__3846;
    wire N__3843;
    wire N__3840;
    wire N__3837;
    wire N__3836;
    wire N__3833;
    wire N__3830;
    wire N__3827;
    wire N__3822;
    wire N__3821;
    wire N__3820;
    wire N__3813;
    wire N__3810;
    wire N__3809;
    wire N__3806;
    wire N__3803;
    wire N__3798;
    wire N__3797;
    wire N__3794;
    wire N__3791;
    wire N__3786;
    wire N__3783;
    wire N__3782;
    wire N__3779;
    wire N__3776;
    wire N__3771;
    wire N__3768;
    wire N__3765;
    wire N__3762;
    wire N__3761;
    wire N__3758;
    wire N__3755;
    wire N__3750;
    wire N__3747;
    wire N__3746;
    wire N__3743;
    wire N__3740;
    wire N__3735;
    wire N__3732;
    wire N__3729;
    wire N__3726;
    wire N__3723;
    wire N__3720;
    wire N__3719;
    wire N__3716;
    wire N__3713;
    wire N__3708;
    wire N__3705;
    wire N__3702;
    wire N__3699;
    wire N__3696;
    wire N__3693;
    wire N__3690;
    wire N__3687;
    wire N__3684;
    wire N__3681;
    wire N__3680;
    wire N__3677;
    wire N__3674;
    wire N__3669;
    wire N__3666;
    wire N__3665;
    wire N__3664;
    wire N__3663;
    wire N__3662;
    wire N__3659;
    wire N__3656;
    wire N__3649;
    wire N__3642;
    wire N__3641;
    wire N__3638;
    wire N__3635;
    wire N__3630;
    wire N__3629;
    wire N__3626;
    wire N__3623;
    wire N__3620;
    wire N__3619;
    wire N__3618;
    wire N__3615;
    wire N__3612;
    wire N__3607;
    wire N__3600;
    wire N__3597;
    wire N__3594;
    wire N__3591;
    wire N__3588;
    wire N__3585;
    wire N__3582;
    wire N__3579;
    wire N__3578;
    wire N__3575;
    wire N__3572;
    wire N__3567;
    wire N__3566;
    wire N__3563;
    wire N__3560;
    wire N__3555;
    wire N__3554;
    wire N__3553;
    wire N__3546;
    wire N__3543;
    wire N__3540;
    wire N__3539;
    wire N__3536;
    wire N__3533;
    wire N__3528;
    wire N__3525;
    wire N__3524;
    wire N__3523;
    wire N__3516;
    wire N__3513;
    wire N__3512;
    wire N__3509;
    wire N__3506;
    wire N__3501;
    wire N__3498;
    wire N__3495;
    wire N__3492;
    wire N__3489;
    wire N__3486;
    wire N__3483;
    wire N__3480;
    wire N__3477;
    wire N__3474;
    wire N__3473;
    wire N__3468;
    wire N__3465;
    wire N__3462;
    wire N__3459;
    wire N__3456;
    wire N__3455;
    wire N__3454;
    wire N__3453;
    wire N__3450;
    wire N__3447;
    wire N__3442;
    wire N__3435;
    wire N__3432;
    wire N__3431;
    wire N__3430;
    wire N__3427;
    wire N__3424;
    wire N__3421;
    wire N__3414;
    wire N__3411;
    wire N__3408;
    wire N__3405;
    wire N__3404;
    wire N__3401;
    wire N__3398;
    wire N__3393;
    wire N__3390;
    wire N__3387;
    wire N__3386;
    wire N__3383;
    wire N__3380;
    wire N__3379;
    wire N__3376;
    wire N__3373;
    wire N__3370;
    wire N__3363;
    wire N__3360;
    wire N__3357;
    wire N__3356;
    wire N__3353;
    wire N__3350;
    wire N__3349;
    wire N__3346;
    wire N__3343;
    wire N__3340;
    wire N__3337;
    wire N__3332;
    wire N__3327;
    wire N__3324;
    wire N__3321;
    wire N__3318;
    wire N__3317;
    wire N__3316;
    wire N__3313;
    wire N__3308;
    wire N__3303;
    wire N__3300;
    wire N__3297;
    wire N__3294;
    wire N__3291;
    wire N__3290;
    wire N__3287;
    wire N__3286;
    wire N__3285;
    wire N__3284;
    wire N__3281;
    wire N__3272;
    wire N__3267;
    wire N__3266;
    wire N__3265;
    wire N__3264;
    wire N__3255;
    wire N__3252;
    wire N__3249;
    wire N__3246;
    wire N__3245;
    wire N__3244;
    wire N__3241;
    wire N__3238;
    wire N__3235;
    wire N__3228;
    wire N__3227;
    wire N__3226;
    wire N__3225;
    wire N__3222;
    wire N__3219;
    wire N__3214;
    wire N__3213;
    wire N__3206;
    wire N__3203;
    wire N__3200;
    wire N__3197;
    wire N__3192;
    wire N__3191;
    wire N__3188;
    wire N__3185;
    wire N__3180;
    wire N__3177;
    wire N__3174;
    wire N__3171;
    wire N__3168;
    wire N__3165;
    wire N__3162;
    wire N__3159;
    wire N__3156;
    wire N__3153;
    wire N__3150;
    wire N__3147;
    wire N__3144;
    wire N__3141;
    wire N__3140;
    wire N__3139;
    wire N__3138;
    wire N__3131;
    wire N__3130;
    wire N__3129;
    wire N__3126;
    wire N__3123;
    wire N__3120;
    wire N__3117;
    wire N__3114;
    wire N__3111;
    wire N__3106;
    wire N__3103;
    wire N__3098;
    wire N__3095;
    wire N__3092;
    wire N__3087;
    wire N__3086;
    wire N__3081;
    wire N__3078;
    wire N__3075;
    wire N__3072;
    wire N__3069;
    wire N__3066;
    wire N__3063;
    wire N__3060;
    wire N__3057;
    wire N__3054;
    wire N__3051;
    wire N__3048;
    wire N__3045;
    wire N__3042;
    wire N__3039;
    wire N__3036;
    wire N__3033;
    wire N__3030;
    wire N__3027;
    wire N__3024;
    wire N__3021;
    wire N__3018;
    wire N__3015;
    wire N__3012;
    wire N__3009;
    wire N__3008;
    wire N__3007;
    wire N__3004;
    wire N__3001;
    wire N__2998;
    wire N__2993;
    wire N__2990;
    wire N__2985;
    wire N__2982;
    wire N__2979;
    wire N__2978;
    wire N__2975;
    wire N__2972;
    wire N__2971;
    wire N__2966;
    wire N__2963;
    wire N__2960;
    wire N__2957;
    wire N__2954;
    wire N__2951;
    wire N__2948;
    wire N__2945;
    wire N__2942;
    wire N__2939;
    wire N__2934;
    wire N__2931;
    wire N__2928;
    wire N__2925;
    wire N__2922;
    wire N__2919;
    wire N__2916;
    wire N__2913;
    wire N__2910;
    wire N__2907;
    wire N__2904;
    wire N__2901;
    wire N__2898;
    wire N__2895;
    wire N__2892;
    wire N__2889;
    wire N__2886;
    wire N__2883;
    wire N__2880;
    wire N__2877;
    wire N__2874;
    wire N__2871;
    wire N__2868;
    wire N__2865;
    wire N__2862;
    wire N__2859;
    wire N__2856;
    wire N__2855;
    wire N__2850;
    wire N__2847;
    wire N__2844;
    wire N__2841;
    wire N__2838;
    wire N__2837;
    wire N__2832;
    wire N__2829;
    wire N__2826;
    wire N__2823;
    wire N__2820;
    wire N__2817;
    wire N__2814;
    wire N__2813;
    wire N__2810;
    wire N__2807;
    wire N__2804;
    wire N__2801;
    wire N__2798;
    wire N__2795;
    wire N__2790;
    wire N__2787;
    wire N__2784;
    wire N__2781;
    wire N__2778;
    wire N__2777;
    wire N__2772;
    wire N__2769;
    wire N__2766;
    wire N__2763;
    wire N__2760;
    wire N__2759;
    wire N__2754;
    wire N__2751;
    wire N__2748;
    wire N__2745;
    wire N__2742;
    wire N__2739;
    wire N__2736;
    wire N__2735;
    wire N__2730;
    wire N__2727;
    wire N__2724;
    wire N__2721;
    wire N__2718;
    wire N__2717;
    wire N__2712;
    wire N__2709;
    wire N__2706;
    wire N__2703;
    wire N__2700;
    wire N__2697;
    wire N__2694;
    wire N__2693;
    wire N__2690;
    wire N__2685;
    wire N__2682;
    wire N__2679;
    wire N__2676;
    wire N__2673;
    wire N__2670;
    wire N__2667;
    wire N__2666;
    wire N__2665;
    wire N__2664;
    wire N__2661;
    wire N__2656;
    wire N__2653;
    wire N__2652;
    wire N__2645;
    wire N__2642;
    wire N__2637;
    wire N__2634;
    wire N__2631;
    wire N__2628;
    wire N__2625;
    wire N__2622;
    wire N__2619;
    wire N__2616;
    wire N__2615;
    wire N__2614;
    wire N__2611;
    wire N__2606;
    wire N__2603;
    wire N__2600;
    wire N__2597;
    wire N__2594;
    wire N__2589;
    wire N__2586;
    wire N__2583;
    wire N__2580;
    wire N__2577;
    wire N__2574;
    wire N__2571;
    wire N__2568;
    wire N__2567;
    wire N__2562;
    wire N__2559;
    wire N__2556;
    wire N__2553;
    wire N__2550;
    wire N__2547;
    wire N__2544;
    wire N__2543;
    wire N__2540;
    wire N__2537;
    wire N__2532;
    wire N__2529;
    wire N__2526;
    wire N__2523;
    wire N__2520;
    wire N__2517;
    wire N__2514;
    wire N__2511;
    wire N__2508;
    wire N__2507;
    wire N__2504;
    wire N__2501;
    wire N__2498;
    wire N__2495;
    wire N__2490;
    wire N__2487;
    wire N__2484;
    wire N__2481;
    wire N__2480;
    wire N__2475;
    wire N__2472;
    wire N__2469;
    wire N__2466;
    wire N__2465;
    wire N__2462;
    wire N__2459;
    wire N__2458;
    wire N__2455;
    wire N__2450;
    wire N__2445;
    wire N__2442;
    wire N__2439;
    wire N__2436;
    wire N__2433;
    wire N__2432;
    wire N__2431;
    wire N__2430;
    wire N__2423;
    wire N__2420;
    wire N__2415;
    wire N__2412;
    wire N__2409;
    wire N__2406;
    wire N__2405;
    wire N__2404;
    wire N__2403;
    wire N__2402;
    wire N__2401;
    wire N__2400;
    wire N__2399;
    wire N__2398;
    wire N__2397;
    wire N__2396;
    wire N__2373;
    wire CLK80_OUT;
    wire GNDG0;
    wire VCCG0;
    wire A_c_18;
    wire A_c_16;
    wire \U409_CIA.g0Z0Z_11 ;
    wire A_c_17;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2_cascade_ ;
    wire \U409_ADDRESS_DECODE.CIA_SPACEm_6 ;
    wire A_c_20;
    wire \U409_CIA.g0Z0Z_8 ;
    wire A_c_21;
    wire A_c_29;
    wire A_c_30;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3 ;
    wire A_c_25;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4 ;
    wire A_c_27;
    wire A_c_26;
    wire A_c_24;
    wire A_c_31;
    wire \U409_CIA.g0Z0Z_2 ;
    wire A_c_28;
    wire \U409_CIA.g0Z0Z_10_cascade_ ;
    wire A_c_22;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2 ;
    wire A_c_19;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3 ;
    wire \U409_ADDRESS_DECODE.un1_REGSPACEnZ0_cascade_ ;
    wire PORTSIZE_0_i;
    wire A_c_23;
    wire \U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_3 ;
    wire U409_ADDRESS_DECODE_un1_REGSPACEn_i;
    wire U409_ADDRESS_DECODE_un1_RAMSPACEn_i;
    wire \U409_ADDRESS_DECODE.un10_ROMENZ0 ;
    wire \U409_ADDRESS_DECODE.un1_REGSPACEnZ0 ;
    wire \U409_ADDRESS_DECODE.un6_ROMENZ0 ;
    wire OVL_c;
    wire A_c_13;
    wire U409_ADDRESS_DECODE_un1_CIACS1n_i;
    wire A_c_12;
    wire U409_ADDRESS_DECODE_un1_CIACS0n_i;
    wire \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ;
    wire \U409_TRANSFER_ACK.RESETn_c_i ;
    wire CIA_ENABLEm;
    wire \U409_CIA.g0Z0Z_14 ;
    wire \U409_CIA.g0Z0Z_13 ;
    wire \U409_CIA.CIA_HOLDZ0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_3_0_cascade_ ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ;
    wire \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa ;
    wire U409_ADDRESS_DECODE_Z2_SPACE;
    wire U409_ADDRESS_DECODE_un1_ROMEN_0;
    wire ROMENm_i;
    wire \U409_TRANSFER_ACK.m9_bm_cascade_ ;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_0C_net ;
    wire \U409_TRANSFER_ACK.N_4_cascade_ ;
    wire \U409_TRANSFER_ACK.m9_am ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_1 ;
    wire \U409_TRANSFER_ACK.N_4 ;
    wire \U409_TRANSFER_ACK.i6_mux_0_cascade_ ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.LASTCLK_1C_net ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ;
    wire \U409_TRANSFER_ACK.N_97 ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_TACK_EN_0_cascade_ ;
    wire \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ;
    wire TACK_OUTn;
    wire \U409_TRANSFER_ACK.CIA_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_ ;
    wire \U409_TRANSFER_ACK.ROM_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_ ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ;
    wire \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ;
    wire \INVU409_TRANSFER_ACK.TACK_EN_iC_net ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0 ;
    wire \U409_TICK.TICK603_11_cascade_ ;
    wire \U409_TICK.TICK603_14_cascade_ ;
    wire \U409_TICK.TICK603_8 ;
    wire bfn_10_6_0_;
    wire \U409_TICK.COUNTER60Z0Z_2 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_1 ;
    wire \U409_TICK.COUNTER60Z0Z_3 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_2 ;
    wire \U409_TICK.COUNTER60Z0Z_4 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_4 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_3 ;
    wire \U409_TICK.COUNTER60Z0Z_5 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_4 ;
    wire \U409_TICK.COUNTER60Z0Z_6 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_6 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_5 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_6 ;
    wire \U409_TICK.COUNTER60Z0Z_8 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_8 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_8 ;
    wire bfn_10_7_0_;
    wire \U409_TICK.un3_COUNTER60_1_cry_9 ;
    wire \U409_TICK.COUNTER60Z0Z_11 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_10 ;
    wire \U409_TICK.COUNTER60Z0Z_12 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_11 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_12 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_13 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_15 ;
    wire \U409_TICK.COUNTER60Z0Z_16 ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_0 ;
    wire \INVU409_TRANSFER_ACK.LASTCLK_0C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ;
    wire \U409_TICK.COUNTER60Z0Z_1 ;
    wire \U409_TICK.COUNTER60Z0Z_0 ;
    wire TICK60_c;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_15 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_9 ;
    wire \U409_TICK.COUNTER60Z0Z_9 ;
    wire \U409_TICK.COUNTER60Z0Z_13 ;
    wire \U409_TICK.COUNTER60Z0Z_10 ;
    wire \U409_TICK.COUNTER60Z0Z_7 ;
    wire \U409_TICK.COUNTER60Z0Z_15 ;
    wire \U409_TICK.TICK603_10 ;
    wire \U409_TICK.TICK603_9 ;
    wire \U409_TICK.TICK603_14 ;
    wire \U409_TICK.TICK603_10_cascade_ ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_14 ;
    wire \U409_TICK.COUNTER60Z0Z_14 ;
    wire \U409_TICK.TICK503_11 ;
    wire \U409_TICK.TICK503_8_cascade_ ;
    wire \U409_TICK.TICK503_14_cascade_ ;
    wire \U409_TICK.TICK503_10_cascade_ ;
    wire \U409_TICK.TICK503_9_cascade_ ;
    wire \U409_TICK.TICK503_14 ;
    wire \U409_TICK.TICK503_10 ;
    wire \U409_TICK.TICK503_9 ;
    wire TICK50_c;
    wire \U409_CIA.N_9_cascade_ ;
    wire \U409_CIA.VMAZ0 ;
    wire \U409_CIA.N_20_cascade_ ;
    wire \U409_CIA.CLKCIA6_0_a2_1 ;
    wire \U409_CIA.CLKCIAZ0_cascade_ ;
    wire CLKCIA_c;
    wire \U409_CIA.CLKCIA8_0_a2_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ;
    wire CLK40_IN_c;
    wire TSn_c;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ;
    wire CONSTANT_ONE_NET;
    wire \U409_TICK.COUNTER50Z0Z_1 ;
    wire \U409_TICK.COUNTER50Z0Z_0 ;
    wire bfn_12_6_0_;
    wire \U409_TICK.COUNTER50Z0Z_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_1 ;
    wire \U409_TICK.COUNTER50Z0Z_3 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_2 ;
    wire \U409_TICK.COUNTER50Z0Z_4 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_3 ;
    wire \U409_TICK.COUNTER50Z0Z_5 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_5 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_4 ;
    wire \U409_TICK.COUNTER50Z0Z_6 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_6 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_5 ;
    wire \U409_TICK.COUNTER50Z0Z_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_6 ;
    wire \U409_TICK.COUNTER50Z0Z_8 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_8 ;
    wire \U409_TICK.COUNTER50Z0Z_9 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_9 ;
    wire bfn_12_7_0_;
    wire \U409_TICK.COUNTER50Z0Z_10 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_9 ;
    wire \U409_TICK.COUNTER50Z0Z_11 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_11 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_10 ;
    wire \U409_TICK.COUNTER50Z0Z_12 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_11 ;
    wire \U409_TICK.COUNTER50Z0Z_13 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_13 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_12 ;
    wire \U409_TICK.COUNTER50Z0Z_14 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_13 ;
    wire \U409_TICK.COUNTER50Z0Z_15 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_15 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_15 ;
    wire \U409_TICK.COUNTER50Z0Z_16 ;
    wire CLK6_c_g;
    wire bfn_12_9_0_;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_1 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_3 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4 ;
    wire \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_2 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_1 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_4 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_5 ;
    wire \U409_CIA.CIA_CLK_COUNT11_0_a2_2 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ;
    wire \U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_0 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_3 ;
    wire CLK28_IN_c_g;
    wire TACK_EN_i;
    wire N_353_i;
    wire BUFENn_c;
    wire TACKn_in;
    wire RESETn_c;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="SIMPLE";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0001111;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE pll (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__4692),
            .RESETB(N__4977),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(CLK80_OUT));
    PRE_IO_GBUF CLK28_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__6077),
            .GLOBALBUFFEROUTPUT(CLK28_IN_c_g));
    IO_PAD CLK28_IN_ibuf_gb_io_iopad (
            .OE(N__6079),
            .DIN(N__6078),
            .DOUT(N__6077),
            .PACKAGEPIN(CLK28_IN));
    defparam CLK28_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK28_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK28_IN_ibuf_gb_io_preio (
            .PADOEN(N__6079),
            .PADOUT(N__6078),
            .PADIN(N__6077),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK6_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__6067),
            .GLOBALBUFFEROUTPUT(CLK6_c_g));
    IO_PAD CLK6_ibuf_gb_io_iopad (
            .OE(N__6069),
            .DIN(N__6068),
            .DOUT(N__6067),
            .PACKAGEPIN(CLK6));
    defparam CLK6_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK6_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK6_ibuf_gb_io_preio (
            .PADOEN(N__6069),
            .PADOUT(N__6068),
            .PADIN(N__6067),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKCIA_obuf_iopad (
            .OE(N__6058),
            .DIN(N__6057),
            .DOUT(N__6056),
            .PACKAGEPIN(CLKCIA));
    defparam CLKCIA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKCIA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKCIA_obuf_preio (
            .PADOEN(N__6058),
            .PADOUT(N__6057),
            .PADIN(N__6056),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4275),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_23_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_23_iopad (
            .OE(N__6049),
            .DIN(N__6048),
            .DOUT(N__6047),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__6049),
            .PADOUT(N__6048),
            .PADIN(N__6047),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_24_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_24_iopad (
            .OE(N__6040),
            .DIN(N__6039),
            .DOUT(N__6038),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__6040),
            .PADOUT(N__6039),
            .PADIN(N__6038),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_31_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_31_iopad (
            .OE(N__6031),
            .DIN(N__6030),
            .DOUT(N__6029),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__6031),
            .PADOUT(N__6030),
            .PADIN(N__6029),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS1n_obuf_iopad (
            .OE(N__6022),
            .DIN(N__6021),
            .DOUT(N__6020),
            .PACKAGEPIN(CIACS1n));
    defparam CIACS1n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS1n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS1n_obuf_preio (
            .PADOEN(N__6022),
            .PADOUT(N__6021),
            .PADIN(N__6020),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2916),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_obuf_iopad (
            .OE(N__6013),
            .DIN(N__6012),
            .DOUT(N__6011),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGSPACEn_obuf_preio (
            .PADOEN(N__6013),
            .PADOUT(N__6012),
            .PADIN(N__6011),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3072),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_17_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_17_iopad (
            .OE(N__6004),
            .DIN(N__6003),
            .DOUT(N__6002),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__6004),
            .PADOUT(N__6003),
            .PADIN(N__6002),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_21_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_21_iopad (
            .OE(N__5995),
            .DIN(N__5994),
            .DOUT(N__5993),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__5995),
            .PADOUT(N__5994),
            .PADIN(N__5993),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_obuf_iopad (
            .OE(N__5986),
            .DIN(N__5985),
            .DOUT(N__5984),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMSPACEn_obuf_preio (
            .PADOEN(N__5986),
            .PADOUT(N__5985),
            .PADIN(N__5984),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3048),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TACKn_iobuf_iopad.PULLUP=1'b1;
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__5977),
            .DIN(N__5976),
            .DOUT(N__5975),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__5977),
            .PADOUT(N__5976),
            .PADIN(N__5975),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5610),
            .DIN0(TACKn_in),
            .DOUT0(N__3597),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_12_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_12_iopad (
            .OE(N__5968),
            .DIN(N__5967),
            .DOUT(N__5966),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__5968),
            .PADOUT(N__5967),
            .PADIN(N__5966),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ROMENn_obuf_iopad (
            .OE(N__5959),
            .DIN(N__5958),
            .DOUT(N__5957),
            .PACKAGEPIN(ROMENn));
    defparam ROMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ROMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ROMENn_obuf_preio (
            .PADOEN(N__5959),
            .PADOUT(N__5958),
            .PADIN(N__5957),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3180),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__5950),
            .DIN(N__5949),
            .DOUT(N__5948),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__5950),
            .PADOUT(N__5949),
            .PADIN(N__5948),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__5941),
            .DIN(N__5940),
            .DOUT(N__5939),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__5941),
            .PADOUT(N__5940),
            .PADIN(N__5939),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5586),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam PORTSIZE_obuf_iopad.PULLUP=1'b1;
    IO_PAD PORTSIZE_obuf_iopad (
            .OE(N__5932),
            .DIN(N__5931),
            .DOUT(N__5930),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PORTSIZE_obuf_preio (
            .PADOEN(N__5932),
            .PADOUT(N__5931),
            .PADIN(N__5930),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3162),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_18_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_18_iopad (
            .OE(N__5923),
            .DIN(N__5922),
            .DOUT(N__5921),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__5923),
            .PADOUT(N__5922),
            .PADIN(N__5921),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_29_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_29_iopad (
            .OE(N__5914),
            .DIN(N__5913),
            .DOUT(N__5912),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__5914),
            .PADOUT(N__5913),
            .PADIN(N__5912),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_22_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_22_iopad (
            .OE(N__5905),
            .DIN(N__5904),
            .DOUT(N__5903),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__5905),
            .PADOUT(N__5904),
            .PADIN(N__5903),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_27_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_27_iopad (
            .OE(N__5896),
            .DIN(N__5895),
            .DOUT(N__5894),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__5896),
            .PADOUT(N__5895),
            .PADIN(N__5894),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__5887),
            .DIN(N__5886),
            .DOUT(N__5885),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__5887),
            .PADOUT(N__5886),
            .PADIN(N__5885),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__5878),
            .DIN(N__5877),
            .DOUT(N__5876),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__5878),
            .PADOUT(N__5877),
            .PADIN(N__5876),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_20_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_20_iopad (
            .OE(N__5869),
            .DIN(N__5868),
            .DOUT(N__5867),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__5869),
            .PADOUT(N__5868),
            .PADIN(N__5867),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_13_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_13_iopad (
            .OE(N__5860),
            .DIN(N__5859),
            .DOUT(N__5858),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__5860),
            .PADOUT(N__5859),
            .PADIN(N__5858),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_25_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_25_iopad (
            .OE(N__5851),
            .DIN(N__5850),
            .DOUT(N__5849),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__5851),
            .PADOUT(N__5850),
            .PADIN(N__5849),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS0n_obuf_iopad (
            .OE(N__5842),
            .DIN(N__5841),
            .DOUT(N__5840),
            .PACKAGEPIN(CIACS0n));
    defparam CIACS0n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS0n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS0n_obuf_preio (
            .PADOEN(N__5842),
            .PADOUT(N__5841),
            .PADIN(N__5840),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2880),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK50_obuf_iopad (
            .OE(N__5833),
            .DIN(N__5832),
            .DOUT(N__5831),
            .PACKAGEPIN(TICK50));
    defparam TICK50_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK50_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK50_obuf_preio (
            .PADOEN(N__5833),
            .PADOUT(N__5832),
            .PADIN(N__5831),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4350),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_19_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_19_iopad (
            .OE(N__5824),
            .DIN(N__5823),
            .DOUT(N__5822),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__5824),
            .PADOUT(N__5823),
            .PADIN(N__5822),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_28_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_28_iopad (
            .OE(N__5815),
            .DIN(N__5814),
            .DOUT(N__5813),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__5815),
            .PADOUT(N__5814),
            .PADIN(N__5813),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_30_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_30_iopad (
            .OE(N__5806),
            .DIN(N__5805),
            .DOUT(N__5804),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__5806),
            .PADOUT(N__5805),
            .PADIN(N__5804),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD OVL_ibuf_iopad (
            .OE(N__5797),
            .DIN(N__5796),
            .DOUT(N__5795),
            .PACKAGEPIN(OVL));
    defparam OVL_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam OVL_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO OVL_ibuf_preio (
            .PADOEN(N__5797),
            .PADOUT(N__5796),
            .PADIN(N__5795),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(OVL_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_16_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_16_iopad (
            .OE(N__5788),
            .DIN(N__5787),
            .DOUT(N__5786),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__5788),
            .PADOUT(N__5787),
            .PADIN(N__5786),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK60_obuf_iopad (
            .OE(N__5779),
            .DIN(N__5778),
            .DOUT(N__5777),
            .PACKAGEPIN(TICK60));
    defparam TICK60_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK60_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK60_obuf_preio (
            .PADOEN(N__5779),
            .PADOUT(N__5778),
            .PADIN(N__5777),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4209),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_26_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_26_iopad (
            .OE(N__5770),
            .DIN(N__5769),
            .DOUT(N__5768),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__5770),
            .PADOUT(N__5769),
            .PADIN(N__5768),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__1333 (
            .O(N__5751),
            .I(N__5746));
    InMux I__1332 (
            .O(N__5750),
            .I(N__5740));
    InMux I__1331 (
            .O(N__5749),
            .I(N__5740));
    InMux I__1330 (
            .O(N__5746),
            .I(N__5737));
    InMux I__1329 (
            .O(N__5745),
            .I(N__5734));
    LocalMux I__1328 (
            .O(N__5740),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__1327 (
            .O(N__5737),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__1326 (
            .O(N__5734),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    InMux I__1325 (
            .O(N__5727),
            .I(N__5724));
    LocalMux I__1324 (
            .O(N__5724),
            .I(\U409_CIA.CIA_CLK_COUNT11_0_a2_2 ));
    InMux I__1323 (
            .O(N__5721),
            .I(N__5718));
    LocalMux I__1322 (
            .O(N__5718),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ));
    CascadeMux I__1321 (
            .O(N__5715),
            .I(\U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_ ));
    CascadeMux I__1320 (
            .O(N__5712),
            .I(N__5702));
    InMux I__1319 (
            .O(N__5711),
            .I(N__5699));
    InMux I__1318 (
            .O(N__5710),
            .I(N__5696));
    InMux I__1317 (
            .O(N__5709),
            .I(N__5689));
    InMux I__1316 (
            .O(N__5708),
            .I(N__5689));
    InMux I__1315 (
            .O(N__5707),
            .I(N__5689));
    InMux I__1314 (
            .O(N__5706),
            .I(N__5682));
    InMux I__1313 (
            .O(N__5705),
            .I(N__5682));
    InMux I__1312 (
            .O(N__5702),
            .I(N__5682));
    LocalMux I__1311 (
            .O(N__5699),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1310 (
            .O(N__5696),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1309 (
            .O(N__5689),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1308 (
            .O(N__5682),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    InMux I__1307 (
            .O(N__5673),
            .I(N__5664));
    InMux I__1306 (
            .O(N__5672),
            .I(N__5657));
    InMux I__1305 (
            .O(N__5671),
            .I(N__5657));
    InMux I__1304 (
            .O(N__5670),
            .I(N__5657));
    InMux I__1303 (
            .O(N__5669),
            .I(N__5650));
    InMux I__1302 (
            .O(N__5668),
            .I(N__5650));
    InMux I__1301 (
            .O(N__5667),
            .I(N__5650));
    LocalMux I__1300 (
            .O(N__5664),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__1299 (
            .O(N__5657),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__1298 (
            .O(N__5650),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    ClkMux I__1297 (
            .O(N__5643),
            .I(N__5631));
    ClkMux I__1296 (
            .O(N__5642),
            .I(N__5631));
    ClkMux I__1295 (
            .O(N__5641),
            .I(N__5631));
    ClkMux I__1294 (
            .O(N__5640),
            .I(N__5631));
    GlobalMux I__1293 (
            .O(N__5631),
            .I(N__5628));
    gio2CtrlBuf I__1292 (
            .O(N__5628),
            .I(CLK28_IN_c_g));
    InMux I__1291 (
            .O(N__5625),
            .I(N__5622));
    LocalMux I__1290 (
            .O(N__5622),
            .I(N__5619));
    Span4Mux_v I__1289 (
            .O(N__5619),
            .I(N__5616));
    Sp12to4 I__1288 (
            .O(N__5616),
            .I(N__5613));
    Odrv12 I__1287 (
            .O(N__5613),
            .I(TACK_EN_i));
    IoInMux I__1286 (
            .O(N__5610),
            .I(N__5607));
    LocalMux I__1285 (
            .O(N__5607),
            .I(N__5604));
    IoSpan4Mux I__1284 (
            .O(N__5604),
            .I(N__5601));
    Span4Mux_s1_v I__1283 (
            .O(N__5601),
            .I(N__5598));
    Span4Mux_v I__1282 (
            .O(N__5598),
            .I(N__5595));
    Span4Mux_v I__1281 (
            .O(N__5595),
            .I(N__5592));
    Span4Mux_v I__1280 (
            .O(N__5592),
            .I(N__5589));
    Odrv4 I__1279 (
            .O(N__5589),
            .I(N_353_i));
    IoInMux I__1278 (
            .O(N__5586),
            .I(N__5583));
    LocalMux I__1277 (
            .O(N__5583),
            .I(N__5580));
    Span4Mux_s1_v I__1276 (
            .O(N__5580),
            .I(N__5577));
    Sp12to4 I__1275 (
            .O(N__5577),
            .I(N__5573));
    InMux I__1274 (
            .O(N__5576),
            .I(N__5570));
    Span12Mux_h I__1273 (
            .O(N__5573),
            .I(N__5567));
    LocalMux I__1272 (
            .O(N__5570),
            .I(N__5564));
    Span12Mux_v I__1271 (
            .O(N__5567),
            .I(N__5559));
    Span12Mux_h I__1270 (
            .O(N__5564),
            .I(N__5559));
    Odrv12 I__1269 (
            .O(N__5559),
            .I(BUFENn_c));
    InMux I__1268 (
            .O(N__5556),
            .I(N__5553));
    LocalMux I__1267 (
            .O(N__5553),
            .I(N__5550));
    Span12Mux_h I__1266 (
            .O(N__5550),
            .I(N__5547));
    Span12Mux_v I__1265 (
            .O(N__5547),
            .I(N__5544));
    Odrv12 I__1264 (
            .O(N__5544),
            .I(TACKn_in));
    InMux I__1263 (
            .O(N__5541),
            .I(N__5538));
    LocalMux I__1262 (
            .O(N__5538),
            .I(N__5534));
    InMux I__1261 (
            .O(N__5537),
            .I(N__5530));
    Span4Mux_v I__1260 (
            .O(N__5534),
            .I(N__5526));
    CascadeMux I__1259 (
            .O(N__5533),
            .I(N__5517));
    LocalMux I__1258 (
            .O(N__5530),
            .I(N__5508));
    InMux I__1257 (
            .O(N__5529),
            .I(N__5505));
    Span4Mux_h I__1256 (
            .O(N__5526),
            .I(N__5501));
    InMux I__1255 (
            .O(N__5525),
            .I(N__5492));
    InMux I__1254 (
            .O(N__5524),
            .I(N__5492));
    InMux I__1253 (
            .O(N__5523),
            .I(N__5492));
    InMux I__1252 (
            .O(N__5522),
            .I(N__5492));
    InMux I__1251 (
            .O(N__5521),
            .I(N__5489));
    InMux I__1250 (
            .O(N__5520),
            .I(N__5486));
    InMux I__1249 (
            .O(N__5517),
            .I(N__5479));
    InMux I__1248 (
            .O(N__5516),
            .I(N__5479));
    InMux I__1247 (
            .O(N__5515),
            .I(N__5479));
    InMux I__1246 (
            .O(N__5514),
            .I(N__5476));
    InMux I__1245 (
            .O(N__5513),
            .I(N__5469));
    InMux I__1244 (
            .O(N__5512),
            .I(N__5469));
    InMux I__1243 (
            .O(N__5511),
            .I(N__5469));
    Span4Mux_h I__1242 (
            .O(N__5508),
            .I(N__5463));
    LocalMux I__1241 (
            .O(N__5505),
            .I(N__5463));
    InMux I__1240 (
            .O(N__5504),
            .I(N__5460));
    Span4Mux_h I__1239 (
            .O(N__5501),
            .I(N__5444));
    LocalMux I__1238 (
            .O(N__5492),
            .I(N__5444));
    LocalMux I__1237 (
            .O(N__5489),
            .I(N__5444));
    LocalMux I__1236 (
            .O(N__5486),
            .I(N__5444));
    LocalMux I__1235 (
            .O(N__5479),
            .I(N__5444));
    LocalMux I__1234 (
            .O(N__5476),
            .I(N__5444));
    LocalMux I__1233 (
            .O(N__5469),
            .I(N__5444));
    InMux I__1232 (
            .O(N__5468),
            .I(N__5441));
    Span4Mux_v I__1231 (
            .O(N__5463),
            .I(N__5436));
    LocalMux I__1230 (
            .O(N__5460),
            .I(N__5436));
    InMux I__1229 (
            .O(N__5459),
            .I(N__5432));
    Span4Mux_v I__1228 (
            .O(N__5444),
            .I(N__5429));
    LocalMux I__1227 (
            .O(N__5441),
            .I(N__5426));
    Span4Mux_v I__1226 (
            .O(N__5436),
            .I(N__5423));
    InMux I__1225 (
            .O(N__5435),
            .I(N__5420));
    LocalMux I__1224 (
            .O(N__5432),
            .I(N__5417));
    Span4Mux_h I__1223 (
            .O(N__5429),
            .I(N__5414));
    Span4Mux_v I__1222 (
            .O(N__5426),
            .I(N__5411));
    Span4Mux_h I__1221 (
            .O(N__5423),
            .I(N__5408));
    LocalMux I__1220 (
            .O(N__5420),
            .I(N__5405));
    Span4Mux_h I__1219 (
            .O(N__5417),
            .I(N__5402));
    Sp12to4 I__1218 (
            .O(N__5414),
            .I(N__5397));
    Sp12to4 I__1217 (
            .O(N__5411),
            .I(N__5397));
    Sp12to4 I__1216 (
            .O(N__5408),
            .I(N__5392));
    Span12Mux_h I__1215 (
            .O(N__5405),
            .I(N__5392));
    Span4Mux_h I__1214 (
            .O(N__5402),
            .I(N__5389));
    Span12Mux_h I__1213 (
            .O(N__5397),
            .I(N__5386));
    Span12Mux_v I__1212 (
            .O(N__5392),
            .I(N__5383));
    Sp12to4 I__1211 (
            .O(N__5389),
            .I(N__5380));
    Span12Mux_v I__1210 (
            .O(N__5386),
            .I(N__5375));
    Span12Mux_h I__1209 (
            .O(N__5383),
            .I(N__5375));
    Span12Mux_v I__1208 (
            .O(N__5380),
            .I(N__5372));
    Odrv12 I__1207 (
            .O(N__5375),
            .I(RESETn_c));
    Odrv12 I__1206 (
            .O(N__5372),
            .I(RESETn_c));
    SRMux I__1205 (
            .O(N__5367),
            .I(N__5362));
    SRMux I__1204 (
            .O(N__5366),
            .I(N__5359));
    SRMux I__1203 (
            .O(N__5365),
            .I(N__5356));
    LocalMux I__1202 (
            .O(N__5362),
            .I(N__5353));
    LocalMux I__1201 (
            .O(N__5359),
            .I(N__5350));
    LocalMux I__1200 (
            .O(N__5356),
            .I(N__5347));
    Span4Mux_v I__1199 (
            .O(N__5353),
            .I(N__5344));
    Span4Mux_h I__1198 (
            .O(N__5350),
            .I(N__5341));
    Span4Mux_v I__1197 (
            .O(N__5347),
            .I(N__5338));
    Sp12to4 I__1196 (
            .O(N__5344),
            .I(N__5335));
    Span4Mux_h I__1195 (
            .O(N__5341),
            .I(N__5332));
    Span4Mux_h I__1194 (
            .O(N__5338),
            .I(N__5329));
    Odrv12 I__1193 (
            .O(N__5335),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    Odrv4 I__1192 (
            .O(N__5332),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    Odrv4 I__1191 (
            .O(N__5329),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    InMux I__1190 (
            .O(N__5322),
            .I(\U409_TICK.un2_COUNTER50_1_cry_15 ));
    InMux I__1189 (
            .O(N__5319),
            .I(N__5315));
    InMux I__1188 (
            .O(N__5318),
            .I(N__5312));
    LocalMux I__1187 (
            .O(N__5315),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    LocalMux I__1186 (
            .O(N__5312),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    ClkMux I__1185 (
            .O(N__5307),
            .I(N__5280));
    ClkMux I__1184 (
            .O(N__5306),
            .I(N__5280));
    ClkMux I__1183 (
            .O(N__5305),
            .I(N__5280));
    ClkMux I__1182 (
            .O(N__5304),
            .I(N__5280));
    ClkMux I__1181 (
            .O(N__5303),
            .I(N__5280));
    ClkMux I__1180 (
            .O(N__5302),
            .I(N__5280));
    ClkMux I__1179 (
            .O(N__5301),
            .I(N__5280));
    ClkMux I__1178 (
            .O(N__5300),
            .I(N__5280));
    ClkMux I__1177 (
            .O(N__5299),
            .I(N__5280));
    GlobalMux I__1176 (
            .O(N__5280),
            .I(N__5277));
    gio2CtrlBuf I__1175 (
            .O(N__5277),
            .I(CLK6_c_g));
    InMux I__1174 (
            .O(N__5274),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ));
    InMux I__1173 (
            .O(N__5271),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ));
    InMux I__1172 (
            .O(N__5268),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ));
    InMux I__1171 (
            .O(N__5265),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ));
    CascadeMux I__1170 (
            .O(N__5262),
            .I(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_ ));
    InMux I__1169 (
            .O(N__5259),
            .I(N__5251));
    InMux I__1168 (
            .O(N__5258),
            .I(N__5251));
    InMux I__1167 (
            .O(N__5257),
            .I(N__5246));
    InMux I__1166 (
            .O(N__5256),
            .I(N__5246));
    LocalMux I__1165 (
            .O(N__5251),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__1164 (
            .O(N__5246),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    InMux I__1163 (
            .O(N__5241),
            .I(N__5227));
    InMux I__1162 (
            .O(N__5240),
            .I(N__5227));
    InMux I__1161 (
            .O(N__5239),
            .I(N__5227));
    InMux I__1160 (
            .O(N__5238),
            .I(N__5227));
    InMux I__1159 (
            .O(N__5237),
            .I(N__5222));
    InMux I__1158 (
            .O(N__5236),
            .I(N__5222));
    LocalMux I__1157 (
            .O(N__5227),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__1156 (
            .O(N__5222),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    CascadeMux I__1155 (
            .O(N__5217),
            .I(N__5213));
    InMux I__1154 (
            .O(N__5216),
            .I(N__5208));
    InMux I__1153 (
            .O(N__5213),
            .I(N__5203));
    InMux I__1152 (
            .O(N__5212),
            .I(N__5203));
    InMux I__1151 (
            .O(N__5211),
            .I(N__5200));
    LocalMux I__1150 (
            .O(N__5208),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__1149 (
            .O(N__5203),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__1148 (
            .O(N__5200),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    InMux I__1147 (
            .O(N__5193),
            .I(N__5190));
    LocalMux I__1146 (
            .O(N__5190),
            .I(N__5186));
    InMux I__1145 (
            .O(N__5189),
            .I(N__5183));
    Odrv4 I__1144 (
            .O(N__5186),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    LocalMux I__1143 (
            .O(N__5183),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    InMux I__1142 (
            .O(N__5178),
            .I(\U409_TICK.un2_COUNTER50_1_cry_7 ));
    InMux I__1141 (
            .O(N__5175),
            .I(N__5171));
    InMux I__1140 (
            .O(N__5174),
            .I(N__5168));
    LocalMux I__1139 (
            .O(N__5171),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    LocalMux I__1138 (
            .O(N__5168),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    CascadeMux I__1137 (
            .O(N__5163),
            .I(N__5160));
    InMux I__1136 (
            .O(N__5160),
            .I(N__5157));
    LocalMux I__1135 (
            .O(N__5157),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ));
    InMux I__1134 (
            .O(N__5154),
            .I(bfn_12_7_0_));
    InMux I__1133 (
            .O(N__5151),
            .I(N__5147));
    InMux I__1132 (
            .O(N__5150),
            .I(N__5144));
    LocalMux I__1131 (
            .O(N__5147),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    LocalMux I__1130 (
            .O(N__5144),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    InMux I__1129 (
            .O(N__5139),
            .I(\U409_TICK.un2_COUNTER50_1_cry_9 ));
    CascadeMux I__1128 (
            .O(N__5136),
            .I(N__5133));
    InMux I__1127 (
            .O(N__5133),
            .I(N__5129));
    InMux I__1126 (
            .O(N__5132),
            .I(N__5126));
    LocalMux I__1125 (
            .O(N__5129),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    LocalMux I__1124 (
            .O(N__5126),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    CascadeMux I__1123 (
            .O(N__5121),
            .I(N__5118));
    InMux I__1122 (
            .O(N__5118),
            .I(N__5115));
    LocalMux I__1121 (
            .O(N__5115),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ));
    InMux I__1120 (
            .O(N__5112),
            .I(\U409_TICK.un2_COUNTER50_1_cry_10 ));
    InMux I__1119 (
            .O(N__5109),
            .I(N__5105));
    InMux I__1118 (
            .O(N__5108),
            .I(N__5102));
    LocalMux I__1117 (
            .O(N__5105),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    LocalMux I__1116 (
            .O(N__5102),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    InMux I__1115 (
            .O(N__5097),
            .I(\U409_TICK.un2_COUNTER50_1_cry_11 ));
    InMux I__1114 (
            .O(N__5094),
            .I(N__5090));
    InMux I__1113 (
            .O(N__5093),
            .I(N__5087));
    LocalMux I__1112 (
            .O(N__5090),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    LocalMux I__1111 (
            .O(N__5087),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    InMux I__1110 (
            .O(N__5082),
            .I(N__5079));
    LocalMux I__1109 (
            .O(N__5079),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ));
    InMux I__1108 (
            .O(N__5076),
            .I(\U409_TICK.un2_COUNTER50_1_cry_12 ));
    InMux I__1107 (
            .O(N__5073),
            .I(N__5069));
    InMux I__1106 (
            .O(N__5072),
            .I(N__5066));
    LocalMux I__1105 (
            .O(N__5069),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    LocalMux I__1104 (
            .O(N__5066),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    InMux I__1103 (
            .O(N__5061),
            .I(N__5058));
    LocalMux I__1102 (
            .O(N__5058),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ));
    InMux I__1101 (
            .O(N__5055),
            .I(\U409_TICK.un2_COUNTER50_1_cry_13 ));
    InMux I__1100 (
            .O(N__5052),
            .I(N__5048));
    InMux I__1099 (
            .O(N__5051),
            .I(N__5045));
    LocalMux I__1098 (
            .O(N__5048),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    LocalMux I__1097 (
            .O(N__5045),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    CascadeMux I__1096 (
            .O(N__5040),
            .I(N__5037));
    InMux I__1095 (
            .O(N__5037),
            .I(N__5034));
    LocalMux I__1094 (
            .O(N__5034),
            .I(N__5031));
    Odrv4 I__1093 (
            .O(N__5031),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ));
    InMux I__1092 (
            .O(N__5028),
            .I(\U409_TICK.un2_COUNTER50_1_cry_14 ));
    InMux I__1091 (
            .O(N__5025),
            .I(N__5014));
    InMux I__1090 (
            .O(N__5024),
            .I(N__5014));
    InMux I__1089 (
            .O(N__5023),
            .I(N__5014));
    InMux I__1088 (
            .O(N__5022),
            .I(N__5009));
    InMux I__1087 (
            .O(N__5021),
            .I(N__5009));
    LocalMux I__1086 (
            .O(N__5014),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__1085 (
            .O(N__5009),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    CascadeMux I__1084 (
            .O(N__5004),
            .I(N__5001));
    InMux I__1083 (
            .O(N__5001),
            .I(N__4995));
    InMux I__1082 (
            .O(N__5000),
            .I(N__4990));
    InMux I__1081 (
            .O(N__4999),
            .I(N__4990));
    InMux I__1080 (
            .O(N__4998),
            .I(N__4987));
    LocalMux I__1079 (
            .O(N__4995),
            .I(N__4984));
    LocalMux I__1078 (
            .O(N__4990),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__1077 (
            .O(N__4987),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    Odrv4 I__1076 (
            .O(N__4984),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    IoInMux I__1075 (
            .O(N__4977),
            .I(N__4974));
    LocalMux I__1074 (
            .O(N__4974),
            .I(N__4971));
    Span4Mux_s2_v I__1073 (
            .O(N__4971),
            .I(N__4968));
    Span4Mux_v I__1072 (
            .O(N__4968),
            .I(N__4965));
    Odrv4 I__1071 (
            .O(N__4965),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__1070 (
            .O(N__4962),
            .I(N__4958));
    InMux I__1069 (
            .O(N__4961),
            .I(N__4952));
    InMux I__1068 (
            .O(N__4958),
            .I(N__4952));
    InMux I__1067 (
            .O(N__4957),
            .I(N__4949));
    LocalMux I__1066 (
            .O(N__4952),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    LocalMux I__1065 (
            .O(N__4949),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    CascadeMux I__1064 (
            .O(N__4944),
            .I(N__4938));
    InMux I__1063 (
            .O(N__4943),
            .I(N__4935));
    InMux I__1062 (
            .O(N__4942),
            .I(N__4930));
    InMux I__1061 (
            .O(N__4941),
            .I(N__4930));
    InMux I__1060 (
            .O(N__4938),
            .I(N__4927));
    LocalMux I__1059 (
            .O(N__4935),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__1058 (
            .O(N__4930),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__1057 (
            .O(N__4927),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    InMux I__1056 (
            .O(N__4920),
            .I(N__4916));
    InMux I__1055 (
            .O(N__4919),
            .I(N__4913));
    LocalMux I__1054 (
            .O(N__4916),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    LocalMux I__1053 (
            .O(N__4913),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    InMux I__1052 (
            .O(N__4908),
            .I(\U409_TICK.un2_COUNTER50_1_cry_1 ));
    InMux I__1051 (
            .O(N__4905),
            .I(N__4901));
    InMux I__1050 (
            .O(N__4904),
            .I(N__4898));
    LocalMux I__1049 (
            .O(N__4901),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    LocalMux I__1048 (
            .O(N__4898),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    InMux I__1047 (
            .O(N__4893),
            .I(\U409_TICK.un2_COUNTER50_1_cry_2 ));
    CascadeMux I__1046 (
            .O(N__4890),
            .I(N__4887));
    InMux I__1045 (
            .O(N__4887),
            .I(N__4884));
    LocalMux I__1044 (
            .O(N__4884),
            .I(N__4881));
    Span4Mux_h I__1043 (
            .O(N__4881),
            .I(N__4877));
    InMux I__1042 (
            .O(N__4880),
            .I(N__4874));
    Odrv4 I__1041 (
            .O(N__4877),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    LocalMux I__1040 (
            .O(N__4874),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    InMux I__1039 (
            .O(N__4869),
            .I(\U409_TICK.un2_COUNTER50_1_cry_3 ));
    InMux I__1038 (
            .O(N__4866),
            .I(N__4862));
    InMux I__1037 (
            .O(N__4865),
            .I(N__4859));
    LocalMux I__1036 (
            .O(N__4862),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    LocalMux I__1035 (
            .O(N__4859),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    InMux I__1034 (
            .O(N__4854),
            .I(N__4851));
    LocalMux I__1033 (
            .O(N__4851),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ));
    InMux I__1032 (
            .O(N__4848),
            .I(\U409_TICK.un2_COUNTER50_1_cry_4 ));
    InMux I__1031 (
            .O(N__4845),
            .I(N__4841));
    InMux I__1030 (
            .O(N__4844),
            .I(N__4838));
    LocalMux I__1029 (
            .O(N__4841),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    LocalMux I__1028 (
            .O(N__4838),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    InMux I__1027 (
            .O(N__4833),
            .I(N__4830));
    LocalMux I__1026 (
            .O(N__4830),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ));
    InMux I__1025 (
            .O(N__4827),
            .I(\U409_TICK.un2_COUNTER50_1_cry_5 ));
    InMux I__1024 (
            .O(N__4824),
            .I(N__4820));
    InMux I__1023 (
            .O(N__4823),
            .I(N__4817));
    LocalMux I__1022 (
            .O(N__4820),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    LocalMux I__1021 (
            .O(N__4817),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    InMux I__1020 (
            .O(N__4812),
            .I(\U409_TICK.un2_COUNTER50_1_cry_6 ));
    InMux I__1019 (
            .O(N__4809),
            .I(N__4803));
    InMux I__1018 (
            .O(N__4808),
            .I(N__4803));
    LocalMux I__1017 (
            .O(N__4803),
            .I(\U409_CIA.CLKCIA8_0_a2_0 ));
    CascadeMux I__1016 (
            .O(N__4800),
            .I(N__4791));
    InMux I__1015 (
            .O(N__4799),
            .I(N__4788));
    InMux I__1014 (
            .O(N__4798),
            .I(N__4785));
    InMux I__1013 (
            .O(N__4797),
            .I(N__4782));
    InMux I__1012 (
            .O(N__4796),
            .I(N__4773));
    InMux I__1011 (
            .O(N__4795),
            .I(N__4773));
    InMux I__1010 (
            .O(N__4794),
            .I(N__4773));
    InMux I__1009 (
            .O(N__4791),
            .I(N__4773));
    LocalMux I__1008 (
            .O(N__4788),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1007 (
            .O(N__4785),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1006 (
            .O(N__4782),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1005 (
            .O(N__4773),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    InMux I__1004 (
            .O(N__4764),
            .I(N__4757));
    InMux I__1003 (
            .O(N__4763),
            .I(N__4754));
    InMux I__1002 (
            .O(N__4762),
            .I(N__4747));
    InMux I__1001 (
            .O(N__4761),
            .I(N__4747));
    InMux I__1000 (
            .O(N__4760),
            .I(N__4747));
    LocalMux I__999 (
            .O(N__4757),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__998 (
            .O(N__4754),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__997 (
            .O(N__4747),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    InMux I__996 (
            .O(N__4740),
            .I(N__4735));
    InMux I__995 (
            .O(N__4739),
            .I(N__4730));
    InMux I__994 (
            .O(N__4738),
            .I(N__4730));
    LocalMux I__993 (
            .O(N__4735),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    LocalMux I__992 (
            .O(N__4730),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    CascadeMux I__991 (
            .O(N__4725),
            .I(N__4722));
    InMux I__990 (
            .O(N__4722),
            .I(N__4719));
    LocalMux I__989 (
            .O(N__4719),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ));
    CascadeMux I__988 (
            .O(N__4716),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_ ));
    InMux I__987 (
            .O(N__4713),
            .I(N__4705));
    InMux I__986 (
            .O(N__4712),
            .I(N__4705));
    InMux I__985 (
            .O(N__4711),
            .I(N__4702));
    InMux I__984 (
            .O(N__4710),
            .I(N__4699));
    LocalMux I__983 (
            .O(N__4705),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__982 (
            .O(N__4702),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__981 (
            .O(N__4699),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    IoInMux I__980 (
            .O(N__4692),
            .I(N__4689));
    LocalMux I__979 (
            .O(N__4689),
            .I(N__4684));
    CascadeMux I__978 (
            .O(N__4688),
            .I(N__4680));
    CascadeMux I__977 (
            .O(N__4687),
            .I(N__4676));
    Span4Mux_s2_v I__976 (
            .O(N__4684),
            .I(N__4673));
    CascadeMux I__975 (
            .O(N__4683),
            .I(N__4670));
    InMux I__974 (
            .O(N__4680),
            .I(N__4667));
    InMux I__973 (
            .O(N__4679),
            .I(N__4662));
    InMux I__972 (
            .O(N__4676),
            .I(N__4662));
    Span4Mux_v I__971 (
            .O(N__4673),
            .I(N__4659));
    InMux I__970 (
            .O(N__4670),
            .I(N__4656));
    LocalMux I__969 (
            .O(N__4667),
            .I(N__4653));
    LocalMux I__968 (
            .O(N__4662),
            .I(N__4649));
    Span4Mux_v I__967 (
            .O(N__4659),
            .I(N__4644));
    LocalMux I__966 (
            .O(N__4656),
            .I(N__4644));
    Span4Mux_v I__965 (
            .O(N__4653),
            .I(N__4641));
    InMux I__964 (
            .O(N__4652),
            .I(N__4638));
    Span4Mux_v I__963 (
            .O(N__4649),
            .I(N__4633));
    Span4Mux_v I__962 (
            .O(N__4644),
            .I(N__4633));
    Sp12to4 I__961 (
            .O(N__4641),
            .I(N__4630));
    LocalMux I__960 (
            .O(N__4638),
            .I(N__4627));
    Sp12to4 I__959 (
            .O(N__4633),
            .I(N__4624));
    Span12Mux_h I__958 (
            .O(N__4630),
            .I(N__4621));
    Sp12to4 I__957 (
            .O(N__4627),
            .I(N__4618));
    Span12Mux_h I__956 (
            .O(N__4624),
            .I(N__4615));
    Span12Mux_v I__955 (
            .O(N__4621),
            .I(N__4612));
    Span12Mux_v I__954 (
            .O(N__4618),
            .I(N__4609));
    Span12Mux_v I__953 (
            .O(N__4615),
            .I(N__4606));
    Odrv12 I__952 (
            .O(N__4612),
            .I(CLK40_IN_c));
    Odrv12 I__951 (
            .O(N__4609),
            .I(CLK40_IN_c));
    Odrv12 I__950 (
            .O(N__4606),
            .I(CLK40_IN_c));
    CascadeMux I__949 (
            .O(N__4599),
            .I(N__4594));
    InMux I__948 (
            .O(N__4598),
            .I(N__4591));
    InMux I__947 (
            .O(N__4597),
            .I(N__4588));
    InMux I__946 (
            .O(N__4594),
            .I(N__4585));
    LocalMux I__945 (
            .O(N__4591),
            .I(N__4580));
    LocalMux I__944 (
            .O(N__4588),
            .I(N__4580));
    LocalMux I__943 (
            .O(N__4585),
            .I(N__4577));
    Span4Mux_v I__942 (
            .O(N__4580),
            .I(N__4574));
    Span4Mux_v I__941 (
            .O(N__4577),
            .I(N__4571));
    Sp12to4 I__940 (
            .O(N__4574),
            .I(N__4568));
    Span4Mux_h I__939 (
            .O(N__4571),
            .I(N__4565));
    Span12Mux_h I__938 (
            .O(N__4568),
            .I(N__4560));
    Sp12to4 I__937 (
            .O(N__4565),
            .I(N__4560));
    Span12Mux_v I__936 (
            .O(N__4560),
            .I(N__4557));
    Odrv12 I__935 (
            .O(N__4557),
            .I(TSn_c));
    CascadeMux I__934 (
            .O(N__4554),
            .I(N__4550));
    InMux I__933 (
            .O(N__4553),
            .I(N__4547));
    InMux I__932 (
            .O(N__4550),
            .I(N__4544));
    LocalMux I__931 (
            .O(N__4547),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ));
    LocalMux I__930 (
            .O(N__4544),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ));
    InMux I__929 (
            .O(N__4539),
            .I(N__4532));
    InMux I__928 (
            .O(N__4538),
            .I(N__4532));
    InMux I__927 (
            .O(N__4537),
            .I(N__4529));
    LocalMux I__926 (
            .O(N__4532),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    LocalMux I__925 (
            .O(N__4529),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    CascadeMux I__924 (
            .O(N__4524),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ));
    InMux I__923 (
            .O(N__4521),
            .I(N__4518));
    LocalMux I__922 (
            .O(N__4518),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0 ));
    InMux I__921 (
            .O(N__4515),
            .I(N__4509));
    InMux I__920 (
            .O(N__4514),
            .I(N__4506));
    InMux I__919 (
            .O(N__4513),
            .I(N__4501));
    InMux I__918 (
            .O(N__4512),
            .I(N__4501));
    LocalMux I__917 (
            .O(N__4509),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__916 (
            .O(N__4506),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__915 (
            .O(N__4501),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    InMux I__914 (
            .O(N__4494),
            .I(N__4485));
    InMux I__913 (
            .O(N__4493),
            .I(N__4485));
    InMux I__912 (
            .O(N__4492),
            .I(N__4485));
    LocalMux I__911 (
            .O(N__4485),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ));
    CascadeMux I__910 (
            .O(N__4482),
            .I(N__4477));
    InMux I__909 (
            .O(N__4481),
            .I(N__4472));
    InMux I__908 (
            .O(N__4480),
            .I(N__4463));
    InMux I__907 (
            .O(N__4477),
            .I(N__4463));
    InMux I__906 (
            .O(N__4476),
            .I(N__4463));
    InMux I__905 (
            .O(N__4475),
            .I(N__4463));
    LocalMux I__904 (
            .O(N__4472),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__903 (
            .O(N__4463),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    CascadeMux I__902 (
            .O(N__4458),
            .I(N__4455));
    InMux I__901 (
            .O(N__4455),
            .I(N__4443));
    InMux I__900 (
            .O(N__4454),
            .I(N__4443));
    InMux I__899 (
            .O(N__4453),
            .I(N__4436));
    InMux I__898 (
            .O(N__4452),
            .I(N__4436));
    InMux I__897 (
            .O(N__4451),
            .I(N__4436));
    InMux I__896 (
            .O(N__4450),
            .I(N__4429));
    InMux I__895 (
            .O(N__4449),
            .I(N__4429));
    InMux I__894 (
            .O(N__4448),
            .I(N__4429));
    LocalMux I__893 (
            .O(N__4443),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__892 (
            .O(N__4436),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__891 (
            .O(N__4429),
            .I(\U409_TICK.TICK503_14 ));
    InMux I__890 (
            .O(N__4422),
            .I(N__4410));
    InMux I__889 (
            .O(N__4421),
            .I(N__4410));
    InMux I__888 (
            .O(N__4420),
            .I(N__4403));
    InMux I__887 (
            .O(N__4419),
            .I(N__4403));
    InMux I__886 (
            .O(N__4418),
            .I(N__4403));
    InMux I__885 (
            .O(N__4417),
            .I(N__4396));
    InMux I__884 (
            .O(N__4416),
            .I(N__4396));
    InMux I__883 (
            .O(N__4415),
            .I(N__4396));
    LocalMux I__882 (
            .O(N__4410),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__881 (
            .O(N__4403),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__880 (
            .O(N__4396),
            .I(\U409_TICK.TICK503_10 ));
    CascadeMux I__879 (
            .O(N__4389),
            .I(N__4384));
    CascadeMux I__878 (
            .O(N__4388),
            .I(N__4379));
    InMux I__877 (
            .O(N__4387),
            .I(N__4371));
    InMux I__876 (
            .O(N__4384),
            .I(N__4371));
    InMux I__875 (
            .O(N__4383),
            .I(N__4364));
    InMux I__874 (
            .O(N__4382),
            .I(N__4364));
    InMux I__873 (
            .O(N__4379),
            .I(N__4364));
    InMux I__872 (
            .O(N__4378),
            .I(N__4357));
    InMux I__871 (
            .O(N__4377),
            .I(N__4357));
    InMux I__870 (
            .O(N__4376),
            .I(N__4357));
    LocalMux I__869 (
            .O(N__4371),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__868 (
            .O(N__4364),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__867 (
            .O(N__4357),
            .I(\U409_TICK.TICK503_9 ));
    IoInMux I__866 (
            .O(N__4350),
            .I(N__4347));
    LocalMux I__865 (
            .O(N__4347),
            .I(N__4344));
    Span4Mux_s1_v I__864 (
            .O(N__4344),
            .I(N__4341));
    Sp12to4 I__863 (
            .O(N__4341),
            .I(N__4338));
    Span12Mux_h I__862 (
            .O(N__4338),
            .I(N__4335));
    Span12Mux_v I__861 (
            .O(N__4335),
            .I(N__4331));
    InMux I__860 (
            .O(N__4334),
            .I(N__4328));
    Odrv12 I__859 (
            .O(N__4331),
            .I(TICK50_c));
    LocalMux I__858 (
            .O(N__4328),
            .I(TICK50_c));
    CascadeMux I__857 (
            .O(N__4323),
            .I(\U409_CIA.N_9_cascade_ ));
    CascadeMux I__856 (
            .O(N__4320),
            .I(N__4317));
    InMux I__855 (
            .O(N__4317),
            .I(N__4313));
    CascadeMux I__854 (
            .O(N__4316),
            .I(N__4309));
    LocalMux I__853 (
            .O(N__4313),
            .I(N__4305));
    InMux I__852 (
            .O(N__4312),
            .I(N__4300));
    InMux I__851 (
            .O(N__4309),
            .I(N__4300));
    InMux I__850 (
            .O(N__4308),
            .I(N__4297));
    Span4Mux_v I__849 (
            .O(N__4305),
            .I(N__4292));
    LocalMux I__848 (
            .O(N__4300),
            .I(N__4292));
    LocalMux I__847 (
            .O(N__4297),
            .I(\U409_CIA.VMAZ0 ));
    Odrv4 I__846 (
            .O(N__4292),
            .I(\U409_CIA.VMAZ0 ));
    CascadeMux I__845 (
            .O(N__4287),
            .I(\U409_CIA.N_20_cascade_ ));
    InMux I__844 (
            .O(N__4284),
            .I(N__4281));
    LocalMux I__843 (
            .O(N__4281),
            .I(\U409_CIA.CLKCIA6_0_a2_1 ));
    CascadeMux I__842 (
            .O(N__4278),
            .I(\U409_CIA.CLKCIAZ0_cascade_ ));
    IoInMux I__841 (
            .O(N__4275),
            .I(N__4272));
    LocalMux I__840 (
            .O(N__4272),
            .I(N__4269));
    Span4Mux_s1_v I__839 (
            .O(N__4269),
            .I(N__4266));
    Span4Mux_v I__838 (
            .O(N__4266),
            .I(N__4263));
    Sp12to4 I__837 (
            .O(N__4263),
            .I(N__4260));
    Span12Mux_h I__836 (
            .O(N__4260),
            .I(N__4257));
    Span12Mux_v I__835 (
            .O(N__4257),
            .I(N__4252));
    InMux I__834 (
            .O(N__4256),
            .I(N__4249));
    InMux I__833 (
            .O(N__4255),
            .I(N__4246));
    Odrv12 I__832 (
            .O(N__4252),
            .I(CLKCIA_c));
    LocalMux I__831 (
            .O(N__4249),
            .I(CLKCIA_c));
    LocalMux I__830 (
            .O(N__4246),
            .I(CLKCIA_c));
    InMux I__829 (
            .O(N__4239),
            .I(N__4235));
    InMux I__828 (
            .O(N__4238),
            .I(N__4232));
    LocalMux I__827 (
            .O(N__4235),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    LocalMux I__826 (
            .O(N__4232),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    InMux I__825 (
            .O(N__4227),
            .I(N__4224));
    LocalMux I__824 (
            .O(N__4224),
            .I(\U409_TICK.TICK503_11 ));
    CascadeMux I__823 (
            .O(N__4221),
            .I(\U409_TICK.TICK503_8_cascade_ ));
    CascadeMux I__822 (
            .O(N__4218),
            .I(\U409_TICK.TICK503_14_cascade_ ));
    CascadeMux I__821 (
            .O(N__4215),
            .I(\U409_TICK.TICK503_10_cascade_ ));
    CascadeMux I__820 (
            .O(N__4212),
            .I(\U409_TICK.TICK503_9_cascade_ ));
    IoInMux I__819 (
            .O(N__4209),
            .I(N__4206));
    LocalMux I__818 (
            .O(N__4206),
            .I(N__4203));
    Span4Mux_s2_v I__817 (
            .O(N__4203),
            .I(N__4200));
    Span4Mux_v I__816 (
            .O(N__4200),
            .I(N__4197));
    Span4Mux_v I__815 (
            .O(N__4197),
            .I(N__4194));
    Span4Mux_h I__814 (
            .O(N__4194),
            .I(N__4190));
    InMux I__813 (
            .O(N__4193),
            .I(N__4187));
    Odrv4 I__812 (
            .O(N__4190),
            .I(TICK60_c));
    LocalMux I__811 (
            .O(N__4187),
            .I(TICK60_c));
    InMux I__810 (
            .O(N__4182),
            .I(N__4179));
    LocalMux I__809 (
            .O(N__4179),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ));
    CascadeMux I__808 (
            .O(N__4176),
            .I(N__4173));
    InMux I__807 (
            .O(N__4173),
            .I(N__4170));
    LocalMux I__806 (
            .O(N__4170),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ));
    InMux I__805 (
            .O(N__4167),
            .I(N__4163));
    InMux I__804 (
            .O(N__4166),
            .I(N__4160));
    LocalMux I__803 (
            .O(N__4163),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    LocalMux I__802 (
            .O(N__4160),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    InMux I__801 (
            .O(N__4155),
            .I(N__4151));
    InMux I__800 (
            .O(N__4154),
            .I(N__4148));
    LocalMux I__799 (
            .O(N__4151),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    LocalMux I__798 (
            .O(N__4148),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    InMux I__797 (
            .O(N__4143),
            .I(N__4139));
    InMux I__796 (
            .O(N__4142),
            .I(N__4136));
    LocalMux I__795 (
            .O(N__4139),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    LocalMux I__794 (
            .O(N__4136),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    CascadeMux I__793 (
            .O(N__4131),
            .I(N__4128));
    InMux I__792 (
            .O(N__4128),
            .I(N__4125));
    LocalMux I__791 (
            .O(N__4125),
            .I(N__4121));
    InMux I__790 (
            .O(N__4124),
            .I(N__4118));
    Odrv4 I__789 (
            .O(N__4121),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    LocalMux I__788 (
            .O(N__4118),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    InMux I__787 (
            .O(N__4113),
            .I(N__4109));
    InMux I__786 (
            .O(N__4112),
            .I(N__4106));
    LocalMux I__785 (
            .O(N__4109),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    LocalMux I__784 (
            .O(N__4106),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    CascadeMux I__783 (
            .O(N__4101),
            .I(N__4096));
    CascadeMux I__782 (
            .O(N__4100),
            .I(N__4092));
    InMux I__781 (
            .O(N__4099),
            .I(N__4084));
    InMux I__780 (
            .O(N__4096),
            .I(N__4084));
    InMux I__779 (
            .O(N__4095),
            .I(N__4079));
    InMux I__778 (
            .O(N__4092),
            .I(N__4079));
    InMux I__777 (
            .O(N__4091),
            .I(N__4072));
    InMux I__776 (
            .O(N__4090),
            .I(N__4072));
    InMux I__775 (
            .O(N__4089),
            .I(N__4072));
    LocalMux I__774 (
            .O(N__4084),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__773 (
            .O(N__4079),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__772 (
            .O(N__4072),
            .I(\U409_TICK.TICK603_10 ));
    CascadeMux I__771 (
            .O(N__4065),
            .I(N__4059));
    InMux I__770 (
            .O(N__4064),
            .I(N__4050));
    InMux I__769 (
            .O(N__4063),
            .I(N__4050));
    InMux I__768 (
            .O(N__4062),
            .I(N__4043));
    InMux I__767 (
            .O(N__4059),
            .I(N__4043));
    InMux I__766 (
            .O(N__4058),
            .I(N__4043));
    InMux I__765 (
            .O(N__4057),
            .I(N__4036));
    InMux I__764 (
            .O(N__4056),
            .I(N__4036));
    InMux I__763 (
            .O(N__4055),
            .I(N__4036));
    LocalMux I__762 (
            .O(N__4050),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__761 (
            .O(N__4043),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__760 (
            .O(N__4036),
            .I(\U409_TICK.TICK603_9 ));
    InMux I__759 (
            .O(N__4029),
            .I(N__4019));
    InMux I__758 (
            .O(N__4028),
            .I(N__4019));
    InMux I__757 (
            .O(N__4027),
            .I(N__4019));
    CascadeMux I__756 (
            .O(N__4026),
            .I(N__4016));
    LocalMux I__755 (
            .O(N__4019),
            .I(N__4010));
    InMux I__754 (
            .O(N__4016),
            .I(N__4007));
    InMux I__753 (
            .O(N__4015),
            .I(N__4004));
    InMux I__752 (
            .O(N__4014),
            .I(N__4001));
    InMux I__751 (
            .O(N__4013),
            .I(N__3998));
    Span4Mux_v I__750 (
            .O(N__4010),
            .I(N__3995));
    LocalMux I__749 (
            .O(N__4007),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__748 (
            .O(N__4004),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__747 (
            .O(N__4001),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__746 (
            .O(N__3998),
            .I(\U409_TICK.TICK603_14 ));
    Odrv4 I__745 (
            .O(N__3995),
            .I(\U409_TICK.TICK603_14 ));
    CascadeMux I__744 (
            .O(N__3984),
            .I(\U409_TICK.TICK603_10_cascade_ ));
    InMux I__743 (
            .O(N__3981),
            .I(N__3978));
    LocalMux I__742 (
            .O(N__3978),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ));
    CascadeMux I__741 (
            .O(N__3975),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_ ));
    CascadeMux I__740 (
            .O(N__3972),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_ ));
    CascadeMux I__739 (
            .O(N__3969),
            .I(N__3964));
    CascadeMux I__738 (
            .O(N__3968),
            .I(N__3961));
    InMux I__737 (
            .O(N__3967),
            .I(N__3957));
    InMux I__736 (
            .O(N__3964),
            .I(N__3950));
    InMux I__735 (
            .O(N__3961),
            .I(N__3950));
    InMux I__734 (
            .O(N__3960),
            .I(N__3950));
    LocalMux I__733 (
            .O(N__3957),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__732 (
            .O(N__3950),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    InMux I__731 (
            .O(N__3945),
            .I(N__3939));
    InMux I__730 (
            .O(N__3944),
            .I(N__3939));
    LocalMux I__729 (
            .O(N__3939),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ));
    InMux I__728 (
            .O(N__3936),
            .I(N__3931));
    InMux I__727 (
            .O(N__3935),
            .I(N__3928));
    InMux I__726 (
            .O(N__3934),
            .I(N__3925));
    LocalMux I__725 (
            .O(N__3931),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__724 (
            .O(N__3928),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__723 (
            .O(N__3925),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    CascadeMux I__722 (
            .O(N__3918),
            .I(N__3914));
    CascadeMux I__721 (
            .O(N__3917),
            .I(N__3909));
    InMux I__720 (
            .O(N__3914),
            .I(N__3904));
    InMux I__719 (
            .O(N__3913),
            .I(N__3904));
    InMux I__718 (
            .O(N__3912),
            .I(N__3901));
    InMux I__717 (
            .O(N__3909),
            .I(N__3898));
    LocalMux I__716 (
            .O(N__3904),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__715 (
            .O(N__3901),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__714 (
            .O(N__3898),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    InMux I__713 (
            .O(N__3891),
            .I(N__3888));
    LocalMux I__712 (
            .O(N__3888),
            .I(N__3884));
    InMux I__711 (
            .O(N__3887),
            .I(N__3881));
    Odrv4 I__710 (
            .O(N__3884),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    LocalMux I__709 (
            .O(N__3881),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    InMux I__708 (
            .O(N__3876),
            .I(\U409_TICK.un3_COUNTER60_1_cry_10 ));
    InMux I__707 (
            .O(N__3873),
            .I(N__3870));
    LocalMux I__706 (
            .O(N__3870),
            .I(N__3866));
    InMux I__705 (
            .O(N__3869),
            .I(N__3863));
    Span4Mux_v I__704 (
            .O(N__3866),
            .I(N__3860));
    LocalMux I__703 (
            .O(N__3863),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    Odrv4 I__702 (
            .O(N__3860),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    InMux I__701 (
            .O(N__3855),
            .I(\U409_TICK.un3_COUNTER60_1_cry_11 ));
    InMux I__700 (
            .O(N__3852),
            .I(\U409_TICK.un3_COUNTER60_1_cry_12 ));
    InMux I__699 (
            .O(N__3849),
            .I(\U409_TICK.un3_COUNTER60_1_cry_13 ));
    InMux I__698 (
            .O(N__3846),
            .I(\U409_TICK.un3_COUNTER60_1_cry_14 ));
    InMux I__697 (
            .O(N__3843),
            .I(\U409_TICK.un3_COUNTER60_1_cry_15 ));
    CascadeMux I__696 (
            .O(N__3840),
            .I(N__3837));
    InMux I__695 (
            .O(N__3837),
            .I(N__3833));
    InMux I__694 (
            .O(N__3836),
            .I(N__3830));
    LocalMux I__693 (
            .O(N__3833),
            .I(N__3827));
    LocalMux I__692 (
            .O(N__3830),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    Odrv4 I__691 (
            .O(N__3827),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    InMux I__690 (
            .O(N__3822),
            .I(N__3813));
    InMux I__689 (
            .O(N__3821),
            .I(N__3813));
    InMux I__688 (
            .O(N__3820),
            .I(N__3813));
    LocalMux I__687 (
            .O(N__3813),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    InMux I__686 (
            .O(N__3810),
            .I(N__3806));
    InMux I__685 (
            .O(N__3809),
            .I(N__3803));
    LocalMux I__684 (
            .O(N__3806),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    LocalMux I__683 (
            .O(N__3803),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    InMux I__682 (
            .O(N__3798),
            .I(N__3794));
    InMux I__681 (
            .O(N__3797),
            .I(N__3791));
    LocalMux I__680 (
            .O(N__3794),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    LocalMux I__679 (
            .O(N__3791),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    InMux I__678 (
            .O(N__3786),
            .I(\U409_TICK.un3_COUNTER60_1_cry_2 ));
    InMux I__677 (
            .O(N__3783),
            .I(N__3779));
    InMux I__676 (
            .O(N__3782),
            .I(N__3776));
    LocalMux I__675 (
            .O(N__3779),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    LocalMux I__674 (
            .O(N__3776),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    InMux I__673 (
            .O(N__3771),
            .I(N__3768));
    LocalMux I__672 (
            .O(N__3768),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ));
    InMux I__671 (
            .O(N__3765),
            .I(\U409_TICK.un3_COUNTER60_1_cry_3 ));
    InMux I__670 (
            .O(N__3762),
            .I(N__3758));
    InMux I__669 (
            .O(N__3761),
            .I(N__3755));
    LocalMux I__668 (
            .O(N__3758),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    LocalMux I__667 (
            .O(N__3755),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    InMux I__666 (
            .O(N__3750),
            .I(\U409_TICK.un3_COUNTER60_1_cry_4 ));
    InMux I__665 (
            .O(N__3747),
            .I(N__3743));
    InMux I__664 (
            .O(N__3746),
            .I(N__3740));
    LocalMux I__663 (
            .O(N__3743),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    LocalMux I__662 (
            .O(N__3740),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    InMux I__661 (
            .O(N__3735),
            .I(N__3732));
    LocalMux I__660 (
            .O(N__3732),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ));
    InMux I__659 (
            .O(N__3729),
            .I(\U409_TICK.un3_COUNTER60_1_cry_5 ));
    InMux I__658 (
            .O(N__3726),
            .I(\U409_TICK.un3_COUNTER60_1_cry_6 ));
    CascadeMux I__657 (
            .O(N__3723),
            .I(N__3720));
    InMux I__656 (
            .O(N__3720),
            .I(N__3716));
    InMux I__655 (
            .O(N__3719),
            .I(N__3713));
    LocalMux I__654 (
            .O(N__3716),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    LocalMux I__653 (
            .O(N__3713),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    InMux I__652 (
            .O(N__3708),
            .I(N__3705));
    LocalMux I__651 (
            .O(N__3705),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ));
    InMux I__650 (
            .O(N__3702),
            .I(\U409_TICK.un3_COUNTER60_1_cry_7 ));
    InMux I__649 (
            .O(N__3699),
            .I(bfn_10_7_0_));
    InMux I__648 (
            .O(N__3696),
            .I(\U409_TICK.un3_COUNTER60_1_cry_9 ));
    CascadeMux I__647 (
            .O(N__3693),
            .I(\U409_TICK.TICK603_11_cascade_ ));
    CascadeMux I__646 (
            .O(N__3690),
            .I(\U409_TICK.TICK603_14_cascade_ ));
    InMux I__645 (
            .O(N__3687),
            .I(N__3684));
    LocalMux I__644 (
            .O(N__3684),
            .I(\U409_TICK.TICK603_8 ));
    InMux I__643 (
            .O(N__3681),
            .I(N__3677));
    InMux I__642 (
            .O(N__3680),
            .I(N__3674));
    LocalMux I__641 (
            .O(N__3677),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    LocalMux I__640 (
            .O(N__3674),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    InMux I__639 (
            .O(N__3669),
            .I(\U409_TICK.un3_COUNTER60_1_cry_1 ));
    InMux I__638 (
            .O(N__3666),
            .I(N__3659));
    InMux I__637 (
            .O(N__3665),
            .I(N__3656));
    InMux I__636 (
            .O(N__3664),
            .I(N__3649));
    InMux I__635 (
            .O(N__3663),
            .I(N__3649));
    InMux I__634 (
            .O(N__3662),
            .I(N__3649));
    LocalMux I__633 (
            .O(N__3659),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__632 (
            .O(N__3656),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__631 (
            .O(N__3649),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    InMux I__630 (
            .O(N__3642),
            .I(N__3638));
    InMux I__629 (
            .O(N__3641),
            .I(N__3635));
    LocalMux I__628 (
            .O(N__3638),
            .I(\U409_TRANSFER_ACK.N_97 ));
    LocalMux I__627 (
            .O(N__3635),
            .I(\U409_TRANSFER_ACK.N_97 ));
    CascadeMux I__626 (
            .O(N__3630),
            .I(N__3626));
    CascadeMux I__625 (
            .O(N__3629),
            .I(N__3623));
    InMux I__624 (
            .O(N__3626),
            .I(N__3620));
    InMux I__623 (
            .O(N__3623),
            .I(N__3615));
    LocalMux I__622 (
            .O(N__3620),
            .I(N__3612));
    InMux I__621 (
            .O(N__3619),
            .I(N__3607));
    InMux I__620 (
            .O(N__3618),
            .I(N__3607));
    LocalMux I__619 (
            .O(N__3615),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    Odrv12 I__618 (
            .O(N__3612),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__617 (
            .O(N__3607),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    CascadeMux I__616 (
            .O(N__3600),
            .I(\U409_TRANSFER_ACK.CIA_TACK_EN_0_cascade_ ));
    IoInMux I__615 (
            .O(N__3597),
            .I(N__3594));
    LocalMux I__614 (
            .O(N__3594),
            .I(N__3591));
    Span4Mux_s2_v I__613 (
            .O(N__3591),
            .I(N__3588));
    Span4Mux_h I__612 (
            .O(N__3588),
            .I(N__3585));
    Span4Mux_v I__611 (
            .O(N__3585),
            .I(N__3582));
    Sp12to4 I__610 (
            .O(N__3582),
            .I(N__3579));
    Span12Mux_h I__609 (
            .O(N__3579),
            .I(N__3575));
    InMux I__608 (
            .O(N__3578),
            .I(N__3572));
    Odrv12 I__607 (
            .O(N__3575),
            .I(TACK_OUTn));
    LocalMux I__606 (
            .O(N__3572),
            .I(TACK_OUTn));
    InMux I__605 (
            .O(N__3567),
            .I(N__3563));
    InMux I__604 (
            .O(N__3566),
            .I(N__3560));
    LocalMux I__603 (
            .O(N__3563),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    LocalMux I__602 (
            .O(N__3560),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    InMux I__601 (
            .O(N__3555),
            .I(N__3546));
    InMux I__600 (
            .O(N__3554),
            .I(N__3546));
    InMux I__599 (
            .O(N__3553),
            .I(N__3546));
    LocalMux I__598 (
            .O(N__3546),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    CascadeMux I__597 (
            .O(N__3543),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_ ));
    InMux I__596 (
            .O(N__3540),
            .I(N__3536));
    InMux I__595 (
            .O(N__3539),
            .I(N__3533));
    LocalMux I__594 (
            .O(N__3536),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    LocalMux I__593 (
            .O(N__3533),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    CascadeMux I__592 (
            .O(N__3528),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_ ));
    InMux I__591 (
            .O(N__3525),
            .I(N__3516));
    InMux I__590 (
            .O(N__3524),
            .I(N__3516));
    InMux I__589 (
            .O(N__3523),
            .I(N__3516));
    LocalMux I__588 (
            .O(N__3516),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    InMux I__587 (
            .O(N__3513),
            .I(N__3509));
    InMux I__586 (
            .O(N__3512),
            .I(N__3506));
    LocalMux I__585 (
            .O(N__3509),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ));
    LocalMux I__584 (
            .O(N__3506),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ));
    CEMux I__583 (
            .O(N__3501),
            .I(N__3498));
    LocalMux I__582 (
            .O(N__3498),
            .I(N__3495));
    Span4Mux_v I__581 (
            .O(N__3495),
            .I(N__3492));
    Span4Mux_h I__580 (
            .O(N__3492),
            .I(N__3489));
    Odrv4 I__579 (
            .O(N__3489),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0 ));
    CascadeMux I__578 (
            .O(N__3486),
            .I(\U409_TRANSFER_ACK.m9_bm_cascade_ ));
    CascadeMux I__577 (
            .O(N__3483),
            .I(\U409_TRANSFER_ACK.N_4_cascade_ ));
    InMux I__576 (
            .O(N__3480),
            .I(N__3477));
    LocalMux I__575 (
            .O(N__3477),
            .I(\U409_TRANSFER_ACK.m9_am ));
    InMux I__574 (
            .O(N__3474),
            .I(N__3468));
    InMux I__573 (
            .O(N__3473),
            .I(N__3468));
    LocalMux I__572 (
            .O(N__3468),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    InMux I__571 (
            .O(N__3465),
            .I(N__3462));
    LocalMux I__570 (
            .O(N__3462),
            .I(\U409_TRANSFER_ACK.N_4 ));
    CascadeMux I__569 (
            .O(N__3459),
            .I(\U409_TRANSFER_ACK.i6_mux_0_cascade_ ));
    InMux I__568 (
            .O(N__3456),
            .I(N__3450));
    InMux I__567 (
            .O(N__3455),
            .I(N__3447));
    InMux I__566 (
            .O(N__3454),
            .I(N__3442));
    InMux I__565 (
            .O(N__3453),
            .I(N__3442));
    LocalMux I__564 (
            .O(N__3450),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__563 (
            .O(N__3447),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__562 (
            .O(N__3442),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    CascadeMux I__561 (
            .O(N__3435),
            .I(N__3432));
    InMux I__560 (
            .O(N__3432),
            .I(N__3427));
    InMux I__559 (
            .O(N__3431),
            .I(N__3424));
    InMux I__558 (
            .O(N__3430),
            .I(N__3421));
    LocalMux I__557 (
            .O(N__3427),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    LocalMux I__556 (
            .O(N__3424),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    LocalMux I__555 (
            .O(N__3421),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    SRMux I__554 (
            .O(N__3414),
            .I(N__3411));
    LocalMux I__553 (
            .O(N__3411),
            .I(N__3408));
    Odrv4 I__552 (
            .O(N__3408),
            .I(\U409_TRANSFER_ACK.RESETn_c_i ));
    InMux I__551 (
            .O(N__3405),
            .I(N__3401));
    InMux I__550 (
            .O(N__3404),
            .I(N__3398));
    LocalMux I__549 (
            .O(N__3401),
            .I(N__3393));
    LocalMux I__548 (
            .O(N__3398),
            .I(N__3393));
    Odrv12 I__547 (
            .O(N__3393),
            .I(CIA_ENABLEm));
    InMux I__546 (
            .O(N__3390),
            .I(N__3387));
    LocalMux I__545 (
            .O(N__3387),
            .I(N__3383));
    CascadeMux I__544 (
            .O(N__3386),
            .I(N__3380));
    Span4Mux_v I__543 (
            .O(N__3383),
            .I(N__3376));
    InMux I__542 (
            .O(N__3380),
            .I(N__3373));
    InMux I__541 (
            .O(N__3379),
            .I(N__3370));
    Sp12to4 I__540 (
            .O(N__3376),
            .I(N__3363));
    LocalMux I__539 (
            .O(N__3373),
            .I(N__3363));
    LocalMux I__538 (
            .O(N__3370),
            .I(N__3363));
    Span12Mux_h I__537 (
            .O(N__3363),
            .I(N__3360));
    Odrv12 I__536 (
            .O(N__3360),
            .I(\U409_CIA.g0Z0Z_14 ));
    InMux I__535 (
            .O(N__3357),
            .I(N__3353));
    InMux I__534 (
            .O(N__3356),
            .I(N__3350));
    LocalMux I__533 (
            .O(N__3353),
            .I(N__3346));
    LocalMux I__532 (
            .O(N__3350),
            .I(N__3343));
    InMux I__531 (
            .O(N__3349),
            .I(N__3340));
    Span4Mux_v I__530 (
            .O(N__3346),
            .I(N__3337));
    Span4Mux_h I__529 (
            .O(N__3343),
            .I(N__3332));
    LocalMux I__528 (
            .O(N__3340),
            .I(N__3332));
    Span4Mux_v I__527 (
            .O(N__3337),
            .I(N__3327));
    Span4Mux_v I__526 (
            .O(N__3332),
            .I(N__3327));
    Sp12to4 I__525 (
            .O(N__3327),
            .I(N__3324));
    Span12Mux_h I__524 (
            .O(N__3324),
            .I(N__3321));
    Odrv12 I__523 (
            .O(N__3321),
            .I(\U409_CIA.g0Z0Z_13 ));
    InMux I__522 (
            .O(N__3318),
            .I(N__3313));
    InMux I__521 (
            .O(N__3317),
            .I(N__3308));
    InMux I__520 (
            .O(N__3316),
            .I(N__3308));
    LocalMux I__519 (
            .O(N__3313),
            .I(\U409_CIA.CIA_HOLDZ0 ));
    LocalMux I__518 (
            .O(N__3308),
            .I(\U409_CIA.CIA_HOLDZ0 ));
    CascadeMux I__517 (
            .O(N__3303),
            .I(\U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0_cascade_ ));
    CascadeMux I__516 (
            .O(N__3300),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_3_0_cascade_ ));
    InMux I__515 (
            .O(N__3297),
            .I(N__3294));
    LocalMux I__514 (
            .O(N__3294),
            .I(\U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0 ));
    CascadeMux I__513 (
            .O(N__3291),
            .I(N__3287));
    InMux I__512 (
            .O(N__3290),
            .I(N__3281));
    InMux I__511 (
            .O(N__3287),
            .I(N__3272));
    InMux I__510 (
            .O(N__3286),
            .I(N__3272));
    InMux I__509 (
            .O(N__3285),
            .I(N__3272));
    InMux I__508 (
            .O(N__3284),
            .I(N__3272));
    LocalMux I__507 (
            .O(N__3281),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__506 (
            .O(N__3272),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    InMux I__505 (
            .O(N__3267),
            .I(N__3255));
    InMux I__504 (
            .O(N__3266),
            .I(N__3255));
    InMux I__503 (
            .O(N__3265),
            .I(N__3255));
    InMux I__502 (
            .O(N__3264),
            .I(N__3255));
    LocalMux I__501 (
            .O(N__3255),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    InMux I__500 (
            .O(N__3252),
            .I(N__3249));
    LocalMux I__499 (
            .O(N__3249),
            .I(\U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa ));
    InMux I__498 (
            .O(N__3246),
            .I(N__3241));
    InMux I__497 (
            .O(N__3245),
            .I(N__3238));
    InMux I__496 (
            .O(N__3244),
            .I(N__3235));
    LocalMux I__495 (
            .O(N__3241),
            .I(N__3228));
    LocalMux I__494 (
            .O(N__3238),
            .I(N__3228));
    LocalMux I__493 (
            .O(N__3235),
            .I(N__3228));
    Span4Mux_v I__492 (
            .O(N__3228),
            .I(N__3222));
    InMux I__491 (
            .O(N__3227),
            .I(N__3219));
    InMux I__490 (
            .O(N__3226),
            .I(N__3214));
    InMux I__489 (
            .O(N__3225),
            .I(N__3214));
    Sp12to4 I__488 (
            .O(N__3222),
            .I(N__3206));
    LocalMux I__487 (
            .O(N__3219),
            .I(N__3206));
    LocalMux I__486 (
            .O(N__3214),
            .I(N__3206));
    InMux I__485 (
            .O(N__3213),
            .I(N__3203));
    Span12Mux_h I__484 (
            .O(N__3206),
            .I(N__3200));
    LocalMux I__483 (
            .O(N__3203),
            .I(N__3197));
    Odrv12 I__482 (
            .O(N__3200),
            .I(U409_ADDRESS_DECODE_Z2_SPACE));
    Odrv12 I__481 (
            .O(N__3197),
            .I(U409_ADDRESS_DECODE_Z2_SPACE));
    InMux I__480 (
            .O(N__3192),
            .I(N__3188));
    InMux I__479 (
            .O(N__3191),
            .I(N__3185));
    LocalMux I__478 (
            .O(N__3188),
            .I(U409_ADDRESS_DECODE_un1_ROMEN_0));
    LocalMux I__477 (
            .O(N__3185),
            .I(U409_ADDRESS_DECODE_un1_ROMEN_0));
    IoInMux I__476 (
            .O(N__3180),
            .I(N__3177));
    LocalMux I__475 (
            .O(N__3177),
            .I(N__3174));
    Span4Mux_s3_v I__474 (
            .O(N__3174),
            .I(N__3171));
    Sp12to4 I__473 (
            .O(N__3171),
            .I(N__3168));
    Span12Mux_h I__472 (
            .O(N__3168),
            .I(N__3165));
    Odrv12 I__471 (
            .O(N__3165),
            .I(ROMENm_i));
    IoInMux I__470 (
            .O(N__3162),
            .I(N__3159));
    LocalMux I__469 (
            .O(N__3159),
            .I(N__3156));
    Span4Mux_s1_v I__468 (
            .O(N__3156),
            .I(N__3153));
    Sp12to4 I__467 (
            .O(N__3153),
            .I(N__3150));
    Span12Mux_h I__466 (
            .O(N__3150),
            .I(N__3147));
    Span12Mux_v I__465 (
            .O(N__3147),
            .I(N__3144));
    Odrv12 I__464 (
            .O(N__3144),
            .I(PORTSIZE_0_i));
    InMux I__463 (
            .O(N__3141),
            .I(N__3131));
    InMux I__462 (
            .O(N__3140),
            .I(N__3131));
    InMux I__461 (
            .O(N__3139),
            .I(N__3131));
    InMux I__460 (
            .O(N__3138),
            .I(N__3126));
    LocalMux I__459 (
            .O(N__3131),
            .I(N__3123));
    InMux I__458 (
            .O(N__3130),
            .I(N__3120));
    InMux I__457 (
            .O(N__3129),
            .I(N__3117));
    LocalMux I__456 (
            .O(N__3126),
            .I(N__3114));
    Span4Mux_v I__455 (
            .O(N__3123),
            .I(N__3111));
    LocalMux I__454 (
            .O(N__3120),
            .I(N__3106));
    LocalMux I__453 (
            .O(N__3117),
            .I(N__3106));
    Span4Mux_v I__452 (
            .O(N__3114),
            .I(N__3103));
    Span4Mux_h I__451 (
            .O(N__3111),
            .I(N__3098));
    Span4Mux_v I__450 (
            .O(N__3106),
            .I(N__3098));
    Span4Mux_h I__449 (
            .O(N__3103),
            .I(N__3095));
    Span4Mux_h I__448 (
            .O(N__3098),
            .I(N__3092));
    Odrv4 I__447 (
            .O(N__3095),
            .I(A_c_23));
    Odrv4 I__446 (
            .O(N__3092),
            .I(A_c_23));
    InMux I__445 (
            .O(N__3087),
            .I(N__3081));
    InMux I__444 (
            .O(N__3086),
            .I(N__3081));
    LocalMux I__443 (
            .O(N__3081),
            .I(N__3078));
    Span4Mux_h I__442 (
            .O(N__3078),
            .I(N__3075));
    Odrv4 I__441 (
            .O(N__3075),
            .I(\U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_3 ));
    IoInMux I__440 (
            .O(N__3072),
            .I(N__3069));
    LocalMux I__439 (
            .O(N__3069),
            .I(N__3066));
    IoSpan4Mux I__438 (
            .O(N__3066),
            .I(N__3063));
    Span4Mux_s2_v I__437 (
            .O(N__3063),
            .I(N__3060));
    Sp12to4 I__436 (
            .O(N__3060),
            .I(N__3057));
    Span12Mux_v I__435 (
            .O(N__3057),
            .I(N__3054));
    Span12Mux_h I__434 (
            .O(N__3054),
            .I(N__3051));
    Odrv12 I__433 (
            .O(N__3051),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn_i));
    IoInMux I__432 (
            .O(N__3048),
            .I(N__3045));
    LocalMux I__431 (
            .O(N__3045),
            .I(N__3042));
    IoSpan4Mux I__430 (
            .O(N__3042),
            .I(N__3039));
    Span4Mux_s2_v I__429 (
            .O(N__3039),
            .I(N__3036));
    Sp12to4 I__428 (
            .O(N__3036),
            .I(N__3033));
    Span12Mux_v I__427 (
            .O(N__3033),
            .I(N__3030));
    Odrv12 I__426 (
            .O(N__3030),
            .I(U409_ADDRESS_DECODE_un1_RAMSPACEn_i));
    InMux I__425 (
            .O(N__3027),
            .I(N__3024));
    LocalMux I__424 (
            .O(N__3024),
            .I(N__3021));
    Odrv12 I__423 (
            .O(N__3021),
            .I(\U409_ADDRESS_DECODE.un10_ROMENZ0 ));
    InMux I__422 (
            .O(N__3018),
            .I(N__3015));
    LocalMux I__421 (
            .O(N__3015),
            .I(N__3012));
    Odrv4 I__420 (
            .O(N__3012),
            .I(\U409_ADDRESS_DECODE.un1_REGSPACEnZ0 ));
    InMux I__419 (
            .O(N__3009),
            .I(N__3004));
    InMux I__418 (
            .O(N__3008),
            .I(N__3001));
    CascadeMux I__417 (
            .O(N__3007),
            .I(N__2998));
    LocalMux I__416 (
            .O(N__3004),
            .I(N__2993));
    LocalMux I__415 (
            .O(N__3001),
            .I(N__2993));
    InMux I__414 (
            .O(N__2998),
            .I(N__2990));
    Span4Mux_v I__413 (
            .O(N__2993),
            .I(N__2985));
    LocalMux I__412 (
            .O(N__2990),
            .I(N__2985));
    Span4Mux_h I__411 (
            .O(N__2985),
            .I(N__2982));
    Odrv4 I__410 (
            .O(N__2982),
            .I(\U409_ADDRESS_DECODE.un6_ROMENZ0 ));
    InMux I__409 (
            .O(N__2979),
            .I(N__2975));
    InMux I__408 (
            .O(N__2978),
            .I(N__2972));
    LocalMux I__407 (
            .O(N__2975),
            .I(N__2966));
    LocalMux I__406 (
            .O(N__2972),
            .I(N__2966));
    InMux I__405 (
            .O(N__2971),
            .I(N__2963));
    Span4Mux_v I__404 (
            .O(N__2966),
            .I(N__2960));
    LocalMux I__403 (
            .O(N__2963),
            .I(N__2957));
    Sp12to4 I__402 (
            .O(N__2960),
            .I(N__2954));
    Span12Mux_h I__401 (
            .O(N__2957),
            .I(N__2951));
    Span12Mux_h I__400 (
            .O(N__2954),
            .I(N__2948));
    Span12Mux_v I__399 (
            .O(N__2951),
            .I(N__2945));
    Span12Mux_v I__398 (
            .O(N__2948),
            .I(N__2942));
    Span12Mux_h I__397 (
            .O(N__2945),
            .I(N__2939));
    Odrv12 I__396 (
            .O(N__2942),
            .I(OVL_c));
    Odrv12 I__395 (
            .O(N__2939),
            .I(OVL_c));
    InMux I__394 (
            .O(N__2934),
            .I(N__2931));
    LocalMux I__393 (
            .O(N__2931),
            .I(N__2928));
    Span4Mux_v I__392 (
            .O(N__2928),
            .I(N__2925));
    Sp12to4 I__391 (
            .O(N__2925),
            .I(N__2922));
    Span12Mux_h I__390 (
            .O(N__2922),
            .I(N__2919));
    Odrv12 I__389 (
            .O(N__2919),
            .I(A_c_13));
    IoInMux I__388 (
            .O(N__2916),
            .I(N__2913));
    LocalMux I__387 (
            .O(N__2913),
            .I(N__2910));
    IoSpan4Mux I__386 (
            .O(N__2910),
            .I(N__2907));
    IoSpan4Mux I__385 (
            .O(N__2907),
            .I(N__2904));
    Span4Mux_s3_h I__384 (
            .O(N__2904),
            .I(N__2901));
    Sp12to4 I__383 (
            .O(N__2901),
            .I(N__2898));
    Span12Mux_s11_h I__382 (
            .O(N__2898),
            .I(N__2895));
    Odrv12 I__381 (
            .O(N__2895),
            .I(U409_ADDRESS_DECODE_un1_CIACS1n_i));
    InMux I__380 (
            .O(N__2892),
            .I(N__2889));
    LocalMux I__379 (
            .O(N__2889),
            .I(N__2886));
    Span12Mux_h I__378 (
            .O(N__2886),
            .I(N__2883));
    Odrv12 I__377 (
            .O(N__2883),
            .I(A_c_12));
    IoInMux I__376 (
            .O(N__2880),
            .I(N__2877));
    LocalMux I__375 (
            .O(N__2877),
            .I(N__2874));
    Span4Mux_s3_h I__374 (
            .O(N__2874),
            .I(N__2871));
    Span4Mux_v I__373 (
            .O(N__2871),
            .I(N__2868));
    Span4Mux_v I__372 (
            .O(N__2868),
            .I(N__2865));
    Sp12to4 I__371 (
            .O(N__2865),
            .I(N__2862));
    Span12Mux_h I__370 (
            .O(N__2862),
            .I(N__2859));
    Odrv12 I__369 (
            .O(N__2859),
            .I(U409_ADDRESS_DECODE_un1_CIACS0n_i));
    InMux I__368 (
            .O(N__2856),
            .I(N__2850));
    InMux I__367 (
            .O(N__2855),
            .I(N__2850));
    LocalMux I__366 (
            .O(N__2850),
            .I(N__2847));
    Span4Mux_h I__365 (
            .O(N__2847),
            .I(N__2844));
    Span4Mux_v I__364 (
            .O(N__2844),
            .I(N__2841));
    Odrv4 I__363 (
            .O(N__2841),
            .I(A_c_29));
    InMux I__362 (
            .O(N__2838),
            .I(N__2832));
    InMux I__361 (
            .O(N__2837),
            .I(N__2832));
    LocalMux I__360 (
            .O(N__2832),
            .I(N__2829));
    Span4Mux_v I__359 (
            .O(N__2829),
            .I(N__2826));
    Span4Mux_h I__358 (
            .O(N__2826),
            .I(N__2823));
    Odrv4 I__357 (
            .O(N__2823),
            .I(A_c_30));
    InMux I__356 (
            .O(N__2820),
            .I(N__2817));
    LocalMux I__355 (
            .O(N__2817),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3 ));
    InMux I__354 (
            .O(N__2814),
            .I(N__2810));
    CascadeMux I__353 (
            .O(N__2813),
            .I(N__2807));
    LocalMux I__352 (
            .O(N__2810),
            .I(N__2804));
    InMux I__351 (
            .O(N__2807),
            .I(N__2801));
    Span4Mux_v I__350 (
            .O(N__2804),
            .I(N__2798));
    LocalMux I__349 (
            .O(N__2801),
            .I(N__2795));
    Span4Mux_v I__348 (
            .O(N__2798),
            .I(N__2790));
    Span4Mux_v I__347 (
            .O(N__2795),
            .I(N__2790));
    Sp12to4 I__346 (
            .O(N__2790),
            .I(N__2787));
    Odrv12 I__345 (
            .O(N__2787),
            .I(A_c_25));
    InMux I__344 (
            .O(N__2784),
            .I(N__2781));
    LocalMux I__343 (
            .O(N__2781),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4 ));
    InMux I__342 (
            .O(N__2778),
            .I(N__2772));
    InMux I__341 (
            .O(N__2777),
            .I(N__2772));
    LocalMux I__340 (
            .O(N__2772),
            .I(N__2769));
    Span4Mux_v I__339 (
            .O(N__2769),
            .I(N__2766));
    Sp12to4 I__338 (
            .O(N__2766),
            .I(N__2763));
    Odrv12 I__337 (
            .O(N__2763),
            .I(A_c_27));
    InMux I__336 (
            .O(N__2760),
            .I(N__2754));
    InMux I__335 (
            .O(N__2759),
            .I(N__2754));
    LocalMux I__334 (
            .O(N__2754),
            .I(N__2751));
    Span4Mux_v I__333 (
            .O(N__2751),
            .I(N__2748));
    Span4Mux_v I__332 (
            .O(N__2748),
            .I(N__2745));
    Sp12to4 I__331 (
            .O(N__2745),
            .I(N__2742));
    Odrv12 I__330 (
            .O(N__2742),
            .I(A_c_26));
    CascadeMux I__329 (
            .O(N__2739),
            .I(N__2736));
    InMux I__328 (
            .O(N__2736),
            .I(N__2730));
    InMux I__327 (
            .O(N__2735),
            .I(N__2730));
    LocalMux I__326 (
            .O(N__2730),
            .I(N__2727));
    Span4Mux_h I__325 (
            .O(N__2727),
            .I(N__2724));
    Span4Mux_v I__324 (
            .O(N__2724),
            .I(N__2721));
    Odrv4 I__323 (
            .O(N__2721),
            .I(A_c_24));
    InMux I__322 (
            .O(N__2718),
            .I(N__2712));
    InMux I__321 (
            .O(N__2717),
            .I(N__2712));
    LocalMux I__320 (
            .O(N__2712),
            .I(N__2709));
    Span4Mux_v I__319 (
            .O(N__2709),
            .I(N__2706));
    Sp12to4 I__318 (
            .O(N__2706),
            .I(N__2703));
    Odrv12 I__317 (
            .O(N__2703),
            .I(A_c_31));
    InMux I__316 (
            .O(N__2700),
            .I(N__2697));
    LocalMux I__315 (
            .O(N__2697),
            .I(\U409_CIA.g0Z0Z_2 ));
    CascadeMux I__314 (
            .O(N__2694),
            .I(N__2690));
    InMux I__313 (
            .O(N__2693),
            .I(N__2685));
    InMux I__312 (
            .O(N__2690),
            .I(N__2685));
    LocalMux I__311 (
            .O(N__2685),
            .I(N__2682));
    Span4Mux_v I__310 (
            .O(N__2682),
            .I(N__2679));
    Span4Mux_v I__309 (
            .O(N__2679),
            .I(N__2676));
    Sp12to4 I__308 (
            .O(N__2676),
            .I(N__2673));
    Odrv12 I__307 (
            .O(N__2673),
            .I(A_c_28));
    CascadeMux I__306 (
            .O(N__2670),
            .I(\U409_CIA.g0Z0Z_10_cascade_ ));
    InMux I__305 (
            .O(N__2667),
            .I(N__2661));
    InMux I__304 (
            .O(N__2666),
            .I(N__2656));
    InMux I__303 (
            .O(N__2665),
            .I(N__2656));
    InMux I__302 (
            .O(N__2664),
            .I(N__2653));
    LocalMux I__301 (
            .O(N__2661),
            .I(N__2645));
    LocalMux I__300 (
            .O(N__2656),
            .I(N__2645));
    LocalMux I__299 (
            .O(N__2653),
            .I(N__2645));
    InMux I__298 (
            .O(N__2652),
            .I(N__2642));
    Span4Mux_v I__297 (
            .O(N__2645),
            .I(N__2637));
    LocalMux I__296 (
            .O(N__2642),
            .I(N__2637));
    Sp12to4 I__295 (
            .O(N__2637),
            .I(N__2634));
    Span12Mux_v I__294 (
            .O(N__2634),
            .I(N__2631));
    Odrv12 I__293 (
            .O(N__2631),
            .I(A_c_22));
    CascadeMux I__292 (
            .O(N__2628),
            .I(N__2625));
    InMux I__291 (
            .O(N__2625),
            .I(N__2622));
    LocalMux I__290 (
            .O(N__2622),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2 ));
    InMux I__289 (
            .O(N__2619),
            .I(N__2616));
    LocalMux I__288 (
            .O(N__2616),
            .I(N__2611));
    InMux I__287 (
            .O(N__2615),
            .I(N__2606));
    InMux I__286 (
            .O(N__2614),
            .I(N__2606));
    Span4Mux_v I__285 (
            .O(N__2611),
            .I(N__2603));
    LocalMux I__284 (
            .O(N__2606),
            .I(N__2600));
    Sp12to4 I__283 (
            .O(N__2603),
            .I(N__2597));
    Span4Mux_h I__282 (
            .O(N__2600),
            .I(N__2594));
    Span12Mux_h I__281 (
            .O(N__2597),
            .I(N__2589));
    Sp12to4 I__280 (
            .O(N__2594),
            .I(N__2589));
    Span12Mux_v I__279 (
            .O(N__2589),
            .I(N__2586));
    Odrv12 I__278 (
            .O(N__2586),
            .I(A_c_19));
    InMux I__277 (
            .O(N__2583),
            .I(N__2580));
    LocalMux I__276 (
            .O(N__2580),
            .I(N__2577));
    Span4Mux_v I__275 (
            .O(N__2577),
            .I(N__2574));
    Odrv4 I__274 (
            .O(N__2574),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3 ));
    CascadeMux I__273 (
            .O(N__2571),
            .I(\U409_ADDRESS_DECODE.un1_REGSPACEnZ0_cascade_ ));
    InMux I__272 (
            .O(N__2568),
            .I(N__2562));
    InMux I__271 (
            .O(N__2567),
            .I(N__2562));
    LocalMux I__270 (
            .O(N__2562),
            .I(N__2559));
    Span4Mux_v I__269 (
            .O(N__2559),
            .I(N__2556));
    Span4Mux_v I__268 (
            .O(N__2556),
            .I(N__2553));
    Span4Mux_v I__267 (
            .O(N__2553),
            .I(N__2550));
    Sp12to4 I__266 (
            .O(N__2550),
            .I(N__2547));
    Odrv12 I__265 (
            .O(N__2547),
            .I(A_c_18));
    CascadeMux I__264 (
            .O(N__2544),
            .I(N__2540));
    CascadeMux I__263 (
            .O(N__2543),
            .I(N__2537));
    InMux I__262 (
            .O(N__2540),
            .I(N__2532));
    InMux I__261 (
            .O(N__2537),
            .I(N__2532));
    LocalMux I__260 (
            .O(N__2532),
            .I(N__2529));
    Span4Mux_h I__259 (
            .O(N__2529),
            .I(N__2526));
    Sp12to4 I__258 (
            .O(N__2526),
            .I(N__2523));
    Span12Mux_v I__257 (
            .O(N__2523),
            .I(N__2520));
    Odrv12 I__256 (
            .O(N__2520),
            .I(A_c_16));
    InMux I__255 (
            .O(N__2517),
            .I(N__2514));
    LocalMux I__254 (
            .O(N__2514),
            .I(\U409_CIA.g0Z0Z_11 ));
    CascadeMux I__253 (
            .O(N__2511),
            .I(N__2508));
    InMux I__252 (
            .O(N__2508),
            .I(N__2504));
    InMux I__251 (
            .O(N__2507),
            .I(N__2501));
    LocalMux I__250 (
            .O(N__2504),
            .I(N__2498));
    LocalMux I__249 (
            .O(N__2501),
            .I(N__2495));
    Span12Mux_s5_h I__248 (
            .O(N__2498),
            .I(N__2490));
    Sp12to4 I__247 (
            .O(N__2495),
            .I(N__2490));
    Span12Mux_v I__246 (
            .O(N__2490),
            .I(N__2487));
    Odrv12 I__245 (
            .O(N__2487),
            .I(A_c_17));
    CascadeMux I__244 (
            .O(N__2484),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2_cascade_ ));
    InMux I__243 (
            .O(N__2481),
            .I(N__2475));
    InMux I__242 (
            .O(N__2480),
            .I(N__2475));
    LocalMux I__241 (
            .O(N__2475),
            .I(N__2472));
    Odrv4 I__240 (
            .O(N__2472),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEm_6 ));
    InMux I__239 (
            .O(N__2469),
            .I(N__2466));
    LocalMux I__238 (
            .O(N__2466),
            .I(N__2462));
    CascadeMux I__237 (
            .O(N__2465),
            .I(N__2459));
    Span4Mux_v I__236 (
            .O(N__2462),
            .I(N__2455));
    InMux I__235 (
            .O(N__2459),
            .I(N__2450));
    InMux I__234 (
            .O(N__2458),
            .I(N__2450));
    Sp12to4 I__233 (
            .O(N__2455),
            .I(N__2445));
    LocalMux I__232 (
            .O(N__2450),
            .I(N__2445));
    Odrv12 I__231 (
            .O(N__2445),
            .I(A_c_20));
    InMux I__230 (
            .O(N__2442),
            .I(N__2439));
    LocalMux I__229 (
            .O(N__2439),
            .I(N__2436));
    Odrv4 I__228 (
            .O(N__2436),
            .I(\U409_CIA.g0Z0Z_8 ));
    InMux I__227 (
            .O(N__2433),
            .I(N__2423));
    InMux I__226 (
            .O(N__2432),
            .I(N__2423));
    InMux I__225 (
            .O(N__2431),
            .I(N__2423));
    InMux I__224 (
            .O(N__2430),
            .I(N__2420));
    LocalMux I__223 (
            .O(N__2423),
            .I(N__2415));
    LocalMux I__222 (
            .O(N__2420),
            .I(N__2415));
    Span4Mux_v I__221 (
            .O(N__2415),
            .I(N__2412));
    Span4Mux_h I__220 (
            .O(N__2412),
            .I(N__2409));
    Odrv4 I__219 (
            .O(N__2409),
            .I(A_c_21));
    ClkMux I__218 (
            .O(N__2406),
            .I(N__2373));
    ClkMux I__217 (
            .O(N__2405),
            .I(N__2373));
    ClkMux I__216 (
            .O(N__2404),
            .I(N__2373));
    ClkMux I__215 (
            .O(N__2403),
            .I(N__2373));
    ClkMux I__214 (
            .O(N__2402),
            .I(N__2373));
    ClkMux I__213 (
            .O(N__2401),
            .I(N__2373));
    ClkMux I__212 (
            .O(N__2400),
            .I(N__2373));
    ClkMux I__211 (
            .O(N__2399),
            .I(N__2373));
    ClkMux I__210 (
            .O(N__2398),
            .I(N__2373));
    ClkMux I__209 (
            .O(N__2397),
            .I(N__2373));
    ClkMux I__208 (
            .O(N__2396),
            .I(N__2373));
    GlobalMux I__207 (
            .O(N__2373),
            .I(CLK80_OUT));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ),
            .I(N__2403));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .I(N__2399));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .I(N__2402));
    INV \INVU409_TRANSFER_ACK.LASTCLK_0C  (
            .O(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .I(N__2397));
    INV \INVU409_TRANSFER_ACK.TACK_EN_iC  (
            .O(\INVU409_TRANSFER_ACK.TACK_EN_iC_net ),
            .I(N__2405));
    INV \INVU409_TRANSFER_ACK.TACK_COUNTER_1C  (
            .O(\INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ),
            .I(N__2404));
    INV \INVU409_TRANSFER_ACK.CIA_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .I(N__2401));
    INV \INVU409_TRANSFER_ACK.LASTCLK_1C  (
            .O(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .I(N__2398));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .I(N__2396));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .I(N__2406));
    INV \INVU409_TRANSFER_ACK.CIA_ENABLED_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .I(N__2400));
    defparam IN_MUX_bfv_10_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_6_0_));
    defparam IN_MUX_bfv_10_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_7_0_ (
            .carryinitin(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .carryinitout(bfn_10_7_0_));
    defparam IN_MUX_bfv_12_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_6_0_));
    defparam IN_MUX_bfv_12_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_7_0_ (
            .carryinitin(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .carryinitout(bfn_12_7_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_9_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U409_CIA.g0_11_LC_1_9_0 .C_ON=1'b0;
    defparam \U409_CIA.g0_11_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_11_LC_1_9_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_CIA.g0_11_LC_1_9_0  (
            .in0(N__2615),
            .in1(N__2814),
            .in2(N__2544),
            .in3(N__2568),
            .lcout(\U409_CIA.g0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_1_9_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_1_9_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_1_9_6  (
            .in0(N__2614),
            .in1(N__2567),
            .in2(N__2543),
            .in3(N__2507),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEm_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_14_LC_1_10_3 .C_ON=1'b0;
    defparam \U409_CIA.g0_14_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_14_LC_1_10_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_CIA.g0_14_LC_1_10_3  (
            .in0(N__2517),
            .in1(N__2469),
            .in2(N__2511),
            .in3(N__2442),
            .lcout(\U409_CIA.g0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_1_12_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_1_12_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(N__2431),
            .in2(_gnd_net_),
            .in3(N__2458),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2 ),
            .ltout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_1_12_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_1_12_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_1_12_4  (
            .in0(N__3213),
            .in1(N__2480),
            .in2(N__2484),
            .in3(N__2665),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_3_LC_1_12_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_3_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_3_LC_1_12_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_3_LC_1_12_6  (
            .in0(N__2432),
            .in1(N__2481),
            .in2(N__2465),
            .in3(N__2666),
            .lcout(\U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_8_LC_1_12_7 .C_ON=1'b0;
    defparam \U409_CIA.g0_8_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_8_LC_1_12_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_CIA.g0_8_LC_1_12_7  (
            .in0(N__5541),
            .in1(N__3130),
            .in2(_gnd_net_),
            .in3(N__2433),
            .lcout(\U409_CIA.g0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un6_ROMEN_LC_1_13_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un6_ROMEN_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un6_ROMEN_LC_1_13_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_ADDRESS_DECODE.un6_ROMEN_LC_1_13_3  (
            .in0(N__2664),
            .in1(N__3129),
            .in2(_gnd_net_),
            .in3(N__2430),
            .lcout(\U409_ADDRESS_DECODE.un6_ROMENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_0  (
            .in0(N__2820),
            .in1(N__2855),
            .in2(N__2694),
            .in3(N__2784),
            .lcout(U409_ADDRESS_DECODE_Z2_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_2_LC_1_17_1 .C_ON=1'b0;
    defparam \U409_CIA.g0_2_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_2_LC_1_17_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_CIA.g0_2_LC_1_17_1  (
            .in0(N__2856),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2838),
            .lcout(\U409_CIA.g0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_17_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_17_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_17_2  (
            .in0(N__2837),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2717),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_5  (
            .in0(N__2759),
            .in1(N__2777),
            .in2(N__2813),
            .in3(N__2735),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_10_LC_1_17_6 .C_ON=1'b0;
    defparam \U409_CIA.g0_10_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_10_LC_1_17_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_CIA.g0_10_LC_1_17_6  (
            .in0(N__2778),
            .in1(N__2760),
            .in2(N__2739),
            .in3(N__2718),
            .lcout(),
            .ltout(\U409_CIA.g0Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_13_LC_1_17_7 .C_ON=1'b0;
    defparam \U409_CIA.g0_13_LC_1_17_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_13_LC_1_17_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_CIA.g0_13_LC_1_17_7  (
            .in0(N__2700),
            .in1(N__2693),
            .in2(N__2670),
            .in3(N__2652),
            .lcout(\U409_CIA.g0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un10_ROMEN_LC_2_12_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un10_ROMEN_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un10_ROMEN_LC_2_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un10_ROMEN_LC_2_12_2  (
            .in0(N__3138),
            .in1(N__2667),
            .in2(N__2628),
            .in3(N__2619),
            .lcout(\U409_ADDRESS_DECODE.un10_ROMENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_5_13_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_5_13_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_5_13_3  (
            .in0(N__3140),
            .in1(N__3225),
            .in2(_gnd_net_),
            .in3(N__3086),
            .lcout(\U409_ADDRESS_DECODE.un1_REGSPACEnZ0 ),
            .ltout(\U409_ADDRESS_DECODE.un1_REGSPACEnZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_5_13_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_5_13_4 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_5_13_4  (
            .in0(N__2583),
            .in1(N__3139),
            .in2(N__2571),
            .in3(N__5537),
            .lcout(PORTSIZE_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_5_13_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_5_13_7 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_5_13_7  (
            .in0(N__3141),
            .in1(N__3226),
            .in2(_gnd_net_),
            .in3(N__3087),
            .lcout(U409_ADDRESS_DECODE_un1_REGSPACEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_RNO_0_LC_7_8_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_RNO_0_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_RNO_0_LC_7_8_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_RNO_0_LC_7_8_2  (
            .in0(N__5504),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.RESETn_c_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_7_11_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_7_11_4 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_7_11_4  (
            .in0(N__2971),
            .in1(N__3245),
            .in2(_gnd_net_),
            .in3(N__3009),
            .lcout(U409_ADDRESS_DECODE_un1_RAMSPACEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_ROMEN_LC_7_12_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_ROMEN_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_ROMEN_LC_7_12_6 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \U409_ADDRESS_DECODE.un1_ROMEN_LC_7_12_6  (
            .in0(N__3008),
            .in1(N__3027),
            .in2(_gnd_net_),
            .in3(N__2978),
            .lcout(U409_ADDRESS_DECODE_un1_ROMEN_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_7_13_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_7_13_0 .LUT_INIT=16'b0101010100010101;
    LogicCell40 \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_7_13_0  (
            .in0(N__3018),
            .in1(N__3227),
            .in2(N__3007),
            .in3(N__2979),
            .lcout(BUFENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_8_4_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_8_4_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_8_4_7 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_8_4_7  (
            .in0(N__2934),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3405),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS1n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_8_5_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_8_5_3 .LUT_INIT=16'b1101110111011101;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_8_5_3  (
            .in0(N__3404),
            .in1(N__2892),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS0n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_8_8_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_8_8_7 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_8_8_7  (
            .in0(N__3356),
            .in1(N__3390),
            .in2(N__4320),
            .in3(N__3318),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .ce(),
            .sr(N__3414));
    defparam \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_8_9_2 .C_ON=1'b0;
    defparam \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_8_9_2 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_8_9_2  (
            .in0(N__3317),
            .in1(N__4312),
            .in2(N__3386),
            .in3(N__3357),
            .lcout(CIA_ENABLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_HOLD_LC_8_9_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_HOLD_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_HOLD_LC_8_9_7 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U409_CIA.CIA_HOLD_LC_8_9_7  (
            .in0(N__3379),
            .in1(N__3349),
            .in2(N__4316),
            .in3(N__3316),
            .lcout(\U409_CIA.CIA_HOLDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5643),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_8_11_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_8_11_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_8_11_0 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_8_11_0  (
            .in0(N__3266),
            .in1(N__5522),
            .in2(N__3291),
            .in3(N__3252),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa_0_LC_8_11_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa_0_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa_0_LC_8_11_1 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa_0_LC_8_11_1  (
            .in0(N__5524),
            .in1(N__3192),
            .in2(N__4599),
            .in3(N__3246),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0 ),
            .ltout(\U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_8_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_8_11_2 .LUT_INIT=16'b1000100110011001;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_8_11_2  (
            .in0(N__3265),
            .in1(N__3290),
            .in2(N__3303),
            .in3(N__4679),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_8_11_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_8_11_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_8_11_3 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_LC_8_11_3  (
            .in0(N__5525),
            .in1(N__3285),
            .in2(N__3300),
            .in3(N__3540),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_8_11_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_8_11_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_8_11_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_8_11_5  (
            .in0(N__5523),
            .in1(N__3286),
            .in2(_gnd_net_),
            .in3(N__3267),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_8_11_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_8_11_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_8_11_7  (
            .in0(N__3297),
            .in1(N__3284),
            .in2(N__4687),
            .in3(N__3264),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMENm_i_LC_8_12_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMENm_i_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMENm_i_LC_8_12_3 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \U409_ADDRESS_DECODE.ROMENm_i_LC_8_12_3  (
            .in0(N__3244),
            .in1(N__3191),
            .in2(_gnd_net_),
            .in3(N__5529),
            .lcout(ROMENm_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_9_7_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_9_7_2 .LUT_INIT=16'b0001000000011111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_9_7_2  (
            .in0(N__3431),
            .in1(N__3455),
            .in2(N__3629),
            .in3(N__3642),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.m9_bm_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_9_7_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_9_7_3 .LUT_INIT=16'b0000100000101010;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_0_LC_9_7_3  (
            .in0(N__5435),
            .in1(N__3666),
            .in2(N__3486),
            .in3(N__3480),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_9_8_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_9_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_9_8_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_1_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__5513),
            .in2(_gnd_net_),
            .in3(N__3822),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_9_8_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_9_8_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__3473),
            .in2(_gnd_net_),
            .in3(N__3820),
            .lcout(\U409_TRANSFER_ACK.N_4 ),
            .ltout(\U409_TRANSFER_ACK.N_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_9_8_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_9_8_3 .LUT_INIT=16'b1011000111110101;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_9_8_3  (
            .in0(N__3618),
            .in1(N__3430),
            .in2(N__3483),
            .in3(N__3453),
            .lcout(\U409_TRANSFER_ACK.m9_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_9_8_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_9_8_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_9_8_4  (
            .in0(N__3662),
            .in1(N__3474),
            .in2(N__4683),
            .in3(N__3821),
            .lcout(\U409_TRANSFER_ACK.N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_9_8_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_9_8_5 .LUT_INIT=16'b0000010100110011;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_9_8_5  (
            .in0(N__3456),
            .in1(N__3465),
            .in2(N__3435),
            .in3(N__3663),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.i6_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_9_8_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_9_8_6 .LUT_INIT=16'b0000110010001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_1_LC_9_8_6  (
            .in0(N__3664),
            .in1(N__5512),
            .in2(N__3459),
            .in3(N__3619),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_9_8_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_9_8_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_9_8_7  (
            .in0(N__5511),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3454),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_9_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_9_9_6 .LUT_INIT=16'b0001101100001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_9_9_6  (
            .in0(N__3665),
            .in1(N__3641),
            .in2(N__3630),
            .in3(N__3567),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.CIA_TACK_EN_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_9_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_9_9_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_LC_9_9_7  (
            .in0(N__5514),
            .in1(_gnd_net_),
            .in2(N__3600),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_9_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_9_10_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_9_10_0  (
            .in0(N__5516),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3525),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_9_10_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_9_10_2 .LUT_INIT=16'b0000110011101100;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_LC_9_10_2  (
            .in0(N__3555),
            .in1(N__3578),
            .in2(N__5533),
            .in3(N__3513),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_9_10_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_9_10_4 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_9_10_4  (
            .in0(N__3554),
            .in1(N__5520),
            .in2(_gnd_net_),
            .in3(N__3524),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIHST5_LC_9_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIHST5_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIHST5_LC_9_10_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNIHST5_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(N__3809),
            .in2(_gnd_net_),
            .in3(N__3566),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNIURL11_LC_9_10_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNIURL11_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNIURL11_LC_9_10_6 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNIURL11_LC_9_10_6  (
            .in0(N__3553),
            .in1(N__3523),
            .in2(N__3543),
            .in3(N__3539),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_9_10_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_9_10_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3528),
            .in3(N__5515),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_9_11_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_9_11_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_9_11_0 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_i_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__5521),
            .in2(_gnd_net_),
            .in3(N__3512),
            .lcout(TACK_EN_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_EN_iC_net ),
            .ce(N__3501),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_6_LC_10_5_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_6_LC_10_5_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_6_LC_10_5_1 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \U409_TICK.COUNTER60_6_LC_10_5_1  (
            .in0(N__4090),
            .in1(N__3735),
            .in2(N__4026),
            .in3(N__4062),
            .lcout(\U409_TICK.COUNTER60Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5301),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_8_LC_10_5_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_8_LC_10_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_8_LC_10_5_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_8_LC_10_5_2  (
            .in0(N__4013),
            .in1(N__4091),
            .in2(N__4065),
            .in3(N__3708),
            .lcout(\U409_TICK.COUNTER60Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5301),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_10_5_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_10_5_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_10_5_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER60_RNIDB4S_16_LC_10_5_3  (
            .in0(N__3873),
            .in1(N__3681),
            .in2(N__3840),
            .in3(N__3935),
            .lcout(),
            .ltout(\U409_TICK.TICK603_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_10_5_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_10_5_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_10_5_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER60_RNI335G2_11_LC_10_5_4  (
            .in0(N__3687),
            .in1(N__3891),
            .in2(N__3693),
            .in3(N__3798),
            .lcout(\U409_TICK.TICK603_14 ),
            .ltout(\U409_TICK.TICK603_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_4_LC_10_5_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_4_LC_10_5_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_4_LC_10_5_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_4_LC_10_5_5  (
            .in0(N__4089),
            .in1(N__4058),
            .in2(N__3690),
            .in3(N__3771),
            .lcout(\U409_TICK.COUNTER60Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5301),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_10_5_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_10_5_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_10_5_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_TICK.COUNTER60_RNIHJU51_4_LC_10_5_6  (
            .in0(N__3762),
            .in1(N__3783),
            .in2(_gnd_net_),
            .in3(N__3912),
            .lcout(\U409_TICK.TICK603_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_10_5_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_10_5_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_10_5_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER60_RNICDC71_14_LC_10_5_7  (
            .in0(N__3747),
            .in1(N__4167),
            .in2(N__3723),
            .in3(N__4239),
            .lcout(\U409_TICK.TICK603_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_10_6_0 .C_ON=1'b1;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_10_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_10_6_0  (
            .in0(_gnd_net_),
            .in1(N__3934),
            .in2(N__3917),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_6_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_2_LC_10_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_2_LC_10_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_2_LC_10_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_2_LC_10_6_1  (
            .in0(_gnd_net_),
            .in1(N__3680),
            .in2(_gnd_net_),
            .in3(N__3669),
            .lcout(\U409_TICK.COUNTER60Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .clk(N__5304),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_3_LC_10_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_3_LC_10_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_3_LC_10_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_3_LC_10_6_2  (
            .in0(_gnd_net_),
            .in1(N__3797),
            .in2(_gnd_net_),
            .in3(N__3786),
            .lcout(\U409_TICK.COUNTER60Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .clk(N__5304),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_10_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_10_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_4_LC_10_6_3  (
            .in0(_gnd_net_),
            .in1(N__3782),
            .in2(_gnd_net_),
            .in3(N__3765),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_5_LC_10_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_5_LC_10_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_5_LC_10_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_5_LC_10_6_4  (
            .in0(_gnd_net_),
            .in1(N__3761),
            .in2(_gnd_net_),
            .in3(N__3750),
            .lcout(\U409_TICK.COUNTER60Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .clk(N__5304),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_10_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_10_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_6_LC_10_6_5  (
            .in0(_gnd_net_),
            .in1(N__3746),
            .in2(_gnd_net_),
            .in3(N__3729),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_7_LC_10_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_7_LC_10_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_7_LC_10_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_7_LC_10_6_6  (
            .in0(_gnd_net_),
            .in1(N__4124),
            .in2(_gnd_net_),
            .in3(N__3726),
            .lcout(\U409_TICK.COUNTER60Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .clk(N__5304),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_10_6_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_10_6_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_10_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_8_LC_10_6_7  (
            .in0(_gnd_net_),
            .in1(N__3719),
            .in2(_gnd_net_),
            .in3(N__3702),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_10_7_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_10_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_9_LC_10_7_0  (
            .in0(_gnd_net_),
            .in1(N__4166),
            .in2(_gnd_net_),
            .in3(N__3699),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_10_7_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_10_LC_10_7_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_10_LC_10_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_10_LC_10_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_10_LC_10_7_1  (
            .in0(_gnd_net_),
            .in1(N__4142),
            .in2(_gnd_net_),
            .in3(N__3696),
            .lcout(\U409_TICK.COUNTER60Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .clk(N__5306),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_11_LC_10_7_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_11_LC_10_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_11_LC_10_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_11_LC_10_7_2  (
            .in0(_gnd_net_),
            .in1(N__3887),
            .in2(_gnd_net_),
            .in3(N__3876),
            .lcout(\U409_TICK.COUNTER60Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .clk(N__5306),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_12_LC_10_7_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_12_LC_10_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_12_LC_10_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_12_LC_10_7_3  (
            .in0(_gnd_net_),
            .in1(N__3869),
            .in2(_gnd_net_),
            .in3(N__3855),
            .lcout(\U409_TICK.COUNTER60Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .clk(N__5306),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_13_LC_10_7_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_13_LC_10_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_13_LC_10_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_13_LC_10_7_4  (
            .in0(_gnd_net_),
            .in1(N__4154),
            .in2(_gnd_net_),
            .in3(N__3852),
            .lcout(\U409_TICK.COUNTER60Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .clk(N__5306),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_10_7_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_10_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_14_LC_10_7_5  (
            .in0(_gnd_net_),
            .in1(N__4238),
            .in2(_gnd_net_),
            .in3(N__3849),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_10_7_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_10_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_15_LC_10_7_6  (
            .in0(_gnd_net_),
            .in1(N__4112),
            .in2(_gnd_net_),
            .in3(N__3846),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_16_LC_10_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_16_LC_10_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_16_LC_10_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER60_16_LC_10_7_7  (
            .in0(_gnd_net_),
            .in1(N__3836),
            .in2(_gnd_net_),
            .in3(N__3843),
            .lcout(\U409_TICK.COUNTER60Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5306),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_10_8_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_10_8_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_10_8_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_0_LC_10_8_6  (
            .in0(_gnd_net_),
            .in1(N__5468),
            .in2(_gnd_net_),
            .in3(N__4256),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_10_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_10_0 .LUT_INIT=16'b0000000001110101;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_10_0  (
            .in0(N__4539),
            .in1(N__4597),
            .in2(N__4688),
            .in3(N__4797),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5367));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_10_10_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_10_10_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_10_10_1 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_10_10_1  (
            .in0(N__3810),
            .in1(N__4538),
            .in2(_gnd_net_),
            .in3(N__4553),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5367));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_10_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_10_4 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_10_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_10_4  (
            .in0(N__4798),
            .in1(N__3967),
            .in2(_gnd_net_),
            .in3(N__4764),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5367));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_10_11_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_10_11_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_10_11_0  (
            .in0(N__4761),
            .in1(N__4514),
            .in2(N__3968),
            .in3(N__4795),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_10_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_10_11_2 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_10_11_2  (
            .in0(N__4762),
            .in1(_gnd_net_),
            .in2(N__3969),
            .in3(N__4796),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_10_11_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_10_11_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_10_11_3  (
            .in0(N__4710),
            .in1(N__4513),
            .in2(N__4800),
            .in3(N__4738),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_10_11_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_10_11_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_10_11_4  (
            .in0(N__4998),
            .in1(N__5022),
            .in2(N__3975),
            .in3(N__3944),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_10_11_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_10_11_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_10_11_5  (
            .in0(N__5021),
            .in1(N__4512),
            .in2(N__5004),
            .in3(N__4739),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_10_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_10_11_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_10_11_6  (
            .in0(N__4711),
            .in1(N__4794),
            .in2(N__3972),
            .in3(N__3945),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_11_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_11_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_11_7  (
            .in0(_gnd_net_),
            .in1(N__4760),
            .in2(_gnd_net_),
            .in3(N__3960),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_1_LC_11_5_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_1_LC_11_5_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_1_LC_11_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_TICK.COUNTER60_1_LC_11_5_1  (
            .in0(_gnd_net_),
            .in1(N__3913),
            .in2(_gnd_net_),
            .in3(N__3936),
            .lcout(\U409_TICK.COUNTER60Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5299),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_0_LC_11_5_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_0_LC_11_5_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_0_LC_11_5_4 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U409_TICK.COUNTER60_0_LC_11_5_4  (
            .in0(N__4095),
            .in1(N__4063),
            .in2(N__3918),
            .in3(N__4014),
            .lcout(\U409_TICK.COUNTER60Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5299),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK60_LC_11_5_6 .C_ON=1'b0;
    defparam \U409_TICK.TICK60_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK60_LC_11_5_6 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \U409_TICK.TICK60_LC_11_5_6  (
            .in0(N__4015),
            .in1(N__4064),
            .in2(N__4100),
            .in3(N__4193),
            .lcout(TICK60_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5299),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_5_LC_11_6_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_5_LC_11_6_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_5_LC_11_6_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_5_LC_11_6_0  (
            .in0(N__4421),
            .in1(N__4454),
            .in2(N__4389),
            .in3(N__4854),
            .lcout(\U409_TICK.COUNTER50Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5302),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_6_LC_11_6_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_6_LC_11_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_6_LC_11_6_1 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \U409_TICK.COUNTER50_6_LC_11_6_1  (
            .in0(N__4833),
            .in1(N__4422),
            .in2(N__4458),
            .in3(N__4387),
            .lcout(\U409_TICK.COUNTER50Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5302),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_1_LC_11_6_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_1_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_1_LC_11_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_TICK.COUNTER50_1_LC_11_6_2  (
            .in0(_gnd_net_),
            .in1(N__4961),
            .in2(_gnd_net_),
            .in3(N__4943),
            .lcout(\U409_TICK.COUNTER50Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5302),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_11_6_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_11_6_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER50_RNIUHF01_16_LC_11_6_3  (
            .in0(N__5193),
            .in1(N__4920),
            .in2(N__4962),
            .in3(N__5318),
            .lcout(\U409_TICK.TICK503_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_15_LC_11_6_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_15_LC_11_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_15_LC_11_6_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_15_LC_11_6_4  (
            .in0(N__4027),
            .in1(N__4057),
            .in2(N__4101),
            .in3(N__4182),
            .lcout(\U409_TICK.COUNTER60Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5302),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_9_LC_11_6_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_9_LC_11_6_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_9_LC_11_6_5 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_9_LC_11_6_5  (
            .in0(N__4056),
            .in1(N__4029),
            .in2(N__4176),
            .in3(N__4099),
            .lcout(\U409_TICK.COUNTER60Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5302),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_11_6_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_11_6_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_TICK.COUNTER60_RNI2USG_10_LC_11_6_6  (
            .in0(N__4155),
            .in1(N__4143),
            .in2(N__4131),
            .in3(N__4113),
            .lcout(\U409_TICK.TICK603_10 ),
            .ltout(\U409_TICK.TICK603_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_14_LC_11_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_14_LC_11_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_14_LC_11_6_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_14_LC_11_6_7  (
            .in0(N__4055),
            .in1(N__4028),
            .in2(N__3984),
            .in3(N__3981),
            .lcout(\U409_TICK.COUNTER60Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5302),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_11_7_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_11_7_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_TICK.COUNTER50_RNID6CP_3_LC_11_7_0  (
            .in0(N__4866),
            .in1(N__4905),
            .in2(_gnd_net_),
            .in3(N__4941),
            .lcout(),
            .ltout(\U409_TICK.TICK503_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_11_7_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_11_7_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER50_RNITU182_10_LC_11_7_1  (
            .in0(N__4227),
            .in1(N__5109),
            .in2(N__4221),
            .in3(N__5151),
            .lcout(\U409_TICK.TICK503_14 ),
            .ltout(\U409_TICK.TICK503_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_14_LC_11_7_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_14_LC_11_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_14_LC_11_7_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_14_LC_11_7_2  (
            .in0(N__4415),
            .in1(N__4378),
            .in2(N__4218),
            .in3(N__5061),
            .lcout(\U409_TICK.COUNTER50Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5305),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_15_LC_11_7_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_15_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_15_LC_11_7_3 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_15_LC_11_7_3  (
            .in0(N__4377),
            .in1(N__4452),
            .in2(N__5040),
            .in3(N__4417),
            .lcout(\U409_TICK.COUNTER50Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5305),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_11_7_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_11_7_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNII24V_14_LC_11_7_4  (
            .in0(N__5073),
            .in1(N__4824),
            .in2(N__4890),
            .in3(N__5052),
            .lcout(\U409_TICK.TICK503_10 ),
            .ltout(\U409_TICK.TICK503_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_13_LC_11_7_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_13_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_13_LC_11_7_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_13_LC_11_7_5  (
            .in0(N__4376),
            .in1(N__4451),
            .in2(N__4215),
            .in3(N__5082),
            .lcout(\U409_TICK.COUNTER50Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5305),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_11_7_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_11_7_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNIH14V_11_LC_11_7_6  (
            .in0(N__5094),
            .in1(N__4845),
            .in2(N__5136),
            .in3(N__5175),
            .lcout(\U409_TICK.TICK503_9 ),
            .ltout(\U409_TICK.TICK503_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_0_LC_11_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_0_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_0_LC_11_7_7 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \U409_TICK.COUNTER50_0_LC_11_7_7  (
            .in0(N__4942),
            .in1(N__4416),
            .in2(N__4212),
            .in3(N__4453),
            .lcout(\U409_TICK.COUNTER50Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5305),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_11_LC_11_8_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_11_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_11_LC_11_8_3 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_11_LC_11_8_3  (
            .in0(N__4418),
            .in1(N__4449),
            .in2(N__5121),
            .in3(N__4382),
            .lcout(\U409_TICK.COUNTER50Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5307),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_9_LC_11_8_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_9_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_9_LC_11_8_5 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_9_LC_11_8_5  (
            .in0(N__4419),
            .in1(N__4383),
            .in2(N__5163),
            .in3(N__4450),
            .lcout(\U409_TICK.COUNTER50Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5307),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK50_LC_11_8_6 .C_ON=1'b0;
    defparam \U409_TICK.TICK50_LC_11_8_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK50_LC_11_8_6 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \U409_TICK.TICK50_LC_11_8_6  (
            .in0(N__4448),
            .in1(N__4420),
            .in2(N__4388),
            .in3(N__4334),
            .lcout(TICK50_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5307),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_RNO_1_LC_11_9_0 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_RNO_1_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLKCIA_RNO_1_LC_11_9_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_CIA.CLKCIA_RNO_1_LC_11_9_0  (
            .in0(N__5259),
            .in1(N__5216),
            .in2(N__5751),
            .in3(N__5673),
            .lcout(\U409_CIA.CLKCIA6_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_11_9_1 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_11_9_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_1_LC_11_9_1  (
            .in0(N__5240),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5711),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5641),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_0_LC_11_9_2 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_0_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_0_LC_11_9_2 .LUT_INIT=16'b0100010000100010;
    LogicCell40 \U409_CIA.VMA_RNO_0_LC_11_9_2  (
            .in0(N__5671),
            .in1(N__5708),
            .in2(_gnd_net_),
            .in3(N__5239),
            .lcout(),
            .ltout(\U409_CIA.N_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_LC_11_9_3 .C_ON=1'b0;
    defparam \U409_CIA.VMA_LC_11_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.VMA_LC_11_9_3 .LUT_INIT=16'b0011101010101010;
    LogicCell40 \U409_CIA.VMA_LC_11_9_3  (
            .in0(N__4308),
            .in1(N__5672),
            .in2(N__4323),
            .in3(N__4809),
            .lcout(\U409_CIA.VMAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5641),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_RNO_2_LC_11_9_4 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_RNO_2_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLKCIA_RNO_2_LC_11_9_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_CIA.CLKCIA_RNO_2_LC_11_9_4  (
            .in0(N__5670),
            .in1(N__5707),
            .in2(_gnd_net_),
            .in3(N__5238),
            .lcout(),
            .ltout(\U409_CIA.N_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_RNO_0_LC_11_9_5 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_RNO_0_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLKCIA_RNO_0_LC_11_9_5 .LUT_INIT=16'b1111110011001100;
    LogicCell40 \U409_CIA.CLKCIA_RNO_0_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__4255),
            .in2(N__4287),
            .in3(N__4808),
            .lcout(),
            .ltout(\U409_CIA.CLKCIAZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_LC_11_9_6 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CLKCIA_LC_11_9_6 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \U409_CIA.CLKCIA_LC_11_9_6  (
            .in0(N__4284),
            .in1(N__5709),
            .in2(N__4278),
            .in3(N__5241),
            .lcout(CLKCIA_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5641),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_11_9_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_11_9_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_11_9_7  (
            .in0(N__5745),
            .in1(N__5211),
            .in2(_gnd_net_),
            .in3(N__5258),
            .lcout(\U409_CIA.CLKCIA8_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_10_5 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_10_5 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_10_5  (
            .in0(N__4799),
            .in1(N__4763),
            .in2(_gnd_net_),
            .in3(N__4481),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__5366));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_11_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_11_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_11_0 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_11_0  (
            .in0(N__4740),
            .in1(N__4713),
            .in2(N__4725),
            .in3(N__4480),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ),
            .ce(),
            .sr(N__5365));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_11_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_11_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_11_1  (
            .in0(N__4492),
            .in1(N__4999),
            .in2(_gnd_net_),
            .in3(N__5023),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_11_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_11_2 .LUT_INIT=16'b0000000000111100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__4712),
            .in2(N__4716),
            .in3(N__4476),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ),
            .ce(),
            .sr(N__5365));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_11_11_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_11_11_3 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_11_11_3  (
            .in0(N__4652),
            .in1(N__4598),
            .in2(N__4554),
            .in3(N__4537),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_11_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_11_4 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_11_4 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_11_4  (
            .in0(N__5024),
            .in1(_gnd_net_),
            .in2(N__4524),
            .in3(N__4493),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ),
            .ce(),
            .sr(N__5365));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_11_6 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_11_6 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_11_6  (
            .in0(N__4521),
            .in1(N__4515),
            .in2(_gnd_net_),
            .in3(N__4475),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ),
            .ce(),
            .sr(N__5365));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_11_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_11_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_11_7 .LUT_INIT=16'b0000011000001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_11_7  (
            .in0(N__4494),
            .in1(N__5000),
            .in2(N__4482),
            .in3(N__5025),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ),
            .ce(),
            .sr(N__5365));
    defparam CONSTANT_ONE_LUT4_LC_12_1_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_1_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_1_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_1_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_12_6_0 .C_ON=1'b1;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_12_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(N__4957),
            .in2(N__4944),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_6_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_2_LC_12_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_2_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_2_LC_12_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_2_LC_12_6_1  (
            .in0(_gnd_net_),
            .in1(N__4919),
            .in2(_gnd_net_),
            .in3(N__4908),
            .lcout(\U409_TICK.COUNTER50Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .clk(N__5300),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_3_LC_12_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_3_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_3_LC_12_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_3_LC_12_6_2  (
            .in0(_gnd_net_),
            .in1(N__4904),
            .in2(_gnd_net_),
            .in3(N__4893),
            .lcout(\U409_TICK.COUNTER50Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .clk(N__5300),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_4_LC_12_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_4_LC_12_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_4_LC_12_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_4_LC_12_6_3  (
            .in0(_gnd_net_),
            .in1(N__4880),
            .in2(_gnd_net_),
            .in3(N__4869),
            .lcout(\U409_TICK.COUNTER50Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .clk(N__5300),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_12_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_12_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_5_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(N__4865),
            .in2(_gnd_net_),
            .in3(N__4848),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_12_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_12_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_6_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(N__4844),
            .in2(_gnd_net_),
            .in3(N__4827),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_7_LC_12_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_7_LC_12_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_7_LC_12_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_7_LC_12_6_6  (
            .in0(_gnd_net_),
            .in1(N__4823),
            .in2(_gnd_net_),
            .in3(N__4812),
            .lcout(\U409_TICK.COUNTER50Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .clk(N__5300),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_8_LC_12_6_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_8_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_8_LC_12_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_8_LC_12_6_7  (
            .in0(_gnd_net_),
            .in1(N__5189),
            .in2(_gnd_net_),
            .in3(N__5178),
            .lcout(\U409_TICK.COUNTER50Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .clk(N__5300),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_12_7_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_12_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_9_LC_12_7_0  (
            .in0(_gnd_net_),
            .in1(N__5174),
            .in2(_gnd_net_),
            .in3(N__5154),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_12_7_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_10_LC_12_7_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_10_LC_12_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_10_LC_12_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_10_LC_12_7_1  (
            .in0(_gnd_net_),
            .in1(N__5150),
            .in2(_gnd_net_),
            .in3(N__5139),
            .lcout(\U409_TICK.COUNTER50Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .clk(N__5303),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_12_7_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_12_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_11_LC_12_7_2  (
            .in0(_gnd_net_),
            .in1(N__5132),
            .in2(_gnd_net_),
            .in3(N__5112),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_12_LC_12_7_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_12_LC_12_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_12_LC_12_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_12_LC_12_7_3  (
            .in0(_gnd_net_),
            .in1(N__5108),
            .in2(_gnd_net_),
            .in3(N__5097),
            .lcout(\U409_TICK.COUNTER50Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .clk(N__5303),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_12_7_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_12_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_13_LC_12_7_4  (
            .in0(_gnd_net_),
            .in1(N__5093),
            .in2(_gnd_net_),
            .in3(N__5076),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_12_7_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_12_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_14_LC_12_7_5  (
            .in0(_gnd_net_),
            .in1(N__5072),
            .in2(_gnd_net_),
            .in3(N__5055),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_12_7_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_12_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_15_LC_12_7_6  (
            .in0(_gnd_net_),
            .in1(N__5051),
            .in2(_gnd_net_),
            .in3(N__5028),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_16_LC_12_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_16_LC_12_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_16_LC_12_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER50_16_LC_12_7_7  (
            .in0(_gnd_net_),
            .in1(N__5319),
            .in2(_gnd_net_),
            .in3(N__5322),
            .lcout(\U409_TICK.COUNTER50Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5303),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_12_8_1 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_12_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_12_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_0_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5710),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5642),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_9_0 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__5236),
            .in2(N__5712),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_12_9_1 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_12_9_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_12_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_2_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(N__5256),
            .in2(_gnd_net_),
            .in3(N__5274),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .clk(N__5640),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_12_9_2 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_12_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(N__5667),
            .in2(_gnd_net_),
            .in3(N__5271),
            .lcout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_12_9_3 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_12_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_12_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_4_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(N__5212),
            .in2(_gnd_net_),
            .in3(N__5268),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .clk(N__5640),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_12_9_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_12_9_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(N__5750),
            .in2(_gnd_net_),
            .in3(N__5265),
            .lcout(),
            .ltout(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_12_9_5 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_12_9_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_12_9_5 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_5_LC_12_9_5  (
            .in0(N__5669),
            .in1(N__5727),
            .in2(N__5262),
            .in3(N__5705),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5640),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_12_9_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_12_9_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_12_9_6  (
            .in0(N__5257),
            .in1(N__5237),
            .in2(N__5217),
            .in3(N__5749),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_0_a2_2 ),
            .ltout(\U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_12_9_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_12_9_7 .LUT_INIT=16'b0010011001100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_3_LC_12_9_7  (
            .in0(N__5668),
            .in1(N__5721),
            .in2(N__5715),
            .in3(N__5706),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5640),
            .ce(),
            .sr(_gnd_net_));
    defparam TACKn_iobuf_RNO_LC_18_13_4.C_ON=1'b0;
    defparam TACKn_iobuf_RNO_LC_18_13_4.SEQ_MODE=4'b0000;
    defparam TACKn_iobuf_RNO_LC_18_13_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 TACKn_iobuf_RNO_LC_18_13_4 (
            .in0(N__5625),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_353_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_18_13_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_18_13_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_18_13_6 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_18_13_6  (
            .in0(N__5576),
            .in1(N__5556),
            .in2(_gnd_net_),
            .in3(N__5459),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U409_TOP

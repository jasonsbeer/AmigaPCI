// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Apr 14 2025 17:39:38

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U409_TOP" view "INTERFACE"

module U409_TOP (
    TM,
    TT,
    D,
    A,
    TICK60,
    CIACS0n,
    CLK6,
    CLK_CIA,
    BUFENn,
    CIACS1n,
    TICK50,
    RAMSPACEn,
    CLK40_IN,
    CLK28_IN,
    REGSPACEn,
    TSn,
    RTC_ENn,
    RESETn,
    OVL,
    TACKn,
    ROMENn,
    PORTSIZE);

    input [1:0] TM;
    input [1:0] TT;
    output [7:0] D;
    input [31:1] A;
    output TICK60;
    output CIACS0n;
    input CLK6;
    output CLK_CIA;
    output BUFENn;
    output CIACS1n;
    output TICK50;
    output RAMSPACEn;
    input CLK40_IN;
    input CLK28_IN;
    output REGSPACEn;
    input TSn;
    output RTC_ENn;
    input RESETn;
    input OVL;
    inout TACKn;
    output ROMENn;
    output PORTSIZE;

    wire N__7448;
    wire N__7447;
    wire N__7446;
    wire N__7438;
    wire N__7437;
    wire N__7436;
    wire N__7427;
    wire N__7426;
    wire N__7425;
    wire N__7418;
    wire N__7417;
    wire N__7416;
    wire N__7409;
    wire N__7408;
    wire N__7407;
    wire N__7400;
    wire N__7399;
    wire N__7398;
    wire N__7391;
    wire N__7390;
    wire N__7389;
    wire N__7382;
    wire N__7381;
    wire N__7380;
    wire N__7373;
    wire N__7372;
    wire N__7371;
    wire N__7364;
    wire N__7363;
    wire N__7362;
    wire N__7355;
    wire N__7354;
    wire N__7353;
    wire N__7346;
    wire N__7345;
    wire N__7344;
    wire N__7337;
    wire N__7336;
    wire N__7335;
    wire N__7328;
    wire N__7327;
    wire N__7326;
    wire N__7319;
    wire N__7318;
    wire N__7317;
    wire N__7310;
    wire N__7309;
    wire N__7308;
    wire N__7301;
    wire N__7300;
    wire N__7299;
    wire N__7292;
    wire N__7291;
    wire N__7290;
    wire N__7283;
    wire N__7282;
    wire N__7281;
    wire N__7274;
    wire N__7273;
    wire N__7272;
    wire N__7265;
    wire N__7264;
    wire N__7263;
    wire N__7256;
    wire N__7255;
    wire N__7254;
    wire N__7247;
    wire N__7246;
    wire N__7245;
    wire N__7238;
    wire N__7237;
    wire N__7236;
    wire N__7229;
    wire N__7228;
    wire N__7227;
    wire N__7220;
    wire N__7219;
    wire N__7218;
    wire N__7211;
    wire N__7210;
    wire N__7209;
    wire N__7202;
    wire N__7201;
    wire N__7200;
    wire N__7193;
    wire N__7192;
    wire N__7191;
    wire N__7184;
    wire N__7183;
    wire N__7182;
    wire N__7175;
    wire N__7174;
    wire N__7173;
    wire N__7166;
    wire N__7165;
    wire N__7164;
    wire N__7157;
    wire N__7156;
    wire N__7155;
    wire N__7148;
    wire N__7147;
    wire N__7146;
    wire N__7139;
    wire N__7138;
    wire N__7137;
    wire N__7130;
    wire N__7129;
    wire N__7128;
    wire N__7121;
    wire N__7120;
    wire N__7119;
    wire N__7112;
    wire N__7111;
    wire N__7110;
    wire N__7103;
    wire N__7102;
    wire N__7101;
    wire N__7094;
    wire N__7093;
    wire N__7092;
    wire N__7085;
    wire N__7084;
    wire N__7083;
    wire N__7076;
    wire N__7075;
    wire N__7074;
    wire N__7067;
    wire N__7066;
    wire N__7065;
    wire N__7058;
    wire N__7057;
    wire N__7056;
    wire N__7049;
    wire N__7048;
    wire N__7047;
    wire N__7040;
    wire N__7039;
    wire N__7038;
    wire N__7031;
    wire N__7030;
    wire N__7029;
    wire N__7022;
    wire N__7021;
    wire N__7020;
    wire N__7003;
    wire N__7002;
    wire N__7001;
    wire N__6998;
    wire N__6997;
    wire N__6996;
    wire N__6995;
    wire N__6994;
    wire N__6989;
    wire N__6986;
    wire N__6977;
    wire N__6970;
    wire N__6969;
    wire N__6968;
    wire N__6965;
    wire N__6964;
    wire N__6963;
    wire N__6962;
    wire N__6959;
    wire N__6954;
    wire N__6947;
    wire N__6940;
    wire N__6939;
    wire N__6938;
    wire N__6931;
    wire N__6928;
    wire N__6925;
    wire N__6922;
    wire N__6919;
    wire N__6916;
    wire N__6913;
    wire N__6910;
    wire N__6907;
    wire N__6904;
    wire N__6901;
    wire N__6898;
    wire N__6895;
    wire N__6892;
    wire N__6891;
    wire N__6890;
    wire N__6887;
    wire N__6882;
    wire N__6877;
    wire N__6874;
    wire N__6873;
    wire N__6872;
    wire N__6869;
    wire N__6864;
    wire N__6859;
    wire N__6856;
    wire N__6853;
    wire N__6850;
    wire N__6847;
    wire N__6844;
    wire N__6843;
    wire N__6840;
    wire N__6837;
    wire N__6836;
    wire N__6833;
    wire N__6830;
    wire N__6827;
    wire N__6820;
    wire N__6817;
    wire N__6814;
    wire N__6811;
    wire N__6808;
    wire N__6805;
    wire N__6802;
    wire N__6799;
    wire N__6796;
    wire N__6795;
    wire N__6792;
    wire N__6789;
    wire N__6786;
    wire N__6783;
    wire N__6782;
    wire N__6777;
    wire N__6774;
    wire N__6769;
    wire N__6766;
    wire N__6765;
    wire N__6760;
    wire N__6757;
    wire N__6754;
    wire N__6753;
    wire N__6752;
    wire N__6751;
    wire N__6748;
    wire N__6745;
    wire N__6742;
    wire N__6739;
    wire N__6730;
    wire N__6729;
    wire N__6728;
    wire N__6727;
    wire N__6724;
    wire N__6721;
    wire N__6716;
    wire N__6709;
    wire N__6706;
    wire N__6703;
    wire N__6702;
    wire N__6701;
    wire N__6700;
    wire N__6699;
    wire N__6696;
    wire N__6693;
    wire N__6686;
    wire N__6679;
    wire N__6676;
    wire N__6675;
    wire N__6674;
    wire N__6671;
    wire N__6666;
    wire N__6661;
    wire N__6658;
    wire N__6655;
    wire N__6652;
    wire N__6649;
    wire N__6646;
    wire N__6643;
    wire N__6640;
    wire N__6637;
    wire N__6636;
    wire N__6633;
    wire N__6632;
    wire N__6629;
    wire N__6624;
    wire N__6619;
    wire N__6618;
    wire N__6615;
    wire N__6612;
    wire N__6607;
    wire N__6604;
    wire N__6601;
    wire N__6598;
    wire N__6597;
    wire N__6594;
    wire N__6591;
    wire N__6586;
    wire N__6583;
    wire N__6582;
    wire N__6579;
    wire N__6576;
    wire N__6571;
    wire N__6568;
    wire N__6565;
    wire N__6562;
    wire N__6561;
    wire N__6558;
    wire N__6555;
    wire N__6550;
    wire N__6547;
    wire N__6546;
    wire N__6543;
    wire N__6540;
    wire N__6535;
    wire N__6532;
    wire N__6529;
    wire N__6526;
    wire N__6525;
    wire N__6522;
    wire N__6519;
    wire N__6514;
    wire N__6511;
    wire N__6508;
    wire N__6505;
    wire N__6502;
    wire N__6499;
    wire N__6498;
    wire N__6495;
    wire N__6492;
    wire N__6487;
    wire N__6484;
    wire N__6481;
    wire N__6478;
    wire N__6475;
    wire N__6474;
    wire N__6471;
    wire N__6468;
    wire N__6463;
    wire N__6462;
    wire N__6461;
    wire N__6460;
    wire N__6459;
    wire N__6458;
    wire N__6457;
    wire N__6456;
    wire N__6439;
    wire N__6436;
    wire N__6433;
    wire N__6432;
    wire N__6429;
    wire N__6428;
    wire N__6423;
    wire N__6420;
    wire N__6415;
    wire N__6414;
    wire N__6413;
    wire N__6410;
    wire N__6409;
    wire N__6406;
    wire N__6403;
    wire N__6400;
    wire N__6397;
    wire N__6394;
    wire N__6385;
    wire N__6384;
    wire N__6381;
    wire N__6378;
    wire N__6373;
    wire N__6370;
    wire N__6369;
    wire N__6366;
    wire N__6363;
    wire N__6358;
    wire N__6355;
    wire N__6352;
    wire N__6351;
    wire N__6348;
    wire N__6345;
    wire N__6340;
    wire N__6337;
    wire N__6336;
    wire N__6333;
    wire N__6330;
    wire N__6327;
    wire N__6322;
    wire N__6319;
    wire N__6316;
    wire N__6313;
    wire N__6310;
    wire N__6307;
    wire N__6306;
    wire N__6303;
    wire N__6300;
    wire N__6295;
    wire N__6292;
    wire N__6289;
    wire N__6286;
    wire N__6283;
    wire N__6280;
    wire N__6279;
    wire N__6276;
    wire N__6273;
    wire N__6268;
    wire N__6265;
    wire N__6264;
    wire N__6261;
    wire N__6258;
    wire N__6253;
    wire N__6250;
    wire N__6249;
    wire N__6246;
    wire N__6243;
    wire N__6238;
    wire N__6235;
    wire N__6232;
    wire N__6229;
    wire N__6228;
    wire N__6225;
    wire N__6222;
    wire N__6217;
    wire N__6214;
    wire N__6213;
    wire N__6210;
    wire N__6207;
    wire N__6202;
    wire N__6199;
    wire N__6198;
    wire N__6195;
    wire N__6192;
    wire N__6187;
    wire N__6184;
    wire N__6183;
    wire N__6180;
    wire N__6177;
    wire N__6172;
    wire N__6169;
    wire N__6168;
    wire N__6165;
    wire N__6162;
    wire N__6157;
    wire N__6154;
    wire N__6151;
    wire N__6148;
    wire N__6147;
    wire N__6144;
    wire N__6141;
    wire N__6136;
    wire N__6133;
    wire N__6130;
    wire N__6127;
    wire N__6124;
    wire N__6123;
    wire N__6120;
    wire N__6117;
    wire N__6112;
    wire N__6111;
    wire N__6108;
    wire N__6107;
    wire N__6104;
    wire N__6101;
    wire N__6098;
    wire N__6091;
    wire N__6090;
    wire N__6087;
    wire N__6086;
    wire N__6085;
    wire N__6082;
    wire N__6079;
    wire N__6076;
    wire N__6073;
    wire N__6070;
    wire N__6061;
    wire N__6060;
    wire N__6057;
    wire N__6054;
    wire N__6049;
    wire N__6046;
    wire N__6045;
    wire N__6042;
    wire N__6039;
    wire N__6034;
    wire N__6031;
    wire N__6030;
    wire N__6027;
    wire N__6024;
    wire N__6019;
    wire N__6016;
    wire N__6013;
    wire N__6010;
    wire N__6007;
    wire N__6006;
    wire N__6003;
    wire N__6000;
    wire N__5995;
    wire N__5992;
    wire N__5991;
    wire N__5988;
    wire N__5985;
    wire N__5982;
    wire N__5979;
    wire N__5974;
    wire N__5971;
    wire N__5968;
    wire N__5965;
    wire N__5962;
    wire N__5959;
    wire N__5958;
    wire N__5955;
    wire N__5952;
    wire N__5947;
    wire N__5944;
    wire N__5943;
    wire N__5940;
    wire N__5937;
    wire N__5932;
    wire N__5929;
    wire N__5926;
    wire N__5923;
    wire N__5920;
    wire N__5917;
    wire N__5914;
    wire N__5911;
    wire N__5910;
    wire N__5909;
    wire N__5908;
    wire N__5907;
    wire N__5906;
    wire N__5905;
    wire N__5904;
    wire N__5895;
    wire N__5886;
    wire N__5881;
    wire N__5880;
    wire N__5879;
    wire N__5878;
    wire N__5877;
    wire N__5876;
    wire N__5875;
    wire N__5874;
    wire N__5863;
    wire N__5856;
    wire N__5851;
    wire N__5850;
    wire N__5849;
    wire N__5846;
    wire N__5845;
    wire N__5844;
    wire N__5843;
    wire N__5842;
    wire N__5833;
    wire N__5832;
    wire N__5829;
    wire N__5826;
    wire N__5823;
    wire N__5820;
    wire N__5813;
    wire N__5806;
    wire N__5803;
    wire N__5800;
    wire N__5797;
    wire N__5794;
    wire N__5791;
    wire N__5790;
    wire N__5787;
    wire N__5784;
    wire N__5779;
    wire N__5776;
    wire N__5775;
    wire N__5774;
    wire N__5773;
    wire N__5770;
    wire N__5767;
    wire N__5766;
    wire N__5765;
    wire N__5764;
    wire N__5755;
    wire N__5748;
    wire N__5743;
    wire N__5740;
    wire N__5737;
    wire N__5736;
    wire N__5735;
    wire N__5734;
    wire N__5733;
    wire N__5732;
    wire N__5731;
    wire N__5728;
    wire N__5721;
    wire N__5714;
    wire N__5707;
    wire N__5706;
    wire N__5703;
    wire N__5702;
    wire N__5701;
    wire N__5700;
    wire N__5699;
    wire N__5698;
    wire N__5689;
    wire N__5682;
    wire N__5677;
    wire N__5674;
    wire N__5671;
    wire N__5668;
    wire N__5665;
    wire N__5664;
    wire N__5661;
    wire N__5658;
    wire N__5653;
    wire N__5650;
    wire N__5649;
    wire N__5646;
    wire N__5645;
    wire N__5642;
    wire N__5641;
    wire N__5640;
    wire N__5637;
    wire N__5634;
    wire N__5631;
    wire N__5628;
    wire N__5625;
    wire N__5624;
    wire N__5621;
    wire N__5618;
    wire N__5615;
    wire N__5612;
    wire N__5609;
    wire N__5606;
    wire N__5593;
    wire N__5590;
    wire N__5587;
    wire N__5584;
    wire N__5581;
    wire N__5578;
    wire N__5575;
    wire N__5574;
    wire N__5573;
    wire N__5570;
    wire N__5569;
    wire N__5568;
    wire N__5565;
    wire N__5562;
    wire N__5555;
    wire N__5548;
    wire N__5547;
    wire N__5546;
    wire N__5545;
    wire N__5544;
    wire N__5541;
    wire N__5536;
    wire N__5533;
    wire N__5528;
    wire N__5521;
    wire N__5520;
    wire N__5519;
    wire N__5518;
    wire N__5517;
    wire N__5516;
    wire N__5515;
    wire N__5508;
    wire N__5505;
    wire N__5502;
    wire N__5497;
    wire N__5488;
    wire N__5487;
    wire N__5486;
    wire N__5485;
    wire N__5482;
    wire N__5479;
    wire N__5474;
    wire N__5467;
    wire N__5466;
    wire N__5463;
    wire N__5462;
    wire N__5459;
    wire N__5456;
    wire N__5453;
    wire N__5452;
    wire N__5449;
    wire N__5444;
    wire N__5441;
    wire N__5436;
    wire N__5433;
    wire N__5428;
    wire N__5425;
    wire N__5422;
    wire N__5419;
    wire N__5416;
    wire N__5413;
    wire N__5410;
    wire N__5407;
    wire N__5404;
    wire N__5401;
    wire N__5398;
    wire N__5395;
    wire N__5392;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5362;
    wire N__5359;
    wire N__5356;
    wire N__5353;
    wire N__5350;
    wire N__5349;
    wire N__5344;
    wire N__5341;
    wire N__5340;
    wire N__5339;
    wire N__5336;
    wire N__5335;
    wire N__5332;
    wire N__5329;
    wire N__5328;
    wire N__5325;
    wire N__5322;
    wire N__5319;
    wire N__5316;
    wire N__5313;
    wire N__5312;
    wire N__5307;
    wire N__5304;
    wire N__5301;
    wire N__5298;
    wire N__5295;
    wire N__5292;
    wire N__5291;
    wire N__5288;
    wire N__5283;
    wire N__5280;
    wire N__5279;
    wire N__5278;
    wire N__5277;
    wire N__5276;
    wire N__5273;
    wire N__5270;
    wire N__5269;
    wire N__5268;
    wire N__5267;
    wire N__5264;
    wire N__5259;
    wire N__5250;
    wire N__5249;
    wire N__5244;
    wire N__5241;
    wire N__5238;
    wire N__5235;
    wire N__5232;
    wire N__5227;
    wire N__5224;
    wire N__5219;
    wire N__5214;
    wire N__5207;
    wire N__5202;
    wire N__5199;
    wire N__5196;
    wire N__5193;
    wire N__5190;
    wire N__5185;
    wire N__5184;
    wire N__5183;
    wire N__5180;
    wire N__5175;
    wire N__5170;
    wire N__5169;
    wire N__5164;
    wire N__5161;
    wire N__5158;
    wire N__5155;
    wire N__5152;
    wire N__5151;
    wire N__5150;
    wire N__5147;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5131;
    wire N__5128;
    wire N__5125;
    wire N__5124;
    wire N__5123;
    wire N__5120;
    wire N__5119;
    wire N__5116;
    wire N__5115;
    wire N__5112;
    wire N__5109;
    wire N__5102;
    wire N__5095;
    wire N__5094;
    wire N__5093;
    wire N__5092;
    wire N__5089;
    wire N__5086;
    wire N__5081;
    wire N__5074;
    wire N__5073;
    wire N__5072;
    wire N__5069;
    wire N__5066;
    wire N__5063;
    wire N__5056;
    wire N__5055;
    wire N__5050;
    wire N__5047;
    wire N__5046;
    wire N__5045;
    wire N__5044;
    wire N__5041;
    wire N__5038;
    wire N__5035;
    wire N__5032;
    wire N__5023;
    wire N__5022;
    wire N__5021;
    wire N__5020;
    wire N__5019;
    wire N__5016;
    wire N__5013;
    wire N__5010;
    wire N__5007;
    wire N__5002;
    wire N__4993;
    wire N__4992;
    wire N__4991;
    wire N__4990;
    wire N__4987;
    wire N__4986;
    wire N__4985;
    wire N__4980;
    wire N__4977;
    wire N__4974;
    wire N__4971;
    wire N__4968;
    wire N__4957;
    wire N__4954;
    wire N__4951;
    wire N__4950;
    wire N__4945;
    wire N__4942;
    wire N__4939;
    wire N__4938;
    wire N__4935;
    wire N__4932;
    wire N__4931;
    wire N__4930;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4918;
    wire N__4913;
    wire N__4910;
    wire N__4907;
    wire N__4904;
    wire N__4901;
    wire N__4898;
    wire N__4891;
    wire N__4888;
    wire N__4885;
    wire N__4882;
    wire N__4879;
    wire N__4878;
    wire N__4875;
    wire N__4872;
    wire N__4871;
    wire N__4868;
    wire N__4865;
    wire N__4862;
    wire N__4861;
    wire N__4860;
    wire N__4859;
    wire N__4856;
    wire N__4853;
    wire N__4850;
    wire N__4847;
    wire N__4844;
    wire N__4841;
    wire N__4840;
    wire N__4837;
    wire N__4834;
    wire N__4829;
    wire N__4826;
    wire N__4823;
    wire N__4820;
    wire N__4811;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4799;
    wire N__4796;
    wire N__4789;
    wire N__4788;
    wire N__4785;
    wire N__4782;
    wire N__4777;
    wire N__4776;
    wire N__4771;
    wire N__4768;
    wire N__4765;
    wire N__4762;
    wire N__4759;
    wire N__4756;
    wire N__4753;
    wire N__4750;
    wire N__4747;
    wire N__4744;
    wire N__4741;
    wire N__4740;
    wire N__4737;
    wire N__4734;
    wire N__4731;
    wire N__4726;
    wire N__4723;
    wire N__4720;
    wire N__4719;
    wire N__4718;
    wire N__4717;
    wire N__4714;
    wire N__4711;
    wire N__4708;
    wire N__4703;
    wire N__4696;
    wire N__4695;
    wire N__4694;
    wire N__4693;
    wire N__4690;
    wire N__4689;
    wire N__4686;
    wire N__4683;
    wire N__4680;
    wire N__4675;
    wire N__4666;
    wire N__4663;
    wire N__4660;
    wire N__4657;
    wire N__4654;
    wire N__4651;
    wire N__4650;
    wire N__4647;
    wire N__4644;
    wire N__4639;
    wire N__4638;
    wire N__4635;
    wire N__4632;
    wire N__4629;
    wire N__4624;
    wire N__4621;
    wire N__4618;
    wire N__4615;
    wire N__4614;
    wire N__4611;
    wire N__4608;
    wire N__4603;
    wire N__4600;
    wire N__4599;
    wire N__4596;
    wire N__4595;
    wire N__4594;
    wire N__4589;
    wire N__4584;
    wire N__4579;
    wire N__4578;
    wire N__4577;
    wire N__4570;
    wire N__4567;
    wire N__4564;
    wire N__4563;
    wire N__4560;
    wire N__4557;
    wire N__4552;
    wire N__4551;
    wire N__4548;
    wire N__4545;
    wire N__4540;
    wire N__4539;
    wire N__4536;
    wire N__4533;
    wire N__4530;
    wire N__4525;
    wire N__4522;
    wire N__4519;
    wire N__4516;
    wire N__4513;
    wire N__4510;
    wire N__4507;
    wire N__4506;
    wire N__4505;
    wire N__4502;
    wire N__4497;
    wire N__4492;
    wire N__4491;
    wire N__4490;
    wire N__4487;
    wire N__4486;
    wire N__4483;
    wire N__4482;
    wire N__4479;
    wire N__4472;
    wire N__4469;
    wire N__4462;
    wire N__4461;
    wire N__4460;
    wire N__4459;
    wire N__4458;
    wire N__4455;
    wire N__4446;
    wire N__4441;
    wire N__4440;
    wire N__4439;
    wire N__4436;
    wire N__4431;
    wire N__4426;
    wire N__4423;
    wire N__4420;
    wire N__4417;
    wire N__4414;
    wire N__4411;
    wire N__4408;
    wire N__4405;
    wire N__4402;
    wire N__4401;
    wire N__4400;
    wire N__4395;
    wire N__4392;
    wire N__4389;
    wire N__4386;
    wire N__4383;
    wire N__4380;
    wire N__4377;
    wire N__4372;
    wire N__4371;
    wire N__4368;
    wire N__4365;
    wire N__4360;
    wire N__4359;
    wire N__4356;
    wire N__4353;
    wire N__4348;
    wire N__4345;
    wire N__4342;
    wire N__4339;
    wire N__4336;
    wire N__4333;
    wire N__4332;
    wire N__4329;
    wire N__4326;
    wire N__4323;
    wire N__4320;
    wire N__4315;
    wire N__4314;
    wire N__4313;
    wire N__4312;
    wire N__4311;
    wire N__4308;
    wire N__4305;
    wire N__4298;
    wire N__4291;
    wire N__4290;
    wire N__4289;
    wire N__4288;
    wire N__4287;
    wire N__4286;
    wire N__4283;
    wire N__4280;
    wire N__4271;
    wire N__4264;
    wire N__4261;
    wire N__4258;
    wire N__4255;
    wire N__4252;
    wire N__4249;
    wire N__4246;
    wire N__4243;
    wire N__4240;
    wire N__4237;
    wire N__4234;
    wire N__4231;
    wire N__4228;
    wire N__4225;
    wire N__4222;
    wire N__4219;
    wire N__4216;
    wire N__4213;
    wire N__4210;
    wire N__4207;
    wire N__4204;
    wire N__4201;
    wire N__4200;
    wire N__4199;
    wire N__4196;
    wire N__4193;
    wire N__4190;
    wire N__4183;
    wire N__4180;
    wire N__4177;
    wire N__4174;
    wire N__4173;
    wire N__4172;
    wire N__4169;
    wire N__4164;
    wire N__4161;
    wire N__4158;
    wire N__4153;
    wire N__4150;
    wire N__4147;
    wire N__4144;
    wire N__4141;
    wire N__4138;
    wire N__4137;
    wire N__4134;
    wire N__4131;
    wire N__4126;
    wire N__4123;
    wire N__4122;
    wire N__4119;
    wire N__4116;
    wire N__4113;
    wire N__4110;
    wire N__4105;
    wire N__4102;
    wire N__4099;
    wire N__4096;
    wire N__4095;
    wire N__4092;
    wire N__4089;
    wire N__4084;
    wire N__4081;
    wire N__4078;
    wire N__4075;
    wire N__4072;
    wire N__4069;
    wire N__4066;
    wire N__4063;
    wire N__4062;
    wire N__4061;
    wire N__4058;
    wire N__4057;
    wire N__4052;
    wire N__4049;
    wire N__4046;
    wire N__4043;
    wire N__4038;
    wire N__4033;
    wire N__4030;
    wire N__4027;
    wire N__4024;
    wire N__4021;
    wire N__4018;
    wire N__4015;
    wire N__4014;
    wire N__4011;
    wire N__4008;
    wire N__4007;
    wire N__4004;
    wire N__4001;
    wire N__4000;
    wire N__3999;
    wire N__3996;
    wire N__3991;
    wire N__3988;
    wire N__3985;
    wire N__3982;
    wire N__3977;
    wire N__3974;
    wire N__3971;
    wire N__3966;
    wire N__3961;
    wire N__3958;
    wire N__3955;
    wire N__3952;
    wire N__3949;
    wire N__3946;
    wire N__3943;
    wire N__3940;
    wire N__3937;
    wire N__3934;
    wire N__3931;
    wire N__3928;
    wire N__3925;
    wire N__3924;
    wire N__3923;
    wire N__3922;
    wire N__3921;
    wire N__3914;
    wire N__3909;
    wire N__3906;
    wire N__3903;
    wire N__3902;
    wire N__3899;
    wire N__3896;
    wire N__3893;
    wire N__3886;
    wire N__3883;
    wire N__3882;
    wire N__3879;
    wire N__3876;
    wire N__3871;
    wire N__3870;
    wire N__3869;
    wire N__3868;
    wire N__3865;
    wire N__3862;
    wire N__3857;
    wire N__3854;
    wire N__3849;
    wire N__3846;
    wire N__3843;
    wire N__3838;
    wire N__3835;
    wire N__3834;
    wire N__3833;
    wire N__3832;
    wire N__3831;
    wire N__3824;
    wire N__3819;
    wire N__3814;
    wire N__3811;
    wire N__3808;
    wire N__3805;
    wire N__3804;
    wire N__3803;
    wire N__3802;
    wire N__3799;
    wire N__3792;
    wire N__3789;
    wire N__3784;
    wire N__3781;
    wire N__3778;
    wire N__3775;
    wire N__3772;
    wire N__3769;
    wire N__3766;
    wire N__3765;
    wire N__3764;
    wire N__3763;
    wire N__3756;
    wire N__3753;
    wire N__3748;
    wire N__3745;
    wire N__3742;
    wire N__3739;
    wire N__3738;
    wire N__3735;
    wire N__3734;
    wire N__3731;
    wire N__3730;
    wire N__3729;
    wire N__3728;
    wire N__3725;
    wire N__3722;
    wire N__3719;
    wire N__3716;
    wire N__3713;
    wire N__3710;
    wire N__3697;
    wire N__3696;
    wire N__3693;
    wire N__3692;
    wire N__3689;
    wire N__3686;
    wire N__3683;
    wire N__3680;
    wire N__3673;
    wire N__3670;
    wire N__3667;
    wire N__3664;
    wire N__3661;
    wire N__3658;
    wire N__3655;
    wire N__3652;
    wire N__3649;
    wire N__3646;
    wire N__3643;
    wire N__3640;
    wire N__3639;
    wire N__3636;
    wire N__3633;
    wire N__3628;
    wire N__3627;
    wire N__3624;
    wire N__3621;
    wire N__3616;
    wire N__3613;
    wire N__3610;
    wire N__3609;
    wire N__3608;
    wire N__3605;
    wire N__3602;
    wire N__3599;
    wire N__3594;
    wire N__3591;
    wire N__3588;
    wire N__3585;
    wire N__3580;
    wire N__3579;
    wire N__3578;
    wire N__3577;
    wire N__3574;
    wire N__3571;
    wire N__3568;
    wire N__3565;
    wire N__3558;
    wire N__3555;
    wire N__3552;
    wire N__3549;
    wire N__3544;
    wire N__3541;
    wire N__3538;
    wire N__3535;
    wire N__3532;
    wire N__3531;
    wire N__3528;
    wire N__3525;
    wire N__3522;
    wire N__3519;
    wire N__3514;
    wire N__3513;
    wire N__3512;
    wire N__3509;
    wire N__3506;
    wire N__3503;
    wire N__3500;
    wire N__3497;
    wire N__3494;
    wire N__3487;
    wire N__3484;
    wire N__3481;
    wire N__3478;
    wire N__3475;
    wire N__3472;
    wire N__3469;
    wire N__3466;
    wire N__3463;
    wire N__3460;
    wire N__3459;
    wire N__3458;
    wire N__3457;
    wire N__3452;
    wire N__3449;
    wire N__3446;
    wire N__3445;
    wire N__3440;
    wire N__3437;
    wire N__3434;
    wire N__3431;
    wire N__3428;
    wire N__3425;
    wire N__3422;
    wire N__3419;
    wire N__3416;
    wire N__3409;
    wire N__3406;
    wire N__3403;
    wire N__3400;
    wire N__3399;
    wire N__3394;
    wire N__3391;
    wire N__3390;
    wire N__3387;
    wire N__3386;
    wire N__3383;
    wire N__3380;
    wire N__3377;
    wire N__3374;
    wire N__3371;
    wire N__3368;
    wire N__3365;
    wire N__3360;
    wire N__3357;
    wire N__3352;
    wire N__3351;
    wire N__3346;
    wire N__3345;
    wire N__3342;
    wire N__3339;
    wire N__3334;
    wire N__3331;
    wire N__3328;
    wire N__3325;
    wire N__3322;
    wire N__3321;
    wire N__3320;
    wire N__3317;
    wire N__3314;
    wire N__3311;
    wire N__3306;
    wire N__3303;
    wire N__3300;
    wire N__3297;
    wire N__3294;
    wire N__3291;
    wire N__3288;
    wire N__3285;
    wire N__3280;
    wire N__3279;
    wire N__3278;
    wire N__3275;
    wire N__3270;
    wire N__3267;
    wire N__3264;
    wire N__3261;
    wire N__3258;
    wire N__3255;
    wire N__3252;
    wire N__3249;
    wire N__3244;
    wire N__3241;
    wire N__3238;
    wire N__3235;
    wire N__3232;
    wire N__3229;
    wire N__3226;
    wire N__3223;
    wire N__3220;
    wire N__3217;
    wire N__3214;
    wire N__3211;
    wire N__3208;
    wire N__3205;
    wire N__3202;
    wire N__3199;
    wire N__3196;
    wire N__3193;
    wire N__3190;
    wire N__3187;
    wire N__3186;
    wire N__3183;
    wire N__3180;
    wire N__3177;
    wire N__3174;
    wire N__3169;
    wire N__3166;
    wire N__3165;
    wire N__3164;
    wire N__3161;
    wire N__3156;
    wire N__3153;
    wire N__3150;
    wire N__3149;
    wire N__3146;
    wire N__3143;
    wire N__3140;
    wire N__3137;
    wire N__3132;
    wire N__3127;
    wire N__3124;
    wire N__3121;
    wire N__3120;
    wire N__3115;
    wire N__3114;
    wire N__3113;
    wire N__3110;
    wire N__3107;
    wire N__3104;
    wire N__3099;
    wire N__3096;
    wire N__3093;
    wire N__3090;
    wire N__3087;
    wire N__3084;
    wire N__3081;
    wire N__3076;
    wire N__3075;
    wire N__3074;
    wire N__3071;
    wire N__3068;
    wire N__3061;
    wire N__3058;
    wire N__3055;
    wire N__3052;
    wire N__3049;
    wire N__3046;
    wire N__3043;
    wire N__3040;
    wire N__3039;
    wire N__3038;
    wire N__3031;
    wire N__3028;
    wire N__3025;
    wire N__3022;
    wire N__3019;
    wire N__3016;
    wire N__3013;
    wire N__3010;
    wire N__3007;
    wire N__3004;
    wire N__3001;
    wire N__2998;
    wire N__2995;
    wire N__2992;
    wire N__2989;
    wire N__2986;
    wire N__2983;
    wire N__2982;
    wire N__2981;
    wire N__2978;
    wire N__2973;
    wire N__2970;
    wire N__2967;
    wire N__2964;
    wire N__2961;
    wire N__2958;
    wire N__2955;
    wire N__2952;
    wire N__2949;
    wire N__2944;
    wire N__2941;
    wire N__2938;
    wire N__2935;
    wire N__2932;
    wire N__2929;
    wire N__2928;
    wire N__2927;
    wire N__2924;
    wire N__2921;
    wire N__2918;
    wire N__2915;
    wire N__2910;
    wire N__2905;
    wire N__2902;
    wire N__2899;
    wire N__2898;
    wire N__2897;
    wire N__2896;
    wire N__2895;
    wire N__2894;
    wire N__2893;
    wire N__2892;
    wire N__2891;
    wire N__2890;
    wire N__2889;
    wire N__2888;
    wire N__2887;
    wire N__2886;
    wire N__2857;
    wire CLK80_OUT;
    wire GNDG0;
    wire VCCG0;
    wire A_c_28;
    wire \U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_7_cascade_ ;
    wire A_c_29;
    wire \U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_8 ;
    wire \U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_9_cascade_ ;
    wire \U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_10 ;
    wire N_31_i;
    wire A_c_31;
    wire TT_c_1;
    wire A_c_30;
    wire A_c_27;
    wire A_c_26;
    wire A_c_24;
    wire A_c_25;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_7 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_8_cascade_ ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_10 ;
    wire N_69_i;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_13 ;
    wire N_101_cascade_;
    wire N_105;
    wire A_c_16;
    wire A_c_17;
    wire N_74_1_cascade_;
    wire N_33_cascade_;
    wire N_99;
    wire U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_a2_5;
    wire N_99_cascade_;
    wire U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_a2_4;
    wire A_c_18;
    wire N_74_1;
    wire N_101;
    wire TT_c_0;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_9 ;
    wire A_c_19;
    wire \U409_ADDRESS_DECODE.HIROMZ0Z_1_cascade_ ;
    wire \U409_TRANSFER_ACK.N_94 ;
    wire \U409_DATA_BUFFERS.un1_BUFENn_iZ0Z_0 ;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_1 ;
    wire A_c_20;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4_cascade_ ;
    wire CIA_SPACE_cascade_;
    wire \U409_ADDRESS_DECODE.N_69 ;
    wire PORTSIZE_0_i;
    wire \U409_ADDRESS_DECODE.un5_RAMSPACEn_cascade_ ;
    wire A_c_21;
    wire A_c_23;
    wire A_c_22;
    wire TM_c_0;
    wire U409_ADDRESS_DECODE_HIROM;
    wire U409_ADDRESS_DECODE_LOWROM_cascade_;
    wire TM_c_1;
    wire N_107;
    wire N_33;
    wire N_68_i;
    wire \U409_TRANSFER_ACK.N_71 ;
    wire TACKn_in;
    wire N_67_i;
    wire N_100;
    wire OVL_c;
    wire N_67;
    wire \INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ;
    wire \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ;
    wire \U409_TRANSFER_ACK.N_106 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER15Z0Z_1 ;
    wire U409_ADDRESS_DECODE_Z2_SPACE;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER20_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_cascade_ ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER20 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ;
    wire ROMENn_c;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ;
    wire \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_ ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.CIA_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ;
    wire \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ;
    wire TACK_OUTn;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_0C_net ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER6 ;
    wire \INVU409_TRANSFER_ACK.TACK_EN_iC_net ;
    wire \U409_TRANSFER_ACK.TACK_OUTn_0_sqmuxa_0_en ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a4_3_cascade_ ;
    wire \U409_TRANSFER_ACK.N_70_cascade_ ;
    wire \U409_TRANSFER_ACK.N_55 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out ;
    wire CONSTANT_ONE_NET;
    wire \U409_TRANSFER_ACK.CO1 ;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0 ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_EN_e_1 ;
    wire \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0 ;
    wire \U409_TRANSFER_ACK.N_17_mux ;
    wire \U409_TRANSFER_ACK.N_3_0 ;
    wire \U409_TRANSFER_ACK.N_3_0_cascade_ ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ;
    wire \U409_TRANSFER_ACK.N_6_0_cascade_ ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_1C_net ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ;
    wire TSn_c;
    wire CLK40_IN_c;
    wire \U409_TRANSFER_ACK.N_70 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ;
    wire A_c_13;
    wire U409_ADDRESS_DECODE_un1_CIACS1n_i;
    wire A_c_12;
    wire U409_ADDRESS_DECODE_un1_CIACS0n_i;
    wire CIA_ENABLE;
    wire RESETn_c;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_0 ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.LASTCLK_0C_net ;
    wire RESETn_c_i;
    wire \U409_TICK.TICK603_8_cascade_ ;
    wire \U409_TICK.TICK603_14_cascade_ ;
    wire \U409_TICK.TICK603_11 ;
    wire \U409_TICK.TICK603_10_cascade_ ;
    wire \U409_TICK.TICK503_10_cascade_ ;
    wire TICK50_c;
    wire \U409_TICK.TICK503_9_cascade_ ;
    wire \U409_TICK.TICK503_11 ;
    wire \U409_TICK.TICK503_8_cascade_ ;
    wire \U409_TICK.TICK503_14_cascade_ ;
    wire \U409_TICK.TICK503_14 ;
    wire \U409_TICK.TICK503_10 ;
    wire \U409_TICK.TICK503_9 ;
    wire TICK60_c;
    wire \U409_TICK.TICK603_9_cascade_ ;
    wire \U409_TICK.TICK603_9 ;
    wire \U409_TICK.TICK603_14 ;
    wire \U409_TICK.TICK603_10 ;
    wire \U409_TICK.COUNTER60Z0Z_1 ;
    wire \U409_TICK.COUNTER60Z0Z_0 ;
    wire bfn_14_8_0_;
    wire \U409_TICK.COUNTER60Z0Z_2 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_1 ;
    wire \U409_TICK.COUNTER60Z0Z_3 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_2 ;
    wire \U409_TICK.COUNTER60Z0Z_4 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_4 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_3 ;
    wire \U409_TICK.COUNTER60Z0Z_5 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_4 ;
    wire \U409_TICK.COUNTER60Z0Z_6 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_6 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_5 ;
    wire \U409_TICK.COUNTER60Z0Z_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_6 ;
    wire \U409_TICK.COUNTER60Z0Z_8 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_8 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_8 ;
    wire \U409_TICK.COUNTER60Z0Z_9 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_9 ;
    wire bfn_14_9_0_;
    wire \U409_TICK.COUNTER60Z0Z_10 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_9 ;
    wire \U409_TICK.COUNTER60Z0Z_11 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_10 ;
    wire \U409_TICK.COUNTER60Z0Z_12 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_11 ;
    wire \U409_TICK.COUNTER60Z0Z_13 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_12 ;
    wire \U409_TICK.COUNTER60Z0Z_14 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_13 ;
    wire \U409_TICK.COUNTER60Z0Z_15 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_15 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_15 ;
    wire \U409_TICK.COUNTER60Z0Z_16 ;
    wire \U409_TICK.COUNTER50Z0Z_1 ;
    wire \U409_TICK.COUNTER50Z0Z_0 ;
    wire bfn_15_3_0_;
    wire \U409_TICK.COUNTER50Z0Z_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_1 ;
    wire \U409_TICK.COUNTER50Z0Z_3 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_2 ;
    wire \U409_TICK.COUNTER50Z0Z_4 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_3 ;
    wire \U409_TICK.COUNTER50Z0Z_5 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_5 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_4 ;
    wire \U409_TICK.COUNTER50Z0Z_6 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_6 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_5 ;
    wire \U409_TICK.COUNTER50Z0Z_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_6 ;
    wire \U409_TICK.COUNTER50Z0Z_8 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_8 ;
    wire \U409_TICK.COUNTER50Z0Z_9 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_9 ;
    wire bfn_15_4_0_;
    wire \U409_TICK.COUNTER50Z0Z_10 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_9 ;
    wire \U409_TICK.COUNTER50Z0Z_11 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_11 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_10 ;
    wire \U409_TICK.COUNTER50Z0Z_12 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_11 ;
    wire \U409_TICK.COUNTER50Z0Z_13 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_13 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_12 ;
    wire \U409_TICK.COUNTER50Z0Z_14 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_13 ;
    wire \U409_TICK.COUNTER50Z0Z_15 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_15 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_15 ;
    wire \U409_TICK.COUNTER50Z0Z_16 ;
    wire CLK6_c_g;
    wire bfn_15_6_0_;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_1 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_3 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_5 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_6 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_3 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_7 ;
    wire \U409_CIA.un1_CIA_CLK_COUNT_2_0_a4_1_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_6 ;
    wire \U409_CIA.CLK_CIA_RNOZ0Z_1_cascade_ ;
    wire CLK_CIA_c;
    wire \U409_CIA.un1_CIA_CLK_COUNT_3_0_a4_0_cascade_ ;
    wire CIA_SPACE;
    wire \U409_CIA.VMA_RNOZ0Z_0_cascade_ ;
    wire \U409_CIA.VMAZ0 ;
    wire \U409_CIA.CIA_CLK_COUNT11_0_a4_2_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNT11 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_2 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_5 ;
    wire \U409_CIA.CLK_CIA6_1 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_4 ;
    wire \U409_CIA.CLK_CIA6_1_cascade_ ;
    wire \U409_CIA.N_104 ;
    wire \U409_CIA.CLK_CIA6 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_1 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_0 ;
    wire CLK28_IN_c_g;
    wire TACK_EN_i;
    wire N_465_i;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="SIMPLE";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0001111;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE pll (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__4882),
            .RESETB(N__4759),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(CLK80_OUT));
    PRE_IO_GBUF CLK28_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__7446),
            .GLOBALBUFFEROUTPUT(CLK28_IN_c_g));
    IO_PAD CLK28_IN_ibuf_gb_io_iopad (
            .OE(N__7448),
            .DIN(N__7447),
            .DOUT(N__7446),
            .PACKAGEPIN(CLK28_IN));
    defparam CLK28_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK28_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK28_IN_ibuf_gb_io_preio (
            .PADOEN(N__7448),
            .PADOUT(N__7447),
            .PADIN(N__7446),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK6_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__7436),
            .GLOBALBUFFEROUTPUT(CLK6_c_g));
    IO_PAD CLK6_ibuf_gb_io_iopad (
            .OE(N__7438),
            .DIN(N__7437),
            .DOUT(N__7436),
            .PACKAGEPIN(CLK6));
    defparam CLK6_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK6_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK6_ibuf_gb_io_preio (
            .PADOEN(N__7438),
            .PADOUT(N__7437),
            .PADIN(N__7436),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_0_iopad (
            .OE(N__7427),
            .DIN(N__7426),
            .DOUT(N__7425),
            .PACKAGEPIN(TT[0]));
    defparam TT_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_0_preio (
            .PADOEN(N__7427),
            .PADOUT(N__7426),
            .PADIN(N__7425),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_6_iopad (
            .OE(N__7418),
            .DIN(N__7417),
            .DOUT(N__7416),
            .PACKAGEPIN(D[6]));
    defparam D_obuft_6_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_6_preio (
            .PADOEN(N__7418),
            .PADOUT(N__7417),
            .PADIN(N__7416),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RTC_ENn_obuf_iopad (
            .OE(N__7409),
            .DIN(N__7408),
            .DOUT(N__7407),
            .PACKAGEPIN(RTC_ENn));
    defparam RTC_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RTC_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RTC_ENn_obuf_preio (
            .PADOEN(N__7409),
            .PADOUT(N__7408),
            .PADIN(N__7407),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3226),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_24_iopad (
            .OE(N__7400),
            .DIN(N__7399),
            .DOUT(N__7398),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__7400),
            .PADOUT(N__7399),
            .PADIN(N__7398),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_5_iopad (
            .OE(N__7391),
            .DIN(N__7390),
            .DOUT(N__7389),
            .PACKAGEPIN(D[5]));
    defparam D_obuft_5_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_5_preio (
            .PADOEN(N__7391),
            .PADOUT(N__7390),
            .PADIN(N__7389),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TM_ibuf_1_iopad (
            .OE(N__7382),
            .DIN(N__7381),
            .DOUT(N__7380),
            .PACKAGEPIN(TM[1]));
    defparam TM_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TM_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TM_ibuf_1_preio (
            .PADOEN(N__7382),
            .PADOUT(N__7381),
            .PADIN(N__7380),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TM_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__7373),
            .DIN(N__7372),
            .DOUT(N__7371),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__7373),
            .PADOUT(N__7372),
            .PADIN(N__7371),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_CIA_obuf_iopad (
            .OE(N__7364),
            .DIN(N__7363),
            .DOUT(N__7362),
            .PACKAGEPIN(CLK_CIA));
    defparam CLK_CIA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_CIA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_CIA_obuf_preio (
            .PADOEN(N__7364),
            .PADOUT(N__7363),
            .PADIN(N__7362),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6856),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_21_iopad (
            .OE(N__7355),
            .DIN(N__7354),
            .DOUT(N__7353),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__7355),
            .PADOUT(N__7354),
            .PADIN(N__7353),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_obuf_iopad (
            .OE(N__7346),
            .DIN(N__7345),
            .DOUT(N__7344),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMSPACEn_obuf_preio (
            .PADOEN(N__7346),
            .PADOUT(N__7345),
            .PADIN(N__7344),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4228),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__7337),
            .DIN(N__7336),
            .DOUT(N__7335),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__7337),
            .PADOUT(N__7336),
            .PADIN(N__7335),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6910),
            .DIN0(TACKn_in),
            .DOUT0(N__4519),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__7328),
            .DIN(N__7327),
            .DOUT(N__7326),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__7328),
            .PADOUT(N__7327),
            .PADIN(N__7326),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ROMENn_obuf_iopad (
            .OE(N__7319),
            .DIN(N__7318),
            .DOUT(N__7317),
            .PACKAGEPIN(ROMENn));
    defparam ROMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ROMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ROMENn_obuf_preio (
            .PADOEN(N__7319),
            .PADOUT(N__7318),
            .PADIN(N__7317),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4348),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_0_iopad (
            .OE(N__7310),
            .DIN(N__7309),
            .DOUT(N__7308),
            .PACKAGEPIN(D[0]));
    defparam D_obuft_0_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_0_preio (
            .PADOEN(N__7310),
            .PADOUT(N__7309),
            .PADIN(N__7308),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_1_iopad (
            .OE(N__7301),
            .DIN(N__7300),
            .DOUT(N__7299),
            .PACKAGEPIN(TT[1]));
    defparam TT_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_1_preio (
            .PADOEN(N__7301),
            .PADOUT(N__7300),
            .PADIN(N__7299),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__7292),
            .DIN(N__7291),
            .DOUT(N__7290),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__7292),
            .PADOUT(N__7291),
            .PADIN(N__7290),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__7283),
            .DIN(N__7282),
            .DOUT(N__7281),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__7283),
            .PADOUT(N__7282),
            .PADIN(N__7281),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3004),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PORTSIZE_obuf_iopad (
            .OE(N__7274),
            .DIN(N__7273),
            .DOUT(N__7272),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PORTSIZE_obuf_preio (
            .PADOEN(N__7274),
            .PADOUT(N__7273),
            .PADIN(N__7272),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3949),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_7_iopad (
            .OE(N__7265),
            .DIN(N__7264),
            .DOUT(N__7263),
            .PACKAGEPIN(D[7]));
    defparam D_obuft_7_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_7_preio (
            .PADOEN(N__7265),
            .PADOUT(N__7264),
            .PADIN(N__7263),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__7256),
            .DIN(N__7255),
            .DOUT(N__7254),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__7256),
            .PADOUT(N__7255),
            .PADIN(N__7254),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_29_iopad (
            .OE(N__7247),
            .DIN(N__7246),
            .DOUT(N__7245),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__7247),
            .PADOUT(N__7246),
            .PADIN(N__7245),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_22_iopad (
            .OE(N__7238),
            .DIN(N__7237),
            .DOUT(N__7236),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__7238),
            .PADOUT(N__7237),
            .PADIN(N__7236),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_27_iopad (
            .OE(N__7229),
            .DIN(N__7228),
            .DOUT(N__7227),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__7229),
            .PADOUT(N__7228),
            .PADIN(N__7227),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__7220),
            .DIN(N__7219),
            .DOUT(N__7218),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__7220),
            .PADOUT(N__7219),
            .PADIN(N__7218),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_2_iopad (
            .OE(N__7211),
            .DIN(N__7210),
            .DOUT(N__7209),
            .PACKAGEPIN(D[2]));
    defparam D_obuft_2_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_2_preio (
            .PADOEN(N__7211),
            .PADOUT(N__7210),
            .PADIN(N__7209),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__7202),
            .DIN(N__7201),
            .DOUT(N__7200),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__7202),
            .PADOUT(N__7201),
            .PADIN(N__7200),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TM_ibuf_0_iopad (
            .OE(N__7193),
            .DIN(N__7192),
            .DOUT(N__7191),
            .PACKAGEPIN(TM[0]));
    defparam TM_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TM_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TM_ibuf_0_preio (
            .PADOEN(N__7193),
            .PADOUT(N__7192),
            .PADIN(N__7191),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TM_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__7184),
            .DIN(N__7183),
            .DOUT(N__7182),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__7184),
            .PADOUT(N__7183),
            .PADIN(N__7182),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__7175),
            .DIN(N__7174),
            .DOUT(N__7173),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__7175),
            .PADOUT(N__7174),
            .PADIN(N__7173),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_25_iopad (
            .OE(N__7166),
            .DIN(N__7165),
            .DOUT(N__7164),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__7166),
            .PADOUT(N__7165),
            .PADIN(N__7164),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_1_iopad (
            .OE(N__7157),
            .DIN(N__7156),
            .DOUT(N__7155),
            .PACKAGEPIN(D[1]));
    defparam D_obuft_1_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_1_preio (
            .PADOEN(N__7157),
            .PADOUT(N__7156),
            .PADIN(N__7155),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS0n_obuf_iopad (
            .OE(N__7148),
            .DIN(N__7147),
            .DOUT(N__7146),
            .PACKAGEPIN(CIACS0n));
    defparam CIACS0n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS0n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS0n_obuf_preio (
            .PADOEN(N__7148),
            .PADOUT(N__7147),
            .PADIN(N__7146),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5371),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_4_iopad (
            .OE(N__7139),
            .DIN(N__7138),
            .DOUT(N__7137),
            .PACKAGEPIN(D[4]));
    defparam D_obuft_4_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_4_preio (
            .PADOEN(N__7139),
            .PADOUT(N__7138),
            .PADIN(N__7137),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK50_obuf_iopad (
            .OE(N__7130),
            .DIN(N__7129),
            .DOUT(N__7128),
            .PACKAGEPIN(TICK50));
    defparam TICK50_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK50_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK50_obuf_preio (
            .PADOEN(N__7130),
            .PADOUT(N__7129),
            .PADIN(N__7128),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5677),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__7121),
            .DIN(N__7120),
            .DOUT(N__7119),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__7121),
            .PADOUT(N__7120),
            .PADIN(N__7119),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_28_iopad (
            .OE(N__7112),
            .DIN(N__7111),
            .DOUT(N__7110),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__7112),
            .PADOUT(N__7111),
            .PADIN(N__7110),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_30_iopad (
            .OE(N__7103),
            .DIN(N__7102),
            .DOUT(N__7101),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__7103),
            .PADOUT(N__7102),
            .PADIN(N__7101),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD OVL_ibuf_iopad (
            .OE(N__7094),
            .DIN(N__7093),
            .DOUT(N__7092),
            .PACKAGEPIN(OVL));
    defparam OVL_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam OVL_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO OVL_ibuf_preio (
            .PADOEN(N__7094),
            .PADOUT(N__7093),
            .PADIN(N__7092),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(OVL_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__7085),
            .DIN(N__7084),
            .DOUT(N__7083),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__7085),
            .PADOUT(N__7084),
            .PADIN(N__7083),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK60_obuf_iopad (
            .OE(N__7076),
            .DIN(N__7075),
            .DOUT(N__7074),
            .PACKAGEPIN(TICK60));
    defparam TICK60_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK60_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK60_obuf_preio (
            .PADOEN(N__7076),
            .PADOUT(N__7075),
            .PADIN(N__7074),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5806),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_26_iopad (
            .OE(N__7067),
            .DIN(N__7066),
            .DOUT(N__7065),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__7067),
            .PADOUT(N__7066),
            .PADIN(N__7065),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_3_iopad (
            .OE(N__7058),
            .DIN(N__7057),
            .DOUT(N__7056),
            .PACKAGEPIN(D[3]));
    defparam D_obuft_3_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_3_preio (
            .PADOEN(N__7058),
            .PADOUT(N__7057),
            .PADIN(N__7056),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_23_iopad (
            .OE(N__7049),
            .DIN(N__7048),
            .DOUT(N__7047),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__7049),
            .PADOUT(N__7048),
            .PADIN(N__7047),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_31_iopad (
            .OE(N__7040),
            .DIN(N__7039),
            .DOUT(N__7038),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__7040),
            .PADOUT(N__7039),
            .PADIN(N__7038),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS1n_obuf_iopad (
            .OE(N__7031),
            .DIN(N__7030),
            .DOUT(N__7029),
            .PACKAGEPIN(CIACS1n));
    defparam CIACS1n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS1n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS1n_obuf_preio (
            .PADOEN(N__7031),
            .PADOUT(N__7030),
            .PADIN(N__7029),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5410),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_obuf_iopad (
            .OE(N__7022),
            .DIN(N__7021),
            .DOUT(N__7020),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGSPACEn_obuf_preio (
            .PADOEN(N__7022),
            .PADOUT(N__7021),
            .PADIN(N__7020),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3673),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__1632 (
            .O(N__7003),
            .I(N__6998));
    InMux I__1631 (
            .O(N__7002),
            .I(N__6989));
    InMux I__1630 (
            .O(N__7001),
            .I(N__6989));
    InMux I__1629 (
            .O(N__6998),
            .I(N__6986));
    InMux I__1628 (
            .O(N__6997),
            .I(N__6977));
    InMux I__1627 (
            .O(N__6996),
            .I(N__6977));
    InMux I__1626 (
            .O(N__6995),
            .I(N__6977));
    InMux I__1625 (
            .O(N__6994),
            .I(N__6977));
    LocalMux I__1624 (
            .O(N__6989),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__1623 (
            .O(N__6986),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__1622 (
            .O(N__6977),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    CascadeMux I__1621 (
            .O(N__6970),
            .I(N__6965));
    InMux I__1620 (
            .O(N__6969),
            .I(N__6959));
    InMux I__1619 (
            .O(N__6968),
            .I(N__6954));
    InMux I__1618 (
            .O(N__6965),
            .I(N__6954));
    InMux I__1617 (
            .O(N__6964),
            .I(N__6947));
    InMux I__1616 (
            .O(N__6963),
            .I(N__6947));
    InMux I__1615 (
            .O(N__6962),
            .I(N__6947));
    LocalMux I__1614 (
            .O(N__6959),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1613 (
            .O(N__6954),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1612 (
            .O(N__6947),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    ClkMux I__1611 (
            .O(N__6940),
            .I(N__6931));
    ClkMux I__1610 (
            .O(N__6939),
            .I(N__6931));
    ClkMux I__1609 (
            .O(N__6938),
            .I(N__6931));
    GlobalMux I__1608 (
            .O(N__6931),
            .I(N__6928));
    gio2CtrlBuf I__1607 (
            .O(N__6928),
            .I(CLK28_IN_c_g));
    InMux I__1606 (
            .O(N__6925),
            .I(N__6922));
    LocalMux I__1605 (
            .O(N__6922),
            .I(N__6919));
    Span4Mux_v I__1604 (
            .O(N__6919),
            .I(N__6916));
    Span4Mux_h I__1603 (
            .O(N__6916),
            .I(N__6913));
    Odrv4 I__1602 (
            .O(N__6913),
            .I(TACK_EN_i));
    IoInMux I__1601 (
            .O(N__6910),
            .I(N__6907));
    LocalMux I__1600 (
            .O(N__6907),
            .I(N__6904));
    Span4Mux_s2_v I__1599 (
            .O(N__6904),
            .I(N__6901));
    Sp12to4 I__1598 (
            .O(N__6901),
            .I(N__6898));
    Span12Mux_h I__1597 (
            .O(N__6898),
            .I(N__6895));
    Odrv12 I__1596 (
            .O(N__6895),
            .I(N_465_i));
    InMux I__1595 (
            .O(N__6892),
            .I(N__6887));
    InMux I__1594 (
            .O(N__6891),
            .I(N__6882));
    InMux I__1593 (
            .O(N__6890),
            .I(N__6882));
    LocalMux I__1592 (
            .O(N__6887),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    LocalMux I__1591 (
            .O(N__6882),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    CascadeMux I__1590 (
            .O(N__6877),
            .I(\U409_CIA.un1_CIA_CLK_COUNT_2_0_a4_1_cascade_ ));
    InMux I__1589 (
            .O(N__6874),
            .I(N__6869));
    InMux I__1588 (
            .O(N__6873),
            .I(N__6864));
    InMux I__1587 (
            .O(N__6872),
            .I(N__6864));
    LocalMux I__1586 (
            .O(N__6869),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__1585 (
            .O(N__6864),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    CascadeMux I__1584 (
            .O(N__6859),
            .I(\U409_CIA.CLK_CIA_RNOZ0Z_1_cascade_ ));
    IoInMux I__1583 (
            .O(N__6856),
            .I(N__6853));
    LocalMux I__1582 (
            .O(N__6853),
            .I(N__6850));
    IoSpan4Mux I__1581 (
            .O(N__6850),
            .I(N__6847));
    Span4Mux_s1_v I__1580 (
            .O(N__6847),
            .I(N__6844));
    Sp12to4 I__1579 (
            .O(N__6844),
            .I(N__6840));
    InMux I__1578 (
            .O(N__6843),
            .I(N__6837));
    Span12Mux_s9_v I__1577 (
            .O(N__6840),
            .I(N__6833));
    LocalMux I__1576 (
            .O(N__6837),
            .I(N__6830));
    InMux I__1575 (
            .O(N__6836),
            .I(N__6827));
    Odrv12 I__1574 (
            .O(N__6833),
            .I(CLK_CIA_c));
    Odrv4 I__1573 (
            .O(N__6830),
            .I(CLK_CIA_c));
    LocalMux I__1572 (
            .O(N__6827),
            .I(CLK_CIA_c));
    CascadeMux I__1571 (
            .O(N__6820),
            .I(\U409_CIA.un1_CIA_CLK_COUNT_3_0_a4_0_cascade_ ));
    InMux I__1570 (
            .O(N__6817),
            .I(N__6814));
    LocalMux I__1569 (
            .O(N__6814),
            .I(N__6811));
    Span4Mux_v I__1568 (
            .O(N__6811),
            .I(N__6808));
    Sp12to4 I__1567 (
            .O(N__6808),
            .I(N__6805));
    Span12Mux_h I__1566 (
            .O(N__6805),
            .I(N__6802));
    Odrv12 I__1565 (
            .O(N__6802),
            .I(CIA_SPACE));
    CascadeMux I__1564 (
            .O(N__6799),
            .I(\U409_CIA.VMA_RNOZ0Z_0_cascade_ ));
    InMux I__1563 (
            .O(N__6796),
            .I(N__6792));
    InMux I__1562 (
            .O(N__6795),
            .I(N__6789));
    LocalMux I__1561 (
            .O(N__6792),
            .I(N__6786));
    LocalMux I__1560 (
            .O(N__6789),
            .I(N__6783));
    Span4Mux_v I__1559 (
            .O(N__6786),
            .I(N__6777));
    Span4Mux_v I__1558 (
            .O(N__6783),
            .I(N__6777));
    InMux I__1557 (
            .O(N__6782),
            .I(N__6774));
    Odrv4 I__1556 (
            .O(N__6777),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__1555 (
            .O(N__6774),
            .I(\U409_CIA.VMAZ0 ));
    CascadeMux I__1554 (
            .O(N__6769),
            .I(\U409_CIA.CIA_CLK_COUNT11_0_a4_2_cascade_ ));
    InMux I__1553 (
            .O(N__6766),
            .I(N__6760));
    InMux I__1552 (
            .O(N__6765),
            .I(N__6760));
    LocalMux I__1551 (
            .O(N__6760),
            .I(\U409_CIA.CIA_CLK_COUNT11 ));
    InMux I__1550 (
            .O(N__6757),
            .I(N__6754));
    LocalMux I__1549 (
            .O(N__6754),
            .I(N__6748));
    InMux I__1548 (
            .O(N__6753),
            .I(N__6745));
    InMux I__1547 (
            .O(N__6752),
            .I(N__6742));
    InMux I__1546 (
            .O(N__6751),
            .I(N__6739));
    Odrv4 I__1545 (
            .O(N__6748),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__1544 (
            .O(N__6745),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__1543 (
            .O(N__6742),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__1542 (
            .O(N__6739),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    InMux I__1541 (
            .O(N__6730),
            .I(N__6724));
    InMux I__1540 (
            .O(N__6729),
            .I(N__6721));
    InMux I__1539 (
            .O(N__6728),
            .I(N__6716));
    InMux I__1538 (
            .O(N__6727),
            .I(N__6716));
    LocalMux I__1537 (
            .O(N__6724),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__1536 (
            .O(N__6721),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__1535 (
            .O(N__6716),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    InMux I__1534 (
            .O(N__6709),
            .I(N__6706));
    LocalMux I__1533 (
            .O(N__6706),
            .I(\U409_CIA.CLK_CIA6_1 ));
    InMux I__1532 (
            .O(N__6703),
            .I(N__6696));
    InMux I__1531 (
            .O(N__6702),
            .I(N__6693));
    InMux I__1530 (
            .O(N__6701),
            .I(N__6686));
    InMux I__1529 (
            .O(N__6700),
            .I(N__6686));
    InMux I__1528 (
            .O(N__6699),
            .I(N__6686));
    LocalMux I__1527 (
            .O(N__6696),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__1526 (
            .O(N__6693),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__1525 (
            .O(N__6686),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    CascadeMux I__1524 (
            .O(N__6679),
            .I(\U409_CIA.CLK_CIA6_1_cascade_ ));
    InMux I__1523 (
            .O(N__6676),
            .I(N__6671));
    InMux I__1522 (
            .O(N__6675),
            .I(N__6666));
    InMux I__1521 (
            .O(N__6674),
            .I(N__6666));
    LocalMux I__1520 (
            .O(N__6671),
            .I(\U409_CIA.N_104 ));
    LocalMux I__1519 (
            .O(N__6666),
            .I(\U409_CIA.N_104 ));
    InMux I__1518 (
            .O(N__6661),
            .I(N__6658));
    LocalMux I__1517 (
            .O(N__6658),
            .I(\U409_CIA.CLK_CIA6 ));
    InMux I__1516 (
            .O(N__6655),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ));
    InMux I__1515 (
            .O(N__6652),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ));
    InMux I__1514 (
            .O(N__6649),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ));
    InMux I__1513 (
            .O(N__6646),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ));
    InMux I__1512 (
            .O(N__6643),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ));
    InMux I__1511 (
            .O(N__6640),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ));
    CascadeMux I__1510 (
            .O(N__6637),
            .I(N__6633));
    InMux I__1509 (
            .O(N__6636),
            .I(N__6629));
    InMux I__1508 (
            .O(N__6633),
            .I(N__6624));
    InMux I__1507 (
            .O(N__6632),
            .I(N__6624));
    LocalMux I__1506 (
            .O(N__6629),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__1505 (
            .O(N__6624),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    InMux I__1504 (
            .O(N__6619),
            .I(N__6615));
    InMux I__1503 (
            .O(N__6618),
            .I(N__6612));
    LocalMux I__1502 (
            .O(N__6615),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    LocalMux I__1501 (
            .O(N__6612),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    InMux I__1500 (
            .O(N__6607),
            .I(N__6604));
    LocalMux I__1499 (
            .O(N__6604),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ));
    InMux I__1498 (
            .O(N__6601),
            .I(bfn_15_4_0_));
    InMux I__1497 (
            .O(N__6598),
            .I(N__6594));
    InMux I__1496 (
            .O(N__6597),
            .I(N__6591));
    LocalMux I__1495 (
            .O(N__6594),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    LocalMux I__1494 (
            .O(N__6591),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    InMux I__1493 (
            .O(N__6586),
            .I(\U409_TICK.un2_COUNTER50_1_cry_9 ));
    InMux I__1492 (
            .O(N__6583),
            .I(N__6579));
    InMux I__1491 (
            .O(N__6582),
            .I(N__6576));
    LocalMux I__1490 (
            .O(N__6579),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    LocalMux I__1489 (
            .O(N__6576),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    InMux I__1488 (
            .O(N__6571),
            .I(N__6568));
    LocalMux I__1487 (
            .O(N__6568),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ));
    InMux I__1486 (
            .O(N__6565),
            .I(\U409_TICK.un2_COUNTER50_1_cry_10 ));
    InMux I__1485 (
            .O(N__6562),
            .I(N__6558));
    InMux I__1484 (
            .O(N__6561),
            .I(N__6555));
    LocalMux I__1483 (
            .O(N__6558),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    LocalMux I__1482 (
            .O(N__6555),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    InMux I__1481 (
            .O(N__6550),
            .I(\U409_TICK.un2_COUNTER50_1_cry_11 ));
    InMux I__1480 (
            .O(N__6547),
            .I(N__6543));
    InMux I__1479 (
            .O(N__6546),
            .I(N__6540));
    LocalMux I__1478 (
            .O(N__6543),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    LocalMux I__1477 (
            .O(N__6540),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    InMux I__1476 (
            .O(N__6535),
            .I(N__6532));
    LocalMux I__1475 (
            .O(N__6532),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ));
    InMux I__1474 (
            .O(N__6529),
            .I(\U409_TICK.un2_COUNTER50_1_cry_12 ));
    InMux I__1473 (
            .O(N__6526),
            .I(N__6522));
    InMux I__1472 (
            .O(N__6525),
            .I(N__6519));
    LocalMux I__1471 (
            .O(N__6522),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    LocalMux I__1470 (
            .O(N__6519),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    CascadeMux I__1469 (
            .O(N__6514),
            .I(N__6511));
    InMux I__1468 (
            .O(N__6511),
            .I(N__6508));
    LocalMux I__1467 (
            .O(N__6508),
            .I(N__6505));
    Odrv4 I__1466 (
            .O(N__6505),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ));
    InMux I__1465 (
            .O(N__6502),
            .I(\U409_TICK.un2_COUNTER50_1_cry_13 ));
    InMux I__1464 (
            .O(N__6499),
            .I(N__6495));
    InMux I__1463 (
            .O(N__6498),
            .I(N__6492));
    LocalMux I__1462 (
            .O(N__6495),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    LocalMux I__1461 (
            .O(N__6492),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    InMux I__1460 (
            .O(N__6487),
            .I(N__6484));
    LocalMux I__1459 (
            .O(N__6484),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ));
    InMux I__1458 (
            .O(N__6481),
            .I(\U409_TICK.un2_COUNTER50_1_cry_14 ));
    InMux I__1457 (
            .O(N__6478),
            .I(\U409_TICK.un2_COUNTER50_1_cry_15 ));
    InMux I__1456 (
            .O(N__6475),
            .I(N__6471));
    InMux I__1455 (
            .O(N__6474),
            .I(N__6468));
    LocalMux I__1454 (
            .O(N__6471),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    LocalMux I__1453 (
            .O(N__6468),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    ClkMux I__1452 (
            .O(N__6463),
            .I(N__6439));
    ClkMux I__1451 (
            .O(N__6462),
            .I(N__6439));
    ClkMux I__1450 (
            .O(N__6461),
            .I(N__6439));
    ClkMux I__1449 (
            .O(N__6460),
            .I(N__6439));
    ClkMux I__1448 (
            .O(N__6459),
            .I(N__6439));
    ClkMux I__1447 (
            .O(N__6458),
            .I(N__6439));
    ClkMux I__1446 (
            .O(N__6457),
            .I(N__6439));
    ClkMux I__1445 (
            .O(N__6456),
            .I(N__6439));
    GlobalMux I__1444 (
            .O(N__6439),
            .I(N__6436));
    gio2CtrlBuf I__1443 (
            .O(N__6436),
            .I(CLK6_c_g));
    CascadeMux I__1442 (
            .O(N__6433),
            .I(N__6429));
    InMux I__1441 (
            .O(N__6432),
            .I(N__6423));
    InMux I__1440 (
            .O(N__6429),
            .I(N__6423));
    InMux I__1439 (
            .O(N__6428),
            .I(N__6420));
    LocalMux I__1438 (
            .O(N__6423),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    LocalMux I__1437 (
            .O(N__6420),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    InMux I__1436 (
            .O(N__6415),
            .I(N__6410));
    CascadeMux I__1435 (
            .O(N__6414),
            .I(N__6406));
    InMux I__1434 (
            .O(N__6413),
            .I(N__6403));
    LocalMux I__1433 (
            .O(N__6410),
            .I(N__6400));
    InMux I__1432 (
            .O(N__6409),
            .I(N__6397));
    InMux I__1431 (
            .O(N__6406),
            .I(N__6394));
    LocalMux I__1430 (
            .O(N__6403),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    Odrv4 I__1429 (
            .O(N__6400),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__1428 (
            .O(N__6397),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__1427 (
            .O(N__6394),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    InMux I__1426 (
            .O(N__6385),
            .I(N__6381));
    InMux I__1425 (
            .O(N__6384),
            .I(N__6378));
    LocalMux I__1424 (
            .O(N__6381),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    LocalMux I__1423 (
            .O(N__6378),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    InMux I__1422 (
            .O(N__6373),
            .I(\U409_TICK.un2_COUNTER50_1_cry_1 ));
    InMux I__1421 (
            .O(N__6370),
            .I(N__6366));
    InMux I__1420 (
            .O(N__6369),
            .I(N__6363));
    LocalMux I__1419 (
            .O(N__6366),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    LocalMux I__1418 (
            .O(N__6363),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    InMux I__1417 (
            .O(N__6358),
            .I(\U409_TICK.un2_COUNTER50_1_cry_2 ));
    CascadeMux I__1416 (
            .O(N__6355),
            .I(N__6352));
    InMux I__1415 (
            .O(N__6352),
            .I(N__6348));
    InMux I__1414 (
            .O(N__6351),
            .I(N__6345));
    LocalMux I__1413 (
            .O(N__6348),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    LocalMux I__1412 (
            .O(N__6345),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    InMux I__1411 (
            .O(N__6340),
            .I(\U409_TICK.un2_COUNTER50_1_cry_3 ));
    CascadeMux I__1410 (
            .O(N__6337),
            .I(N__6333));
    InMux I__1409 (
            .O(N__6336),
            .I(N__6330));
    InMux I__1408 (
            .O(N__6333),
            .I(N__6327));
    LocalMux I__1407 (
            .O(N__6330),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    LocalMux I__1406 (
            .O(N__6327),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    CascadeMux I__1405 (
            .O(N__6322),
            .I(N__6319));
    InMux I__1404 (
            .O(N__6319),
            .I(N__6316));
    LocalMux I__1403 (
            .O(N__6316),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ));
    InMux I__1402 (
            .O(N__6313),
            .I(\U409_TICK.un2_COUNTER50_1_cry_4 ));
    CascadeMux I__1401 (
            .O(N__6310),
            .I(N__6307));
    InMux I__1400 (
            .O(N__6307),
            .I(N__6303));
    InMux I__1399 (
            .O(N__6306),
            .I(N__6300));
    LocalMux I__1398 (
            .O(N__6303),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    LocalMux I__1397 (
            .O(N__6300),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    CascadeMux I__1396 (
            .O(N__6295),
            .I(N__6292));
    InMux I__1395 (
            .O(N__6292),
            .I(N__6289));
    LocalMux I__1394 (
            .O(N__6289),
            .I(N__6286));
    Odrv4 I__1393 (
            .O(N__6286),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ));
    InMux I__1392 (
            .O(N__6283),
            .I(\U409_TICK.un2_COUNTER50_1_cry_5 ));
    InMux I__1391 (
            .O(N__6280),
            .I(N__6276));
    InMux I__1390 (
            .O(N__6279),
            .I(N__6273));
    LocalMux I__1389 (
            .O(N__6276),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    LocalMux I__1388 (
            .O(N__6273),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    InMux I__1387 (
            .O(N__6268),
            .I(\U409_TICK.un2_COUNTER50_1_cry_6 ));
    InMux I__1386 (
            .O(N__6265),
            .I(N__6261));
    InMux I__1385 (
            .O(N__6264),
            .I(N__6258));
    LocalMux I__1384 (
            .O(N__6261),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    LocalMux I__1383 (
            .O(N__6258),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    InMux I__1382 (
            .O(N__6253),
            .I(\U409_TICK.un2_COUNTER50_1_cry_7 ));
    InMux I__1381 (
            .O(N__6250),
            .I(N__6246));
    InMux I__1380 (
            .O(N__6249),
            .I(N__6243));
    LocalMux I__1379 (
            .O(N__6246),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    LocalMux I__1378 (
            .O(N__6243),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    InMux I__1377 (
            .O(N__6238),
            .I(N__6235));
    LocalMux I__1376 (
            .O(N__6235),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ));
    InMux I__1375 (
            .O(N__6232),
            .I(bfn_14_9_0_));
    InMux I__1374 (
            .O(N__6229),
            .I(N__6225));
    InMux I__1373 (
            .O(N__6228),
            .I(N__6222));
    LocalMux I__1372 (
            .O(N__6225),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    LocalMux I__1371 (
            .O(N__6222),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    InMux I__1370 (
            .O(N__6217),
            .I(\U409_TICK.un3_COUNTER60_1_cry_9 ));
    InMux I__1369 (
            .O(N__6214),
            .I(N__6210));
    InMux I__1368 (
            .O(N__6213),
            .I(N__6207));
    LocalMux I__1367 (
            .O(N__6210),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    LocalMux I__1366 (
            .O(N__6207),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    InMux I__1365 (
            .O(N__6202),
            .I(\U409_TICK.un3_COUNTER60_1_cry_10 ));
    InMux I__1364 (
            .O(N__6199),
            .I(N__6195));
    InMux I__1363 (
            .O(N__6198),
            .I(N__6192));
    LocalMux I__1362 (
            .O(N__6195),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    LocalMux I__1361 (
            .O(N__6192),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    InMux I__1360 (
            .O(N__6187),
            .I(\U409_TICK.un3_COUNTER60_1_cry_11 ));
    InMux I__1359 (
            .O(N__6184),
            .I(N__6180));
    InMux I__1358 (
            .O(N__6183),
            .I(N__6177));
    LocalMux I__1357 (
            .O(N__6180),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    LocalMux I__1356 (
            .O(N__6177),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    InMux I__1355 (
            .O(N__6172),
            .I(\U409_TICK.un3_COUNTER60_1_cry_12 ));
    InMux I__1354 (
            .O(N__6169),
            .I(N__6165));
    InMux I__1353 (
            .O(N__6168),
            .I(N__6162));
    LocalMux I__1352 (
            .O(N__6165),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    LocalMux I__1351 (
            .O(N__6162),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    InMux I__1350 (
            .O(N__6157),
            .I(N__6154));
    LocalMux I__1349 (
            .O(N__6154),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ));
    InMux I__1348 (
            .O(N__6151),
            .I(\U409_TICK.un3_COUNTER60_1_cry_13 ));
    InMux I__1347 (
            .O(N__6148),
            .I(N__6144));
    InMux I__1346 (
            .O(N__6147),
            .I(N__6141));
    LocalMux I__1345 (
            .O(N__6144),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    LocalMux I__1344 (
            .O(N__6141),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    InMux I__1343 (
            .O(N__6136),
            .I(N__6133));
    LocalMux I__1342 (
            .O(N__6133),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ));
    InMux I__1341 (
            .O(N__6130),
            .I(\U409_TICK.un3_COUNTER60_1_cry_14 ));
    InMux I__1340 (
            .O(N__6127),
            .I(\U409_TICK.un3_COUNTER60_1_cry_15 ));
    InMux I__1339 (
            .O(N__6124),
            .I(N__6120));
    InMux I__1338 (
            .O(N__6123),
            .I(N__6117));
    LocalMux I__1337 (
            .O(N__6120),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    LocalMux I__1336 (
            .O(N__6117),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    CascadeMux I__1335 (
            .O(N__6112),
            .I(N__6108));
    InMux I__1334 (
            .O(N__6111),
            .I(N__6104));
    InMux I__1333 (
            .O(N__6108),
            .I(N__6101));
    InMux I__1332 (
            .O(N__6107),
            .I(N__6098));
    LocalMux I__1331 (
            .O(N__6104),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__1330 (
            .O(N__6101),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__1329 (
            .O(N__6098),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    CascadeMux I__1328 (
            .O(N__6091),
            .I(N__6087));
    CascadeMux I__1327 (
            .O(N__6090),
            .I(N__6082));
    InMux I__1326 (
            .O(N__6087),
            .I(N__6079));
    InMux I__1325 (
            .O(N__6086),
            .I(N__6076));
    InMux I__1324 (
            .O(N__6085),
            .I(N__6073));
    InMux I__1323 (
            .O(N__6082),
            .I(N__6070));
    LocalMux I__1322 (
            .O(N__6079),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__1321 (
            .O(N__6076),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__1320 (
            .O(N__6073),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__1319 (
            .O(N__6070),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    InMux I__1318 (
            .O(N__6061),
            .I(N__6057));
    InMux I__1317 (
            .O(N__6060),
            .I(N__6054));
    LocalMux I__1316 (
            .O(N__6057),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    LocalMux I__1315 (
            .O(N__6054),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    InMux I__1314 (
            .O(N__6049),
            .I(\U409_TICK.un3_COUNTER60_1_cry_1 ));
    InMux I__1313 (
            .O(N__6046),
            .I(N__6042));
    InMux I__1312 (
            .O(N__6045),
            .I(N__6039));
    LocalMux I__1311 (
            .O(N__6042),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    LocalMux I__1310 (
            .O(N__6039),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    InMux I__1309 (
            .O(N__6034),
            .I(\U409_TICK.un3_COUNTER60_1_cry_2 ));
    InMux I__1308 (
            .O(N__6031),
            .I(N__6027));
    InMux I__1307 (
            .O(N__6030),
            .I(N__6024));
    LocalMux I__1306 (
            .O(N__6027),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    LocalMux I__1305 (
            .O(N__6024),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    InMux I__1304 (
            .O(N__6019),
            .I(N__6016));
    LocalMux I__1303 (
            .O(N__6016),
            .I(N__6013));
    Odrv4 I__1302 (
            .O(N__6013),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ));
    InMux I__1301 (
            .O(N__6010),
            .I(\U409_TICK.un3_COUNTER60_1_cry_3 ));
    InMux I__1300 (
            .O(N__6007),
            .I(N__6003));
    InMux I__1299 (
            .O(N__6006),
            .I(N__6000));
    LocalMux I__1298 (
            .O(N__6003),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    LocalMux I__1297 (
            .O(N__6000),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    InMux I__1296 (
            .O(N__5995),
            .I(\U409_TICK.un3_COUNTER60_1_cry_4 ));
    CascadeMux I__1295 (
            .O(N__5992),
            .I(N__5988));
    CascadeMux I__1294 (
            .O(N__5991),
            .I(N__5985));
    InMux I__1293 (
            .O(N__5988),
            .I(N__5982));
    InMux I__1292 (
            .O(N__5985),
            .I(N__5979));
    LocalMux I__1291 (
            .O(N__5982),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    LocalMux I__1290 (
            .O(N__5979),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    InMux I__1289 (
            .O(N__5974),
            .I(N__5971));
    LocalMux I__1288 (
            .O(N__5971),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ));
    InMux I__1287 (
            .O(N__5968),
            .I(\U409_TICK.un3_COUNTER60_1_cry_5 ));
    CascadeMux I__1286 (
            .O(N__5965),
            .I(N__5962));
    InMux I__1285 (
            .O(N__5962),
            .I(N__5959));
    LocalMux I__1284 (
            .O(N__5959),
            .I(N__5955));
    InMux I__1283 (
            .O(N__5958),
            .I(N__5952));
    Odrv4 I__1282 (
            .O(N__5955),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    LocalMux I__1281 (
            .O(N__5952),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    InMux I__1280 (
            .O(N__5947),
            .I(\U409_TICK.un3_COUNTER60_1_cry_6 ));
    InMux I__1279 (
            .O(N__5944),
            .I(N__5940));
    InMux I__1278 (
            .O(N__5943),
            .I(N__5937));
    LocalMux I__1277 (
            .O(N__5940),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    LocalMux I__1276 (
            .O(N__5937),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    InMux I__1275 (
            .O(N__5932),
            .I(N__5929));
    LocalMux I__1274 (
            .O(N__5929),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ));
    InMux I__1273 (
            .O(N__5926),
            .I(\U409_TICK.un3_COUNTER60_1_cry_7 ));
    InMux I__1272 (
            .O(N__5923),
            .I(N__5920));
    LocalMux I__1271 (
            .O(N__5920),
            .I(\U409_TICK.TICK503_11 ));
    CascadeMux I__1270 (
            .O(N__5917),
            .I(\U409_TICK.TICK503_8_cascade_ ));
    CascadeMux I__1269 (
            .O(N__5914),
            .I(\U409_TICK.TICK503_14_cascade_ ));
    InMux I__1268 (
            .O(N__5911),
            .I(N__5895));
    InMux I__1267 (
            .O(N__5910),
            .I(N__5895));
    InMux I__1266 (
            .O(N__5909),
            .I(N__5895));
    InMux I__1265 (
            .O(N__5908),
            .I(N__5895));
    InMux I__1264 (
            .O(N__5907),
            .I(N__5886));
    InMux I__1263 (
            .O(N__5906),
            .I(N__5886));
    InMux I__1262 (
            .O(N__5905),
            .I(N__5886));
    InMux I__1261 (
            .O(N__5904),
            .I(N__5886));
    LocalMux I__1260 (
            .O(N__5895),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__1259 (
            .O(N__5886),
            .I(\U409_TICK.TICK503_14 ));
    InMux I__1258 (
            .O(N__5881),
            .I(N__5863));
    InMux I__1257 (
            .O(N__5880),
            .I(N__5863));
    InMux I__1256 (
            .O(N__5879),
            .I(N__5863));
    InMux I__1255 (
            .O(N__5878),
            .I(N__5863));
    InMux I__1254 (
            .O(N__5877),
            .I(N__5863));
    InMux I__1253 (
            .O(N__5876),
            .I(N__5856));
    InMux I__1252 (
            .O(N__5875),
            .I(N__5856));
    InMux I__1251 (
            .O(N__5874),
            .I(N__5856));
    LocalMux I__1250 (
            .O(N__5863),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__1249 (
            .O(N__5856),
            .I(\U409_TICK.TICK503_10 ));
    CascadeMux I__1248 (
            .O(N__5851),
            .I(N__5846));
    InMux I__1247 (
            .O(N__5850),
            .I(N__5833));
    InMux I__1246 (
            .O(N__5849),
            .I(N__5833));
    InMux I__1245 (
            .O(N__5846),
            .I(N__5833));
    InMux I__1244 (
            .O(N__5845),
            .I(N__5833));
    CascadeMux I__1243 (
            .O(N__5844),
            .I(N__5829));
    CascadeMux I__1242 (
            .O(N__5843),
            .I(N__5826));
    InMux I__1241 (
            .O(N__5842),
            .I(N__5823));
    LocalMux I__1240 (
            .O(N__5833),
            .I(N__5820));
    InMux I__1239 (
            .O(N__5832),
            .I(N__5813));
    InMux I__1238 (
            .O(N__5829),
            .I(N__5813));
    InMux I__1237 (
            .O(N__5826),
            .I(N__5813));
    LocalMux I__1236 (
            .O(N__5823),
            .I(\U409_TICK.TICK503_9 ));
    Odrv4 I__1235 (
            .O(N__5820),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__1234 (
            .O(N__5813),
            .I(\U409_TICK.TICK503_9 ));
    IoInMux I__1233 (
            .O(N__5806),
            .I(N__5803));
    LocalMux I__1232 (
            .O(N__5803),
            .I(N__5800));
    Span4Mux_s0_v I__1231 (
            .O(N__5800),
            .I(N__5797));
    Span4Mux_v I__1230 (
            .O(N__5797),
            .I(N__5794));
    Span4Mux_v I__1229 (
            .O(N__5794),
            .I(N__5791));
    Span4Mux_v I__1228 (
            .O(N__5791),
            .I(N__5787));
    InMux I__1227 (
            .O(N__5790),
            .I(N__5784));
    Odrv4 I__1226 (
            .O(N__5787),
            .I(TICK60_c));
    LocalMux I__1225 (
            .O(N__5784),
            .I(TICK60_c));
    CascadeMux I__1224 (
            .O(N__5779),
            .I(\U409_TICK.TICK603_9_cascade_ ));
    CascadeMux I__1223 (
            .O(N__5776),
            .I(N__5770));
    CascadeMux I__1222 (
            .O(N__5775),
            .I(N__5767));
    InMux I__1221 (
            .O(N__5774),
            .I(N__5755));
    InMux I__1220 (
            .O(N__5773),
            .I(N__5755));
    InMux I__1219 (
            .O(N__5770),
            .I(N__5755));
    InMux I__1218 (
            .O(N__5767),
            .I(N__5755));
    InMux I__1217 (
            .O(N__5766),
            .I(N__5748));
    InMux I__1216 (
            .O(N__5765),
            .I(N__5748));
    InMux I__1215 (
            .O(N__5764),
            .I(N__5748));
    LocalMux I__1214 (
            .O(N__5755),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__1213 (
            .O(N__5748),
            .I(\U409_TICK.TICK603_9 ));
    CascadeMux I__1212 (
            .O(N__5743),
            .I(N__5740));
    InMux I__1211 (
            .O(N__5740),
            .I(N__5737));
    LocalMux I__1210 (
            .O(N__5737),
            .I(N__5728));
    InMux I__1209 (
            .O(N__5736),
            .I(N__5721));
    InMux I__1208 (
            .O(N__5735),
            .I(N__5721));
    InMux I__1207 (
            .O(N__5734),
            .I(N__5721));
    InMux I__1206 (
            .O(N__5733),
            .I(N__5714));
    InMux I__1205 (
            .O(N__5732),
            .I(N__5714));
    InMux I__1204 (
            .O(N__5731),
            .I(N__5714));
    Odrv4 I__1203 (
            .O(N__5728),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__1202 (
            .O(N__5721),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__1201 (
            .O(N__5714),
            .I(\U409_TICK.TICK603_14 ));
    CascadeMux I__1200 (
            .O(N__5707),
            .I(N__5703));
    InMux I__1199 (
            .O(N__5706),
            .I(N__5689));
    InMux I__1198 (
            .O(N__5703),
            .I(N__5689));
    InMux I__1197 (
            .O(N__5702),
            .I(N__5689));
    InMux I__1196 (
            .O(N__5701),
            .I(N__5689));
    InMux I__1195 (
            .O(N__5700),
            .I(N__5682));
    InMux I__1194 (
            .O(N__5699),
            .I(N__5682));
    InMux I__1193 (
            .O(N__5698),
            .I(N__5682));
    LocalMux I__1192 (
            .O(N__5689),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__1191 (
            .O(N__5682),
            .I(\U409_TICK.TICK603_10 ));
    IoInMux I__1190 (
            .O(N__5677),
            .I(N__5674));
    LocalMux I__1189 (
            .O(N__5674),
            .I(N__5671));
    Span4Mux_s1_v I__1188 (
            .O(N__5671),
            .I(N__5668));
    Sp12to4 I__1187 (
            .O(N__5668),
            .I(N__5665));
    Span12Mux_h I__1186 (
            .O(N__5665),
            .I(N__5661));
    InMux I__1185 (
            .O(N__5664),
            .I(N__5658));
    Odrv12 I__1184 (
            .O(N__5661),
            .I(TICK50_c));
    LocalMux I__1183 (
            .O(N__5658),
            .I(TICK50_c));
    CascadeMux I__1182 (
            .O(N__5653),
            .I(\U409_TICK.TICK503_9_cascade_ ));
    SRMux I__1181 (
            .O(N__5650),
            .I(N__5646));
    SRMux I__1180 (
            .O(N__5649),
            .I(N__5642));
    LocalMux I__1179 (
            .O(N__5646),
            .I(N__5637));
    SRMux I__1178 (
            .O(N__5645),
            .I(N__5634));
    LocalMux I__1177 (
            .O(N__5642),
            .I(N__5631));
    SRMux I__1176 (
            .O(N__5641),
            .I(N__5628));
    SRMux I__1175 (
            .O(N__5640),
            .I(N__5625));
    Span4Mux_v I__1174 (
            .O(N__5637),
            .I(N__5621));
    LocalMux I__1173 (
            .O(N__5634),
            .I(N__5618));
    Span4Mux_v I__1172 (
            .O(N__5631),
            .I(N__5615));
    LocalMux I__1171 (
            .O(N__5628),
            .I(N__5612));
    LocalMux I__1170 (
            .O(N__5625),
            .I(N__5609));
    SRMux I__1169 (
            .O(N__5624),
            .I(N__5606));
    Odrv4 I__1168 (
            .O(N__5621),
            .I(RESETn_c_i));
    Odrv4 I__1167 (
            .O(N__5618),
            .I(RESETn_c_i));
    Odrv4 I__1166 (
            .O(N__5615),
            .I(RESETn_c_i));
    Odrv12 I__1165 (
            .O(N__5612),
            .I(RESETn_c_i));
    Odrv12 I__1164 (
            .O(N__5609),
            .I(RESETn_c_i));
    LocalMux I__1163 (
            .O(N__5606),
            .I(RESETn_c_i));
    CascadeMux I__1162 (
            .O(N__5593),
            .I(\U409_TICK.TICK603_8_cascade_ ));
    CascadeMux I__1161 (
            .O(N__5590),
            .I(\U409_TICK.TICK603_14_cascade_ ));
    InMux I__1160 (
            .O(N__5587),
            .I(N__5584));
    LocalMux I__1159 (
            .O(N__5584),
            .I(\U409_TICK.TICK603_11 ));
    CascadeMux I__1158 (
            .O(N__5581),
            .I(\U409_TICK.TICK603_10_cascade_ ));
    CascadeMux I__1157 (
            .O(N__5578),
            .I(\U409_TICK.TICK503_10_cascade_ ));
    CascadeMux I__1156 (
            .O(N__5575),
            .I(N__5570));
    InMux I__1155 (
            .O(N__5574),
            .I(N__5565));
    InMux I__1154 (
            .O(N__5573),
            .I(N__5562));
    InMux I__1153 (
            .O(N__5570),
            .I(N__5555));
    InMux I__1152 (
            .O(N__5569),
            .I(N__5555));
    InMux I__1151 (
            .O(N__5568),
            .I(N__5555));
    LocalMux I__1150 (
            .O(N__5565),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__1149 (
            .O(N__5562),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__1148 (
            .O(N__5555),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    CascadeMux I__1147 (
            .O(N__5548),
            .I(N__5541));
    InMux I__1146 (
            .O(N__5547),
            .I(N__5536));
    InMux I__1145 (
            .O(N__5546),
            .I(N__5536));
    InMux I__1144 (
            .O(N__5545),
            .I(N__5533));
    InMux I__1143 (
            .O(N__5544),
            .I(N__5528));
    InMux I__1142 (
            .O(N__5541),
            .I(N__5528));
    LocalMux I__1141 (
            .O(N__5536),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1140 (
            .O(N__5533),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1139 (
            .O(N__5528),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    InMux I__1138 (
            .O(N__5521),
            .I(N__5508));
    InMux I__1137 (
            .O(N__5520),
            .I(N__5508));
    InMux I__1136 (
            .O(N__5519),
            .I(N__5508));
    InMux I__1135 (
            .O(N__5518),
            .I(N__5505));
    InMux I__1134 (
            .O(N__5517),
            .I(N__5502));
    InMux I__1133 (
            .O(N__5516),
            .I(N__5497));
    InMux I__1132 (
            .O(N__5515),
            .I(N__5497));
    LocalMux I__1131 (
            .O(N__5508),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1130 (
            .O(N__5505),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1129 (
            .O(N__5502),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1128 (
            .O(N__5497),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    InMux I__1127 (
            .O(N__5488),
            .I(N__5482));
    InMux I__1126 (
            .O(N__5487),
            .I(N__5479));
    InMux I__1125 (
            .O(N__5486),
            .I(N__5474));
    InMux I__1124 (
            .O(N__5485),
            .I(N__5474));
    LocalMux I__1123 (
            .O(N__5482),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1122 (
            .O(N__5479),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1121 (
            .O(N__5474),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    SRMux I__1120 (
            .O(N__5467),
            .I(N__5463));
    SRMux I__1119 (
            .O(N__5466),
            .I(N__5459));
    LocalMux I__1118 (
            .O(N__5463),
            .I(N__5456));
    SRMux I__1117 (
            .O(N__5462),
            .I(N__5453));
    LocalMux I__1116 (
            .O(N__5459),
            .I(N__5449));
    Span4Mux_v I__1115 (
            .O(N__5456),
            .I(N__5444));
    LocalMux I__1114 (
            .O(N__5453),
            .I(N__5444));
    SRMux I__1113 (
            .O(N__5452),
            .I(N__5441));
    Span4Mux_v I__1112 (
            .O(N__5449),
            .I(N__5436));
    Span4Mux_h I__1111 (
            .O(N__5444),
            .I(N__5436));
    LocalMux I__1110 (
            .O(N__5441),
            .I(N__5433));
    Odrv4 I__1109 (
            .O(N__5436),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    Odrv4 I__1108 (
            .O(N__5433),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    InMux I__1107 (
            .O(N__5428),
            .I(N__5425));
    LocalMux I__1106 (
            .O(N__5425),
            .I(N__5422));
    Span4Mux_v I__1105 (
            .O(N__5422),
            .I(N__5419));
    Sp12to4 I__1104 (
            .O(N__5419),
            .I(N__5416));
    Span12Mux_h I__1103 (
            .O(N__5416),
            .I(N__5413));
    Odrv12 I__1102 (
            .O(N__5413),
            .I(A_c_13));
    IoInMux I__1101 (
            .O(N__5410),
            .I(N__5407));
    LocalMux I__1100 (
            .O(N__5407),
            .I(N__5404));
    IoSpan4Mux I__1099 (
            .O(N__5404),
            .I(N__5401));
    IoSpan4Mux I__1098 (
            .O(N__5401),
            .I(N__5398));
    Sp12to4 I__1097 (
            .O(N__5398),
            .I(N__5395));
    Span12Mux_s7_h I__1096 (
            .O(N__5395),
            .I(N__5392));
    Odrv12 I__1095 (
            .O(N__5392),
            .I(U409_ADDRESS_DECODE_un1_CIACS1n_i));
    InMux I__1094 (
            .O(N__5389),
            .I(N__5386));
    LocalMux I__1093 (
            .O(N__5386),
            .I(N__5383));
    Span4Mux_v I__1092 (
            .O(N__5383),
            .I(N__5380));
    Sp12to4 I__1091 (
            .O(N__5380),
            .I(N__5377));
    Span12Mux_h I__1090 (
            .O(N__5377),
            .I(N__5374));
    Odrv12 I__1089 (
            .O(N__5374),
            .I(A_c_12));
    IoInMux I__1088 (
            .O(N__5371),
            .I(N__5368));
    LocalMux I__1087 (
            .O(N__5368),
            .I(N__5365));
    IoSpan4Mux I__1086 (
            .O(N__5365),
            .I(N__5362));
    IoSpan4Mux I__1085 (
            .O(N__5362),
            .I(N__5359));
    Span4Mux_s2_h I__1084 (
            .O(N__5359),
            .I(N__5356));
    Sp12to4 I__1083 (
            .O(N__5356),
            .I(N__5353));
    Odrv12 I__1082 (
            .O(N__5353),
            .I(U409_ADDRESS_DECODE_un1_CIACS0n_i));
    InMux I__1081 (
            .O(N__5350),
            .I(N__5344));
    InMux I__1080 (
            .O(N__5349),
            .I(N__5344));
    LocalMux I__1079 (
            .O(N__5344),
            .I(CIA_ENABLE));
    CascadeMux I__1078 (
            .O(N__5341),
            .I(N__5336));
    InMux I__1077 (
            .O(N__5340),
            .I(N__5332));
    InMux I__1076 (
            .O(N__5339),
            .I(N__5329));
    InMux I__1075 (
            .O(N__5336),
            .I(N__5325));
    InMux I__1074 (
            .O(N__5335),
            .I(N__5322));
    LocalMux I__1073 (
            .O(N__5332),
            .I(N__5319));
    LocalMux I__1072 (
            .O(N__5329),
            .I(N__5316));
    InMux I__1071 (
            .O(N__5328),
            .I(N__5313));
    LocalMux I__1070 (
            .O(N__5325),
            .I(N__5307));
    LocalMux I__1069 (
            .O(N__5322),
            .I(N__5307));
    Span4Mux_h I__1068 (
            .O(N__5319),
            .I(N__5304));
    Span4Mux_v I__1067 (
            .O(N__5316),
            .I(N__5301));
    LocalMux I__1066 (
            .O(N__5313),
            .I(N__5298));
    CascadeMux I__1065 (
            .O(N__5312),
            .I(N__5295));
    Span4Mux_v I__1064 (
            .O(N__5307),
            .I(N__5292));
    Span4Mux_h I__1063 (
            .O(N__5304),
            .I(N__5288));
    Span4Mux_h I__1062 (
            .O(N__5301),
            .I(N__5283));
    Span4Mux_v I__1061 (
            .O(N__5298),
            .I(N__5283));
    InMux I__1060 (
            .O(N__5295),
            .I(N__5280));
    Span4Mux_h I__1059 (
            .O(N__5292),
            .I(N__5273));
    InMux I__1058 (
            .O(N__5291),
            .I(N__5270));
    Span4Mux_h I__1057 (
            .O(N__5288),
            .I(N__5264));
    Span4Mux_h I__1056 (
            .O(N__5283),
            .I(N__5259));
    LocalMux I__1055 (
            .O(N__5280),
            .I(N__5259));
    InMux I__1054 (
            .O(N__5279),
            .I(N__5250));
    InMux I__1053 (
            .O(N__5278),
            .I(N__5250));
    InMux I__1052 (
            .O(N__5277),
            .I(N__5250));
    InMux I__1051 (
            .O(N__5276),
            .I(N__5250));
    Span4Mux_v I__1050 (
            .O(N__5273),
            .I(N__5244));
    LocalMux I__1049 (
            .O(N__5270),
            .I(N__5244));
    InMux I__1048 (
            .O(N__5269),
            .I(N__5241));
    InMux I__1047 (
            .O(N__5268),
            .I(N__5238));
    InMux I__1046 (
            .O(N__5267),
            .I(N__5235));
    Span4Mux_v I__1045 (
            .O(N__5264),
            .I(N__5232));
    Span4Mux_v I__1044 (
            .O(N__5259),
            .I(N__5227));
    LocalMux I__1043 (
            .O(N__5250),
            .I(N__5227));
    InMux I__1042 (
            .O(N__5249),
            .I(N__5224));
    Span4Mux_h I__1041 (
            .O(N__5244),
            .I(N__5219));
    LocalMux I__1040 (
            .O(N__5241),
            .I(N__5219));
    LocalMux I__1039 (
            .O(N__5238),
            .I(N__5214));
    LocalMux I__1038 (
            .O(N__5235),
            .I(N__5214));
    Sp12to4 I__1037 (
            .O(N__5232),
            .I(N__5207));
    Sp12to4 I__1036 (
            .O(N__5227),
            .I(N__5207));
    LocalMux I__1035 (
            .O(N__5224),
            .I(N__5207));
    Span4Mux_v I__1034 (
            .O(N__5219),
            .I(N__5202));
    Span4Mux_v I__1033 (
            .O(N__5214),
            .I(N__5202));
    Span12Mux_v I__1032 (
            .O(N__5207),
            .I(N__5199));
    Sp12to4 I__1031 (
            .O(N__5202),
            .I(N__5196));
    Span12Mux_h I__1030 (
            .O(N__5199),
            .I(N__5193));
    Span12Mux_h I__1029 (
            .O(N__5196),
            .I(N__5190));
    Odrv12 I__1028 (
            .O(N__5193),
            .I(RESETn_c));
    Odrv12 I__1027 (
            .O(N__5190),
            .I(RESETn_c));
    InMux I__1026 (
            .O(N__5185),
            .I(N__5180));
    InMux I__1025 (
            .O(N__5184),
            .I(N__5175));
    InMux I__1024 (
            .O(N__5183),
            .I(N__5175));
    LocalMux I__1023 (
            .O(N__5180),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    LocalMux I__1022 (
            .O(N__5175),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    InMux I__1021 (
            .O(N__5170),
            .I(N__5164));
    InMux I__1020 (
            .O(N__5169),
            .I(N__5164));
    LocalMux I__1019 (
            .O(N__5164),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    InMux I__1018 (
            .O(N__5161),
            .I(N__5158));
    LocalMux I__1017 (
            .O(N__5158),
            .I(\U409_TRANSFER_ACK.N_3_0 ));
    CascadeMux I__1016 (
            .O(N__5155),
            .I(\U409_TRANSFER_ACK.N_3_0_cascade_ ));
    CascadeMux I__1015 (
            .O(N__5152),
            .I(N__5147));
    InMux I__1014 (
            .O(N__5151),
            .I(N__5144));
    InMux I__1013 (
            .O(N__5150),
            .I(N__5141));
    InMux I__1012 (
            .O(N__5147),
            .I(N__5138));
    LocalMux I__1011 (
            .O(N__5144),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__1010 (
            .O(N__5141),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__1009 (
            .O(N__5138),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    CascadeMux I__1008 (
            .O(N__5131),
            .I(\U409_TRANSFER_ACK.N_6_0_cascade_ ));
    CascadeMux I__1007 (
            .O(N__5128),
            .I(N__5125));
    InMux I__1006 (
            .O(N__5125),
            .I(N__5120));
    CascadeMux I__1005 (
            .O(N__5124),
            .I(N__5116));
    InMux I__1004 (
            .O(N__5123),
            .I(N__5112));
    LocalMux I__1003 (
            .O(N__5120),
            .I(N__5109));
    InMux I__1002 (
            .O(N__5119),
            .I(N__5102));
    InMux I__1001 (
            .O(N__5116),
            .I(N__5102));
    InMux I__1000 (
            .O(N__5115),
            .I(N__5102));
    LocalMux I__999 (
            .O(N__5112),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    Odrv4 I__998 (
            .O(N__5109),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__997 (
            .O(N__5102),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    InMux I__996 (
            .O(N__5095),
            .I(N__5089));
    InMux I__995 (
            .O(N__5094),
            .I(N__5086));
    InMux I__994 (
            .O(N__5093),
            .I(N__5081));
    InMux I__993 (
            .O(N__5092),
            .I(N__5081));
    LocalMux I__992 (
            .O(N__5089),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__991 (
            .O(N__5086),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__990 (
            .O(N__5081),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    InMux I__989 (
            .O(N__5074),
            .I(N__5069));
    InMux I__988 (
            .O(N__5073),
            .I(N__5066));
    InMux I__987 (
            .O(N__5072),
            .I(N__5063));
    LocalMux I__986 (
            .O(N__5069),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    LocalMux I__985 (
            .O(N__5066),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    LocalMux I__984 (
            .O(N__5063),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    InMux I__983 (
            .O(N__5056),
            .I(N__5050));
    InMux I__982 (
            .O(N__5055),
            .I(N__5050));
    LocalMux I__981 (
            .O(N__5050),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ));
    InMux I__980 (
            .O(N__5047),
            .I(N__5041));
    InMux I__979 (
            .O(N__5046),
            .I(N__5038));
    InMux I__978 (
            .O(N__5045),
            .I(N__5035));
    InMux I__977 (
            .O(N__5044),
            .I(N__5032));
    LocalMux I__976 (
            .O(N__5041),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__975 (
            .O(N__5038),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__974 (
            .O(N__5035),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__973 (
            .O(N__5032),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    CascadeMux I__972 (
            .O(N__5023),
            .I(N__5016));
    InMux I__971 (
            .O(N__5022),
            .I(N__5013));
    InMux I__970 (
            .O(N__5021),
            .I(N__5010));
    InMux I__969 (
            .O(N__5020),
            .I(N__5007));
    InMux I__968 (
            .O(N__5019),
            .I(N__5002));
    InMux I__967 (
            .O(N__5016),
            .I(N__5002));
    LocalMux I__966 (
            .O(N__5013),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__965 (
            .O(N__5010),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__964 (
            .O(N__5007),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__963 (
            .O(N__5002),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    CascadeMux I__962 (
            .O(N__4993),
            .I(N__4987));
    InMux I__961 (
            .O(N__4992),
            .I(N__4980));
    InMux I__960 (
            .O(N__4991),
            .I(N__4980));
    InMux I__959 (
            .O(N__4990),
            .I(N__4977));
    InMux I__958 (
            .O(N__4987),
            .I(N__4974));
    InMux I__957 (
            .O(N__4986),
            .I(N__4971));
    InMux I__956 (
            .O(N__4985),
            .I(N__4968));
    LocalMux I__955 (
            .O(N__4980),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__954 (
            .O(N__4977),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__953 (
            .O(N__4974),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__952 (
            .O(N__4971),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__951 (
            .O(N__4968),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    CascadeMux I__950 (
            .O(N__4957),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1_cascade_ ));
    CascadeMux I__949 (
            .O(N__4954),
            .I(N__4951));
    InMux I__948 (
            .O(N__4951),
            .I(N__4945));
    InMux I__947 (
            .O(N__4950),
            .I(N__4945));
    LocalMux I__946 (
            .O(N__4945),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ));
    InMux I__945 (
            .O(N__4942),
            .I(N__4939));
    LocalMux I__944 (
            .O(N__4939),
            .I(N__4935));
    InMux I__943 (
            .O(N__4938),
            .I(N__4932));
    Span4Mux_v I__942 (
            .O(N__4935),
            .I(N__4925));
    LocalMux I__941 (
            .O(N__4932),
            .I(N__4925));
    InMux I__940 (
            .O(N__4931),
            .I(N__4922));
    InMux I__939 (
            .O(N__4930),
            .I(N__4919));
    Span4Mux_h I__938 (
            .O(N__4925),
            .I(N__4913));
    LocalMux I__937 (
            .O(N__4922),
            .I(N__4913));
    LocalMux I__936 (
            .O(N__4919),
            .I(N__4910));
    CascadeMux I__935 (
            .O(N__4918),
            .I(N__4907));
    Span4Mux_v I__934 (
            .O(N__4913),
            .I(N__4904));
    Span4Mux_v I__933 (
            .O(N__4910),
            .I(N__4901));
    InMux I__932 (
            .O(N__4907),
            .I(N__4898));
    Sp12to4 I__931 (
            .O(N__4904),
            .I(N__4891));
    Sp12to4 I__930 (
            .O(N__4901),
            .I(N__4891));
    LocalMux I__929 (
            .O(N__4898),
            .I(N__4891));
    Span12Mux_h I__928 (
            .O(N__4891),
            .I(N__4888));
    Span12Mux_v I__927 (
            .O(N__4888),
            .I(N__4885));
    Odrv12 I__926 (
            .O(N__4885),
            .I(TSn_c));
    IoInMux I__925 (
            .O(N__4882),
            .I(N__4879));
    LocalMux I__924 (
            .O(N__4879),
            .I(N__4875));
    InMux I__923 (
            .O(N__4878),
            .I(N__4872));
    IoSpan4Mux I__922 (
            .O(N__4875),
            .I(N__4868));
    LocalMux I__921 (
            .O(N__4872),
            .I(N__4865));
    InMux I__920 (
            .O(N__4871),
            .I(N__4862));
    Span4Mux_s0_v I__919 (
            .O(N__4868),
            .I(N__4856));
    Span4Mux_v I__918 (
            .O(N__4865),
            .I(N__4853));
    LocalMux I__917 (
            .O(N__4862),
            .I(N__4850));
    InMux I__916 (
            .O(N__4861),
            .I(N__4847));
    CascadeMux I__915 (
            .O(N__4860),
            .I(N__4844));
    InMux I__914 (
            .O(N__4859),
            .I(N__4841));
    Sp12to4 I__913 (
            .O(N__4856),
            .I(N__4837));
    Sp12to4 I__912 (
            .O(N__4853),
            .I(N__4834));
    Span4Mux_h I__911 (
            .O(N__4850),
            .I(N__4829));
    LocalMux I__910 (
            .O(N__4847),
            .I(N__4829));
    InMux I__909 (
            .O(N__4844),
            .I(N__4826));
    LocalMux I__908 (
            .O(N__4841),
            .I(N__4823));
    InMux I__907 (
            .O(N__4840),
            .I(N__4820));
    Span12Mux_v I__906 (
            .O(N__4837),
            .I(N__4811));
    Span12Mux_h I__905 (
            .O(N__4834),
            .I(N__4811));
    Sp12to4 I__904 (
            .O(N__4829),
            .I(N__4811));
    LocalMux I__903 (
            .O(N__4826),
            .I(N__4811));
    Span12Mux_h I__902 (
            .O(N__4823),
            .I(N__4808));
    LocalMux I__901 (
            .O(N__4820),
            .I(N__4805));
    Span12Mux_v I__900 (
            .O(N__4811),
            .I(N__4802));
    Span12Mux_v I__899 (
            .O(N__4808),
            .I(N__4799));
    Span12Mux_v I__898 (
            .O(N__4805),
            .I(N__4796));
    Odrv12 I__897 (
            .O(N__4802),
            .I(CLK40_IN_c));
    Odrv12 I__896 (
            .O(N__4799),
            .I(CLK40_IN_c));
    Odrv12 I__895 (
            .O(N__4796),
            .I(CLK40_IN_c));
    InMux I__894 (
            .O(N__4789),
            .I(N__4785));
    InMux I__893 (
            .O(N__4788),
            .I(N__4782));
    LocalMux I__892 (
            .O(N__4785),
            .I(\U409_TRANSFER_ACK.N_70 ));
    LocalMux I__891 (
            .O(N__4782),
            .I(\U409_TRANSFER_ACK.N_70 ));
    InMux I__890 (
            .O(N__4777),
            .I(N__4771));
    InMux I__889 (
            .O(N__4776),
            .I(N__4771));
    LocalMux I__888 (
            .O(N__4771),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ));
    CascadeMux I__887 (
            .O(N__4768),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ));
    InMux I__886 (
            .O(N__4765),
            .I(N__4762));
    LocalMux I__885 (
            .O(N__4762),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out ));
    IoInMux I__884 (
            .O(N__4759),
            .I(N__4756));
    LocalMux I__883 (
            .O(N__4756),
            .I(N__4753));
    Span4Mux_s3_v I__882 (
            .O(N__4753),
            .I(N__4750));
    Span4Mux_h I__881 (
            .O(N__4750),
            .I(N__4747));
    Odrv4 I__880 (
            .O(N__4747),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__879 (
            .O(N__4744),
            .I(N__4741));
    InMux I__878 (
            .O(N__4741),
            .I(N__4737));
    InMux I__877 (
            .O(N__4740),
            .I(N__4734));
    LocalMux I__876 (
            .O(N__4737),
            .I(N__4731));
    LocalMux I__875 (
            .O(N__4734),
            .I(\U409_TRANSFER_ACK.CO1 ));
    Odrv4 I__874 (
            .O(N__4731),
            .I(\U409_TRANSFER_ACK.CO1 ));
    InMux I__873 (
            .O(N__4726),
            .I(N__4723));
    LocalMux I__872 (
            .O(N__4723),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0 ));
    CascadeMux I__871 (
            .O(N__4720),
            .I(N__4714));
    InMux I__870 (
            .O(N__4719),
            .I(N__4711));
    InMux I__869 (
            .O(N__4718),
            .I(N__4708));
    InMux I__868 (
            .O(N__4717),
            .I(N__4703));
    InMux I__867 (
            .O(N__4714),
            .I(N__4703));
    LocalMux I__866 (
            .O(N__4711),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__865 (
            .O(N__4708),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__864 (
            .O(N__4703),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    CascadeMux I__863 (
            .O(N__4696),
            .I(N__4690));
    InMux I__862 (
            .O(N__4695),
            .I(N__4686));
    InMux I__861 (
            .O(N__4694),
            .I(N__4683));
    InMux I__860 (
            .O(N__4693),
            .I(N__4680));
    InMux I__859 (
            .O(N__4690),
            .I(N__4675));
    InMux I__858 (
            .O(N__4689),
            .I(N__4675));
    LocalMux I__857 (
            .O(N__4686),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__856 (
            .O(N__4683),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__855 (
            .O(N__4680),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__854 (
            .O(N__4675),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    CascadeMux I__853 (
            .O(N__4666),
            .I(N__4663));
    InMux I__852 (
            .O(N__4663),
            .I(N__4660));
    LocalMux I__851 (
            .O(N__4660),
            .I(\U409_TRANSFER_ACK.ROM_TACK_EN_e_1 ));
    InMux I__850 (
            .O(N__4657),
            .I(N__4654));
    LocalMux I__849 (
            .O(N__4654),
            .I(\U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0 ));
    InMux I__848 (
            .O(N__4651),
            .I(N__4647));
    InMux I__847 (
            .O(N__4650),
            .I(N__4644));
    LocalMux I__846 (
            .O(N__4647),
            .I(\U409_TRANSFER_ACK.N_17_mux ));
    LocalMux I__845 (
            .O(N__4644),
            .I(\U409_TRANSFER_ACK.N_17_mux ));
    InMux I__844 (
            .O(N__4639),
            .I(N__4635));
    InMux I__843 (
            .O(N__4638),
            .I(N__4632));
    LocalMux I__842 (
            .O(N__4635),
            .I(N__4629));
    LocalMux I__841 (
            .O(N__4632),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    Odrv4 I__840 (
            .O(N__4629),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    CascadeMux I__839 (
            .O(N__4624),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3_cascade_ ));
    CascadeMux I__838 (
            .O(N__4621),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a4_3_cascade_ ));
    CascadeMux I__837 (
            .O(N__4618),
            .I(\U409_TRANSFER_ACK.N_70_cascade_ ));
    InMux I__836 (
            .O(N__4615),
            .I(N__4611));
    InMux I__835 (
            .O(N__4614),
            .I(N__4608));
    LocalMux I__834 (
            .O(N__4611),
            .I(\U409_TRANSFER_ACK.N_55 ));
    LocalMux I__833 (
            .O(N__4608),
            .I(\U409_TRANSFER_ACK.N_55 ));
    CascadeMux I__832 (
            .O(N__4603),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ));
    CascadeMux I__831 (
            .O(N__4600),
            .I(N__4596));
    InMux I__830 (
            .O(N__4599),
            .I(N__4589));
    InMux I__829 (
            .O(N__4596),
            .I(N__4589));
    InMux I__828 (
            .O(N__4595),
            .I(N__4584));
    InMux I__827 (
            .O(N__4594),
            .I(N__4584));
    LocalMux I__826 (
            .O(N__4589),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__825 (
            .O(N__4584),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    InMux I__824 (
            .O(N__4579),
            .I(N__4570));
    InMux I__823 (
            .O(N__4578),
            .I(N__4570));
    InMux I__822 (
            .O(N__4577),
            .I(N__4570));
    LocalMux I__821 (
            .O(N__4570),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    CascadeMux I__820 (
            .O(N__4567),
            .I(\U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_ ));
    InMux I__819 (
            .O(N__4564),
            .I(N__4560));
    InMux I__818 (
            .O(N__4563),
            .I(N__4557));
    LocalMux I__817 (
            .O(N__4560),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    LocalMux I__816 (
            .O(N__4557),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    InMux I__815 (
            .O(N__4552),
            .I(N__4548));
    InMux I__814 (
            .O(N__4551),
            .I(N__4545));
    LocalMux I__813 (
            .O(N__4548),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    LocalMux I__812 (
            .O(N__4545),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    CascadeMux I__811 (
            .O(N__4540),
            .I(N__4536));
    InMux I__810 (
            .O(N__4539),
            .I(N__4533));
    InMux I__809 (
            .O(N__4536),
            .I(N__4530));
    LocalMux I__808 (
            .O(N__4533),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    LocalMux I__807 (
            .O(N__4530),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    CascadeMux I__806 (
            .O(N__4525),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ));
    CascadeMux I__805 (
            .O(N__4522),
            .I(\U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ));
    IoInMux I__804 (
            .O(N__4519),
            .I(N__4516));
    LocalMux I__803 (
            .O(N__4516),
            .I(N__4513));
    Span12Mux_s7_v I__802 (
            .O(N__4513),
            .I(N__4510));
    Span12Mux_v I__801 (
            .O(N__4510),
            .I(N__4507));
    Span12Mux_h I__800 (
            .O(N__4507),
            .I(N__4502));
    InMux I__799 (
            .O(N__4506),
            .I(N__4497));
    InMux I__798 (
            .O(N__4505),
            .I(N__4497));
    Odrv12 I__797 (
            .O(N__4502),
            .I(TACK_OUTn));
    LocalMux I__796 (
            .O(N__4497),
            .I(TACK_OUTn));
    CascadeMux I__795 (
            .O(N__4492),
            .I(N__4487));
    CascadeMux I__794 (
            .O(N__4491),
            .I(N__4483));
    InMux I__793 (
            .O(N__4490),
            .I(N__4479));
    InMux I__792 (
            .O(N__4487),
            .I(N__4472));
    InMux I__791 (
            .O(N__4486),
            .I(N__4472));
    InMux I__790 (
            .O(N__4483),
            .I(N__4472));
    InMux I__789 (
            .O(N__4482),
            .I(N__4469));
    LocalMux I__788 (
            .O(N__4479),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    LocalMux I__787 (
            .O(N__4472),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    LocalMux I__786 (
            .O(N__4469),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    InMux I__785 (
            .O(N__4462),
            .I(N__4455));
    InMux I__784 (
            .O(N__4461),
            .I(N__4446));
    InMux I__783 (
            .O(N__4460),
            .I(N__4446));
    InMux I__782 (
            .O(N__4459),
            .I(N__4446));
    InMux I__781 (
            .O(N__4458),
            .I(N__4446));
    LocalMux I__780 (
            .O(N__4455),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    LocalMux I__779 (
            .O(N__4446),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    InMux I__778 (
            .O(N__4441),
            .I(N__4436));
    InMux I__777 (
            .O(N__4440),
            .I(N__4431));
    InMux I__776 (
            .O(N__4439),
            .I(N__4431));
    LocalMux I__775 (
            .O(N__4436),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    LocalMux I__774 (
            .O(N__4431),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    CEMux I__773 (
            .O(N__4426),
            .I(N__4423));
    LocalMux I__772 (
            .O(N__4423),
            .I(N__4420));
    Span4Mux_v I__771 (
            .O(N__4420),
            .I(N__4417));
    Span4Mux_h I__770 (
            .O(N__4417),
            .I(N__4414));
    Odrv4 I__769 (
            .O(N__4414),
            .I(\U409_TRANSFER_ACK.TACK_OUTn_0_sqmuxa_0_en ));
    CascadeMux I__768 (
            .O(N__4411),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20_cascade_ ));
    CascadeMux I__767 (
            .O(N__4408),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_cascade_ ));
    CascadeMux I__766 (
            .O(N__4405),
            .I(N__4402));
    InMux I__765 (
            .O(N__4402),
            .I(N__4395));
    InMux I__764 (
            .O(N__4401),
            .I(N__4395));
    InMux I__763 (
            .O(N__4400),
            .I(N__4392));
    LocalMux I__762 (
            .O(N__4395),
            .I(N__4389));
    LocalMux I__761 (
            .O(N__4392),
            .I(N__4386));
    Span4Mux_h I__760 (
            .O(N__4389),
            .I(N__4383));
    Span4Mux_v I__759 (
            .O(N__4386),
            .I(N__4380));
    Span4Mux_v I__758 (
            .O(N__4383),
            .I(N__4377));
    Odrv4 I__757 (
            .O(N__4380),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15 ));
    Odrv4 I__756 (
            .O(N__4377),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15 ));
    InMux I__755 (
            .O(N__4372),
            .I(N__4368));
    InMux I__754 (
            .O(N__4371),
            .I(N__4365));
    LocalMux I__753 (
            .O(N__4368),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20 ));
    LocalMux I__752 (
            .O(N__4365),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20 ));
    InMux I__751 (
            .O(N__4360),
            .I(N__4356));
    InMux I__750 (
            .O(N__4359),
            .I(N__4353));
    LocalMux I__749 (
            .O(N__4356),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ));
    LocalMux I__748 (
            .O(N__4353),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ));
    IoInMux I__747 (
            .O(N__4348),
            .I(N__4345));
    LocalMux I__746 (
            .O(N__4345),
            .I(N__4342));
    IoSpan4Mux I__745 (
            .O(N__4342),
            .I(N__4339));
    IoSpan4Mux I__744 (
            .O(N__4339),
            .I(N__4336));
    Span4Mux_s0_v I__743 (
            .O(N__4336),
            .I(N__4333));
    Sp12to4 I__742 (
            .O(N__4333),
            .I(N__4329));
    CascadeMux I__741 (
            .O(N__4332),
            .I(N__4326));
    Span12Mux_s11_v I__740 (
            .O(N__4329),
            .I(N__4323));
    InMux I__739 (
            .O(N__4326),
            .I(N__4320));
    Odrv12 I__738 (
            .O(N__4323),
            .I(ROMENn_c));
    LocalMux I__737 (
            .O(N__4320),
            .I(ROMENn_c));
    InMux I__736 (
            .O(N__4315),
            .I(N__4308));
    InMux I__735 (
            .O(N__4314),
            .I(N__4305));
    InMux I__734 (
            .O(N__4313),
            .I(N__4298));
    InMux I__733 (
            .O(N__4312),
            .I(N__4298));
    InMux I__732 (
            .O(N__4311),
            .I(N__4298));
    LocalMux I__731 (
            .O(N__4308),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__730 (
            .O(N__4305),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__729 (
            .O(N__4298),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    InMux I__728 (
            .O(N__4291),
            .I(N__4283));
    InMux I__727 (
            .O(N__4290),
            .I(N__4280));
    InMux I__726 (
            .O(N__4289),
            .I(N__4271));
    InMux I__725 (
            .O(N__4288),
            .I(N__4271));
    InMux I__724 (
            .O(N__4287),
            .I(N__4271));
    InMux I__723 (
            .O(N__4286),
            .I(N__4271));
    LocalMux I__722 (
            .O(N__4283),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__721 (
            .O(N__4280),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__720 (
            .O(N__4271),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    InMux I__719 (
            .O(N__4264),
            .I(N__4261));
    LocalMux I__718 (
            .O(N__4261),
            .I(N__4258));
    Odrv12 I__717 (
            .O(N__4258),
            .I(\U409_TRANSFER_ACK.N_71 ));
    CascadeMux I__716 (
            .O(N__4255),
            .I(N__4252));
    InMux I__715 (
            .O(N__4252),
            .I(N__4249));
    LocalMux I__714 (
            .O(N__4249),
            .I(N__4246));
    Span4Mux_v I__713 (
            .O(N__4246),
            .I(N__4243));
    Span4Mux_h I__712 (
            .O(N__4243),
            .I(N__4240));
    Sp12to4 I__711 (
            .O(N__4240),
            .I(N__4237));
    Span12Mux_h I__710 (
            .O(N__4237),
            .I(N__4234));
    Span12Mux_v I__709 (
            .O(N__4234),
            .I(N__4231));
    Odrv12 I__708 (
            .O(N__4231),
            .I(TACKn_in));
    IoInMux I__707 (
            .O(N__4228),
            .I(N__4225));
    LocalMux I__706 (
            .O(N__4225),
            .I(N__4222));
    Span4Mux_s2_v I__705 (
            .O(N__4222),
            .I(N__4219));
    Span4Mux_h I__704 (
            .O(N__4219),
            .I(N__4216));
    Sp12to4 I__703 (
            .O(N__4216),
            .I(N__4213));
    Span12Mux_v I__702 (
            .O(N__4213),
            .I(N__4210));
    Odrv12 I__701 (
            .O(N__4210),
            .I(N_67_i));
    InMux I__700 (
            .O(N__4207),
            .I(N__4204));
    LocalMux I__699 (
            .O(N__4204),
            .I(N__4201));
    Span4Mux_v I__698 (
            .O(N__4201),
            .I(N__4196));
    InMux I__697 (
            .O(N__4200),
            .I(N__4193));
    InMux I__696 (
            .O(N__4199),
            .I(N__4190));
    Span4Mux_h I__695 (
            .O(N__4196),
            .I(N__4183));
    LocalMux I__694 (
            .O(N__4193),
            .I(N__4183));
    LocalMux I__693 (
            .O(N__4190),
            .I(N__4183));
    Odrv4 I__692 (
            .O(N__4183),
            .I(N_100));
    InMux I__691 (
            .O(N__4180),
            .I(N__4177));
    LocalMux I__690 (
            .O(N__4177),
            .I(N__4174));
    Span4Mux_h I__689 (
            .O(N__4174),
            .I(N__4169));
    InMux I__688 (
            .O(N__4173),
            .I(N__4164));
    InMux I__687 (
            .O(N__4172),
            .I(N__4164));
    Span4Mux_v I__686 (
            .O(N__4169),
            .I(N__4161));
    LocalMux I__685 (
            .O(N__4164),
            .I(N__4158));
    Sp12to4 I__684 (
            .O(N__4161),
            .I(N__4153));
    Span12Mux_v I__683 (
            .O(N__4158),
            .I(N__4153));
    Span12Mux_v I__682 (
            .O(N__4153),
            .I(N__4150));
    Span12Mux_h I__681 (
            .O(N__4150),
            .I(N__4147));
    Odrv12 I__680 (
            .O(N__4147),
            .I(OVL_c));
    InMux I__679 (
            .O(N__4144),
            .I(N__4141));
    LocalMux I__678 (
            .O(N__4141),
            .I(N__4138));
    Span4Mux_v I__677 (
            .O(N__4138),
            .I(N__4134));
    InMux I__676 (
            .O(N__4137),
            .I(N__4131));
    Odrv4 I__675 (
            .O(N__4134),
            .I(N_67));
    LocalMux I__674 (
            .O(N__4131),
            .I(N_67));
    CascadeMux I__673 (
            .O(N__4126),
            .I(N__4123));
    InMux I__672 (
            .O(N__4123),
            .I(N__4119));
    CascadeMux I__671 (
            .O(N__4122),
            .I(N__4116));
    LocalMux I__670 (
            .O(N__4119),
            .I(N__4113));
    InMux I__669 (
            .O(N__4116),
            .I(N__4110));
    Span4Mux_h I__668 (
            .O(N__4113),
            .I(N__4105));
    LocalMux I__667 (
            .O(N__4110),
            .I(N__4105));
    Span4Mux_v I__666 (
            .O(N__4105),
            .I(N__4102));
    Span4Mux_h I__665 (
            .O(N__4102),
            .I(N__4099));
    Odrv4 I__664 (
            .O(N__4099),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz ));
    InMux I__663 (
            .O(N__4096),
            .I(N__4092));
    InMux I__662 (
            .O(N__4095),
            .I(N__4089));
    LocalMux I__661 (
            .O(N__4092),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ));
    LocalMux I__660 (
            .O(N__4089),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ));
    InMux I__659 (
            .O(N__4084),
            .I(N__4081));
    LocalMux I__658 (
            .O(N__4081),
            .I(N__4078));
    Odrv4 I__657 (
            .O(N__4078),
            .I(\U409_TRANSFER_ACK.N_106 ));
    InMux I__656 (
            .O(N__4075),
            .I(N__4072));
    LocalMux I__655 (
            .O(N__4072),
            .I(N__4069));
    Span4Mux_h I__654 (
            .O(N__4069),
            .I(N__4066));
    Odrv4 I__653 (
            .O(N__4066),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER15Z0Z_1 ));
    InMux I__652 (
            .O(N__4063),
            .I(N__4058));
    InMux I__651 (
            .O(N__4062),
            .I(N__4052));
    InMux I__650 (
            .O(N__4061),
            .I(N__4052));
    LocalMux I__649 (
            .O(N__4058),
            .I(N__4049));
    InMux I__648 (
            .O(N__4057),
            .I(N__4046));
    LocalMux I__647 (
            .O(N__4052),
            .I(N__4043));
    Span4Mux_h I__646 (
            .O(N__4049),
            .I(N__4038));
    LocalMux I__645 (
            .O(N__4046),
            .I(N__4038));
    Odrv12 I__644 (
            .O(N__4043),
            .I(U409_ADDRESS_DECODE_Z2_SPACE));
    Odrv4 I__643 (
            .O(N__4038),
            .I(U409_ADDRESS_DECODE_Z2_SPACE));
    InMux I__642 (
            .O(N__4033),
            .I(N__4030));
    LocalMux I__641 (
            .O(N__4030),
            .I(N__4027));
    Odrv12 I__640 (
            .O(N__4027),
            .I(\U409_DATA_BUFFERS.un1_BUFENn_iZ0Z_0 ));
    CascadeMux I__639 (
            .O(N__4024),
            .I(N__4021));
    InMux I__638 (
            .O(N__4021),
            .I(N__4018));
    LocalMux I__637 (
            .O(N__4018),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_1 ));
    InMux I__636 (
            .O(N__4015),
            .I(N__4011));
    InMux I__635 (
            .O(N__4014),
            .I(N__4008));
    LocalMux I__634 (
            .O(N__4011),
            .I(N__4004));
    LocalMux I__633 (
            .O(N__4008),
            .I(N__4001));
    InMux I__632 (
            .O(N__4007),
            .I(N__3996));
    Span4Mux_v I__631 (
            .O(N__4004),
            .I(N__3991));
    Span4Mux_v I__630 (
            .O(N__4001),
            .I(N__3991));
    InMux I__629 (
            .O(N__4000),
            .I(N__3988));
    InMux I__628 (
            .O(N__3999),
            .I(N__3985));
    LocalMux I__627 (
            .O(N__3996),
            .I(N__3982));
    Sp12to4 I__626 (
            .O(N__3991),
            .I(N__3977));
    LocalMux I__625 (
            .O(N__3988),
            .I(N__3977));
    LocalMux I__624 (
            .O(N__3985),
            .I(N__3974));
    Span12Mux_v I__623 (
            .O(N__3982),
            .I(N__3971));
    Span12Mux_h I__622 (
            .O(N__3977),
            .I(N__3966));
    Span12Mux_v I__621 (
            .O(N__3974),
            .I(N__3966));
    Odrv12 I__620 (
            .O(N__3971),
            .I(A_c_20));
    Odrv12 I__619 (
            .O(N__3966),
            .I(A_c_20));
    CascadeMux I__618 (
            .O(N__3961),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4_cascade_ ));
    CascadeMux I__617 (
            .O(N__3958),
            .I(CIA_SPACE_cascade_));
    InMux I__616 (
            .O(N__3955),
            .I(N__3952));
    LocalMux I__615 (
            .O(N__3952),
            .I(\U409_ADDRESS_DECODE.N_69 ));
    IoInMux I__614 (
            .O(N__3949),
            .I(N__3946));
    LocalMux I__613 (
            .O(N__3946),
            .I(N__3943));
    IoSpan4Mux I__612 (
            .O(N__3943),
            .I(N__3940));
    Span4Mux_s2_v I__611 (
            .O(N__3940),
            .I(N__3937));
    Span4Mux_v I__610 (
            .O(N__3937),
            .I(N__3934));
    Span4Mux_v I__609 (
            .O(N__3934),
            .I(N__3931));
    Odrv4 I__608 (
            .O(N__3931),
            .I(PORTSIZE_0_i));
    CascadeMux I__607 (
            .O(N__3928),
            .I(\U409_ADDRESS_DECODE.un5_RAMSPACEn_cascade_ ));
    InMux I__606 (
            .O(N__3925),
            .I(N__3914));
    InMux I__605 (
            .O(N__3924),
            .I(N__3914));
    InMux I__604 (
            .O(N__3923),
            .I(N__3914));
    InMux I__603 (
            .O(N__3922),
            .I(N__3909));
    InMux I__602 (
            .O(N__3921),
            .I(N__3909));
    LocalMux I__601 (
            .O(N__3914),
            .I(N__3906));
    LocalMux I__600 (
            .O(N__3909),
            .I(N__3903));
    Span4Mux_v I__599 (
            .O(N__3906),
            .I(N__3899));
    Span4Mux_v I__598 (
            .O(N__3903),
            .I(N__3896));
    InMux I__597 (
            .O(N__3902),
            .I(N__3893));
    Sp12to4 I__596 (
            .O(N__3899),
            .I(N__3886));
    Sp12to4 I__595 (
            .O(N__3896),
            .I(N__3886));
    LocalMux I__594 (
            .O(N__3893),
            .I(N__3886));
    Odrv12 I__593 (
            .O(N__3886),
            .I(A_c_21));
    CascadeMux I__592 (
            .O(N__3883),
            .I(N__3879));
    CascadeMux I__591 (
            .O(N__3882),
            .I(N__3876));
    InMux I__590 (
            .O(N__3879),
            .I(N__3871));
    InMux I__589 (
            .O(N__3876),
            .I(N__3871));
    LocalMux I__588 (
            .O(N__3871),
            .I(N__3865));
    InMux I__587 (
            .O(N__3870),
            .I(N__3862));
    InMux I__586 (
            .O(N__3869),
            .I(N__3857));
    InMux I__585 (
            .O(N__3868),
            .I(N__3857));
    Span4Mux_v I__584 (
            .O(N__3865),
            .I(N__3854));
    LocalMux I__583 (
            .O(N__3862),
            .I(N__3849));
    LocalMux I__582 (
            .O(N__3857),
            .I(N__3849));
    Span4Mux_h I__581 (
            .O(N__3854),
            .I(N__3846));
    Span4Mux_v I__580 (
            .O(N__3849),
            .I(N__3843));
    Sp12to4 I__579 (
            .O(N__3846),
            .I(N__3838));
    Sp12to4 I__578 (
            .O(N__3843),
            .I(N__3838));
    Odrv12 I__577 (
            .O(N__3838),
            .I(A_c_23));
    InMux I__576 (
            .O(N__3835),
            .I(N__3824));
    InMux I__575 (
            .O(N__3834),
            .I(N__3824));
    InMux I__574 (
            .O(N__3833),
            .I(N__3824));
    InMux I__573 (
            .O(N__3832),
            .I(N__3819));
    InMux I__572 (
            .O(N__3831),
            .I(N__3819));
    LocalMux I__571 (
            .O(N__3824),
            .I(N__3814));
    LocalMux I__570 (
            .O(N__3819),
            .I(N__3814));
    Sp12to4 I__569 (
            .O(N__3814),
            .I(N__3811));
    Span12Mux_v I__568 (
            .O(N__3811),
            .I(N__3808));
    Odrv12 I__567 (
            .O(N__3808),
            .I(A_c_22));
    CascadeMux I__566 (
            .O(N__3805),
            .I(N__3799));
    InMux I__565 (
            .O(N__3804),
            .I(N__3792));
    InMux I__564 (
            .O(N__3803),
            .I(N__3792));
    InMux I__563 (
            .O(N__3802),
            .I(N__3792));
    InMux I__562 (
            .O(N__3799),
            .I(N__3789));
    LocalMux I__561 (
            .O(N__3792),
            .I(N__3784));
    LocalMux I__560 (
            .O(N__3789),
            .I(N__3784));
    Span12Mux_h I__559 (
            .O(N__3784),
            .I(N__3781));
    Span12Mux_v I__558 (
            .O(N__3781),
            .I(N__3778));
    Odrv12 I__557 (
            .O(N__3778),
            .I(TM_c_0));
    InMux I__556 (
            .O(N__3775),
            .I(N__3772));
    LocalMux I__555 (
            .O(N__3772),
            .I(U409_ADDRESS_DECODE_HIROM));
    CascadeMux I__554 (
            .O(N__3769),
            .I(U409_ADDRESS_DECODE_LOWROM_cascade_));
    InMux I__553 (
            .O(N__3766),
            .I(N__3756));
    InMux I__552 (
            .O(N__3765),
            .I(N__3756));
    InMux I__551 (
            .O(N__3764),
            .I(N__3756));
    InMux I__550 (
            .O(N__3763),
            .I(N__3753));
    LocalMux I__549 (
            .O(N__3756),
            .I(N__3748));
    LocalMux I__548 (
            .O(N__3753),
            .I(N__3748));
    Span4Mux_h I__547 (
            .O(N__3748),
            .I(N__3745));
    Sp12to4 I__546 (
            .O(N__3745),
            .I(N__3742));
    Odrv12 I__545 (
            .O(N__3742),
            .I(TM_c_1));
    InMux I__544 (
            .O(N__3739),
            .I(N__3735));
    InMux I__543 (
            .O(N__3738),
            .I(N__3731));
    LocalMux I__542 (
            .O(N__3735),
            .I(N__3725));
    InMux I__541 (
            .O(N__3734),
            .I(N__3722));
    LocalMux I__540 (
            .O(N__3731),
            .I(N__3719));
    InMux I__539 (
            .O(N__3730),
            .I(N__3716));
    InMux I__538 (
            .O(N__3729),
            .I(N__3713));
    InMux I__537 (
            .O(N__3728),
            .I(N__3710));
    Odrv12 I__536 (
            .O(N__3725),
            .I(N_107));
    LocalMux I__535 (
            .O(N__3722),
            .I(N_107));
    Odrv4 I__534 (
            .O(N__3719),
            .I(N_107));
    LocalMux I__533 (
            .O(N__3716),
            .I(N_107));
    LocalMux I__532 (
            .O(N__3713),
            .I(N_107));
    LocalMux I__531 (
            .O(N__3710),
            .I(N_107));
    InMux I__530 (
            .O(N__3697),
            .I(N__3693));
    InMux I__529 (
            .O(N__3696),
            .I(N__3689));
    LocalMux I__528 (
            .O(N__3693),
            .I(N__3686));
    InMux I__527 (
            .O(N__3692),
            .I(N__3683));
    LocalMux I__526 (
            .O(N__3689),
            .I(N__3680));
    Odrv4 I__525 (
            .O(N__3686),
            .I(N_33));
    LocalMux I__524 (
            .O(N__3683),
            .I(N_33));
    Odrv4 I__523 (
            .O(N__3680),
            .I(N_33));
    IoInMux I__522 (
            .O(N__3673),
            .I(N__3670));
    LocalMux I__521 (
            .O(N__3670),
            .I(N__3667));
    IoSpan4Mux I__520 (
            .O(N__3667),
            .I(N__3664));
    IoSpan4Mux I__519 (
            .O(N__3664),
            .I(N__3661));
    Sp12to4 I__518 (
            .O(N__3661),
            .I(N__3658));
    Span12Mux_v I__517 (
            .O(N__3658),
            .I(N__3655));
    Odrv12 I__516 (
            .O(N__3655),
            .I(N_68_i));
    CascadeMux I__515 (
            .O(N__3652),
            .I(N_74_1_cascade_));
    CascadeMux I__514 (
            .O(N__3649),
            .I(N_33_cascade_));
    InMux I__513 (
            .O(N__3646),
            .I(N__3643));
    LocalMux I__512 (
            .O(N__3643),
            .I(N_99));
    InMux I__511 (
            .O(N__3640),
            .I(N__3636));
    InMux I__510 (
            .O(N__3639),
            .I(N__3633));
    LocalMux I__509 (
            .O(N__3636),
            .I(N__3628));
    LocalMux I__508 (
            .O(N__3633),
            .I(N__3628));
    Span4Mux_v I__507 (
            .O(N__3628),
            .I(N__3624));
    InMux I__506 (
            .O(N__3627),
            .I(N__3621));
    Odrv4 I__505 (
            .O(N__3624),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_a2_5));
    LocalMux I__504 (
            .O(N__3621),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_a2_5));
    CascadeMux I__503 (
            .O(N__3616),
            .I(N_99_cascade_));
    InMux I__502 (
            .O(N__3613),
            .I(N__3610));
    LocalMux I__501 (
            .O(N__3610),
            .I(N__3605));
    InMux I__500 (
            .O(N__3609),
            .I(N__3602));
    InMux I__499 (
            .O(N__3608),
            .I(N__3599));
    Span4Mux_v I__498 (
            .O(N__3605),
            .I(N__3594));
    LocalMux I__497 (
            .O(N__3602),
            .I(N__3594));
    LocalMux I__496 (
            .O(N__3599),
            .I(N__3591));
    Span4Mux_h I__495 (
            .O(N__3594),
            .I(N__3588));
    Span4Mux_v I__494 (
            .O(N__3591),
            .I(N__3585));
    Odrv4 I__493 (
            .O(N__3588),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_a2_4));
    Odrv4 I__492 (
            .O(N__3585),
            .I(U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_a2_4));
    InMux I__491 (
            .O(N__3580),
            .I(N__3574));
    InMux I__490 (
            .O(N__3579),
            .I(N__3571));
    InMux I__489 (
            .O(N__3578),
            .I(N__3568));
    InMux I__488 (
            .O(N__3577),
            .I(N__3565));
    LocalMux I__487 (
            .O(N__3574),
            .I(N__3558));
    LocalMux I__486 (
            .O(N__3571),
            .I(N__3558));
    LocalMux I__485 (
            .O(N__3568),
            .I(N__3558));
    LocalMux I__484 (
            .O(N__3565),
            .I(N__3555));
    Span4Mux_v I__483 (
            .O(N__3558),
            .I(N__3552));
    Span4Mux_v I__482 (
            .O(N__3555),
            .I(N__3549));
    Sp12to4 I__481 (
            .O(N__3552),
            .I(N__3544));
    Sp12to4 I__480 (
            .O(N__3549),
            .I(N__3544));
    Span12Mux_h I__479 (
            .O(N__3544),
            .I(N__3541));
    Span12Mux_v I__478 (
            .O(N__3541),
            .I(N__3538));
    Odrv12 I__477 (
            .O(N__3538),
            .I(A_c_18));
    InMux I__476 (
            .O(N__3535),
            .I(N__3532));
    LocalMux I__475 (
            .O(N__3532),
            .I(N__3528));
    CascadeMux I__474 (
            .O(N__3531),
            .I(N__3525));
    Span4Mux_v I__473 (
            .O(N__3528),
            .I(N__3522));
    InMux I__472 (
            .O(N__3525),
            .I(N__3519));
    Odrv4 I__471 (
            .O(N__3522),
            .I(N_74_1));
    LocalMux I__470 (
            .O(N__3519),
            .I(N_74_1));
    InMux I__469 (
            .O(N__3514),
            .I(N__3509));
    InMux I__468 (
            .O(N__3513),
            .I(N__3506));
    CascadeMux I__467 (
            .O(N__3512),
            .I(N__3503));
    LocalMux I__466 (
            .O(N__3509),
            .I(N__3500));
    LocalMux I__465 (
            .O(N__3506),
            .I(N__3497));
    InMux I__464 (
            .O(N__3503),
            .I(N__3494));
    Odrv4 I__463 (
            .O(N__3500),
            .I(N_101));
    Odrv4 I__462 (
            .O(N__3497),
            .I(N_101));
    LocalMux I__461 (
            .O(N__3494),
            .I(N_101));
    InMux I__460 (
            .O(N__3487),
            .I(N__3484));
    LocalMux I__459 (
            .O(N__3484),
            .I(N__3481));
    Span12Mux_h I__458 (
            .O(N__3481),
            .I(N__3478));
    Span12Mux_v I__457 (
            .O(N__3478),
            .I(N__3475));
    Odrv12 I__456 (
            .O(N__3475),
            .I(TT_c_0));
    InMux I__455 (
            .O(N__3472),
            .I(N__3469));
    LocalMux I__454 (
            .O(N__3469),
            .I(N__3466));
    Span4Mux_h I__453 (
            .O(N__3466),
            .I(N__3463));
    Odrv4 I__452 (
            .O(N__3463),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_9 ));
    InMux I__451 (
            .O(N__3460),
            .I(N__3452));
    InMux I__450 (
            .O(N__3459),
            .I(N__3452));
    InMux I__449 (
            .O(N__3458),
            .I(N__3449));
    InMux I__448 (
            .O(N__3457),
            .I(N__3446));
    LocalMux I__447 (
            .O(N__3452),
            .I(N__3440));
    LocalMux I__446 (
            .O(N__3449),
            .I(N__3440));
    LocalMux I__445 (
            .O(N__3446),
            .I(N__3437));
    InMux I__444 (
            .O(N__3445),
            .I(N__3434));
    Span4Mux_v I__443 (
            .O(N__3440),
            .I(N__3431));
    Span4Mux_h I__442 (
            .O(N__3437),
            .I(N__3428));
    LocalMux I__441 (
            .O(N__3434),
            .I(N__3425));
    Sp12to4 I__440 (
            .O(N__3431),
            .I(N__3422));
    Span4Mux_h I__439 (
            .O(N__3428),
            .I(N__3419));
    Span4Mux_h I__438 (
            .O(N__3425),
            .I(N__3416));
    Span12Mux_h I__437 (
            .O(N__3422),
            .I(N__3409));
    Sp12to4 I__436 (
            .O(N__3419),
            .I(N__3409));
    Sp12to4 I__435 (
            .O(N__3416),
            .I(N__3409));
    Span12Mux_v I__434 (
            .O(N__3409),
            .I(N__3406));
    Odrv12 I__433 (
            .O(N__3406),
            .I(A_c_19));
    CascadeMux I__432 (
            .O(N__3403),
            .I(\U409_ADDRESS_DECODE.HIROMZ0Z_1_cascade_ ));
    InMux I__431 (
            .O(N__3400),
            .I(N__3394));
    InMux I__430 (
            .O(N__3399),
            .I(N__3394));
    LocalMux I__429 (
            .O(N__3394),
            .I(\U409_TRANSFER_ACK.N_94 ));
    InMux I__428 (
            .O(N__3391),
            .I(N__3387));
    InMux I__427 (
            .O(N__3390),
            .I(N__3383));
    LocalMux I__426 (
            .O(N__3387),
            .I(N__3380));
    InMux I__425 (
            .O(N__3386),
            .I(N__3377));
    LocalMux I__424 (
            .O(N__3383),
            .I(N__3374));
    Span4Mux_v I__423 (
            .O(N__3380),
            .I(N__3371));
    LocalMux I__422 (
            .O(N__3377),
            .I(N__3368));
    Span4Mux_v I__421 (
            .O(N__3374),
            .I(N__3365));
    Sp12to4 I__420 (
            .O(N__3371),
            .I(N__3360));
    Span12Mux_v I__419 (
            .O(N__3368),
            .I(N__3360));
    Span4Mux_h I__418 (
            .O(N__3365),
            .I(N__3357));
    Odrv12 I__417 (
            .O(N__3360),
            .I(A_c_27));
    Odrv4 I__416 (
            .O(N__3357),
            .I(A_c_27));
    InMux I__415 (
            .O(N__3352),
            .I(N__3346));
    InMux I__414 (
            .O(N__3351),
            .I(N__3346));
    LocalMux I__413 (
            .O(N__3346),
            .I(N__3342));
    InMux I__412 (
            .O(N__3345),
            .I(N__3339));
    Span4Mux_h I__411 (
            .O(N__3342),
            .I(N__3334));
    LocalMux I__410 (
            .O(N__3339),
            .I(N__3334));
    Span4Mux_h I__409 (
            .O(N__3334),
            .I(N__3331));
    Span4Mux_v I__408 (
            .O(N__3331),
            .I(N__3328));
    Span4Mux_v I__407 (
            .O(N__3328),
            .I(N__3325));
    Odrv4 I__406 (
            .O(N__3325),
            .I(A_c_26));
    CascadeMux I__405 (
            .O(N__3322),
            .I(N__3317));
    CascadeMux I__404 (
            .O(N__3321),
            .I(N__3314));
    InMux I__403 (
            .O(N__3320),
            .I(N__3311));
    InMux I__402 (
            .O(N__3317),
            .I(N__3306));
    InMux I__401 (
            .O(N__3314),
            .I(N__3306));
    LocalMux I__400 (
            .O(N__3311),
            .I(N__3303));
    LocalMux I__399 (
            .O(N__3306),
            .I(N__3300));
    Span4Mux_v I__398 (
            .O(N__3303),
            .I(N__3297));
    Sp12to4 I__397 (
            .O(N__3300),
            .I(N__3294));
    Span4Mux_v I__396 (
            .O(N__3297),
            .I(N__3291));
    Span12Mux_v I__395 (
            .O(N__3294),
            .I(N__3288));
    Span4Mux_h I__394 (
            .O(N__3291),
            .I(N__3285));
    Odrv12 I__393 (
            .O(N__3288),
            .I(A_c_24));
    Odrv4 I__392 (
            .O(N__3285),
            .I(A_c_24));
    CascadeMux I__391 (
            .O(N__3280),
            .I(N__3275));
    InMux I__390 (
            .O(N__3279),
            .I(N__3270));
    InMux I__389 (
            .O(N__3278),
            .I(N__3270));
    InMux I__388 (
            .O(N__3275),
            .I(N__3267));
    LocalMux I__387 (
            .O(N__3270),
            .I(N__3264));
    LocalMux I__386 (
            .O(N__3267),
            .I(N__3261));
    Span4Mux_v I__385 (
            .O(N__3264),
            .I(N__3258));
    Span4Mux_v I__384 (
            .O(N__3261),
            .I(N__3255));
    Sp12to4 I__383 (
            .O(N__3258),
            .I(N__3252));
    Span4Mux_h I__382 (
            .O(N__3255),
            .I(N__3249));
    Odrv12 I__381 (
            .O(N__3252),
            .I(A_c_25));
    Odrv4 I__380 (
            .O(N__3249),
            .I(A_c_25));
    InMux I__379 (
            .O(N__3244),
            .I(N__3241));
    LocalMux I__378 (
            .O(N__3241),
            .I(N__3238));
    Odrv4 I__377 (
            .O(N__3238),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_7 ));
    CascadeMux I__376 (
            .O(N__3235),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_8_cascade_ ));
    InMux I__375 (
            .O(N__3232),
            .I(N__3229));
    LocalMux I__374 (
            .O(N__3229),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_10 ));
    IoInMux I__373 (
            .O(N__3226),
            .I(N__3223));
    LocalMux I__372 (
            .O(N__3223),
            .I(N__3220));
    IoSpan4Mux I__371 (
            .O(N__3220),
            .I(N__3217));
    Span4Mux_s3_h I__370 (
            .O(N__3217),
            .I(N__3214));
    Sp12to4 I__369 (
            .O(N__3214),
            .I(N__3211));
    Span12Mux_v I__368 (
            .O(N__3211),
            .I(N__3208));
    Span12Mux_h I__367 (
            .O(N__3208),
            .I(N__3205));
    Odrv12 I__366 (
            .O(N__3205),
            .I(N_69_i));
    InMux I__365 (
            .O(N__3202),
            .I(N__3199));
    LocalMux I__364 (
            .O(N__3199),
            .I(N__3196));
    Span4Mux_v I__363 (
            .O(N__3196),
            .I(N__3193));
    Odrv4 I__362 (
            .O(N__3193),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_13 ));
    CascadeMux I__361 (
            .O(N__3190),
            .I(N_101_cascade_));
    InMux I__360 (
            .O(N__3187),
            .I(N__3183));
    InMux I__359 (
            .O(N__3186),
            .I(N__3180));
    LocalMux I__358 (
            .O(N__3183),
            .I(N__3177));
    LocalMux I__357 (
            .O(N__3180),
            .I(N__3174));
    Odrv12 I__356 (
            .O(N__3177),
            .I(N_105));
    Odrv4 I__355 (
            .O(N__3174),
            .I(N_105));
    CascadeMux I__354 (
            .O(N__3169),
            .I(N__3166));
    InMux I__353 (
            .O(N__3166),
            .I(N__3161));
    InMux I__352 (
            .O(N__3165),
            .I(N__3156));
    InMux I__351 (
            .O(N__3164),
            .I(N__3156));
    LocalMux I__350 (
            .O(N__3161),
            .I(N__3153));
    LocalMux I__349 (
            .O(N__3156),
            .I(N__3150));
    Span4Mux_h I__348 (
            .O(N__3153),
            .I(N__3146));
    Span4Mux_v I__347 (
            .O(N__3150),
            .I(N__3143));
    InMux I__346 (
            .O(N__3149),
            .I(N__3140));
    Span4Mux_h I__345 (
            .O(N__3146),
            .I(N__3137));
    Sp12to4 I__344 (
            .O(N__3143),
            .I(N__3132));
    LocalMux I__343 (
            .O(N__3140),
            .I(N__3132));
    Sp12to4 I__342 (
            .O(N__3137),
            .I(N__3127));
    Span12Mux_h I__341 (
            .O(N__3132),
            .I(N__3127));
    Span12Mux_v I__340 (
            .O(N__3127),
            .I(N__3124));
    Odrv12 I__339 (
            .O(N__3124),
            .I(A_c_16));
    InMux I__338 (
            .O(N__3121),
            .I(N__3115));
    InMux I__337 (
            .O(N__3120),
            .I(N__3115));
    LocalMux I__336 (
            .O(N__3115),
            .I(N__3110));
    InMux I__335 (
            .O(N__3114),
            .I(N__3107));
    InMux I__334 (
            .O(N__3113),
            .I(N__3104));
    Span4Mux_h I__333 (
            .O(N__3110),
            .I(N__3099));
    LocalMux I__332 (
            .O(N__3107),
            .I(N__3099));
    LocalMux I__331 (
            .O(N__3104),
            .I(N__3096));
    Span4Mux_v I__330 (
            .O(N__3099),
            .I(N__3093));
    Sp12to4 I__329 (
            .O(N__3096),
            .I(N__3090));
    Sp12to4 I__328 (
            .O(N__3093),
            .I(N__3087));
    Span12Mux_v I__327 (
            .O(N__3090),
            .I(N__3084));
    Span12Mux_v I__326 (
            .O(N__3087),
            .I(N__3081));
    Odrv12 I__325 (
            .O(N__3084),
            .I(A_c_17));
    Odrv12 I__324 (
            .O(N__3081),
            .I(A_c_17));
    CascadeMux I__323 (
            .O(N__3076),
            .I(N__3071));
    CascadeMux I__322 (
            .O(N__3075),
            .I(N__3068));
    InMux I__321 (
            .O(N__3074),
            .I(N__3061));
    InMux I__320 (
            .O(N__3071),
            .I(N__3061));
    InMux I__319 (
            .O(N__3068),
            .I(N__3061));
    LocalMux I__318 (
            .O(N__3061),
            .I(N__3058));
    Span4Mux_h I__317 (
            .O(N__3058),
            .I(N__3055));
    Sp12to4 I__316 (
            .O(N__3055),
            .I(N__3052));
    Span12Mux_v I__315 (
            .O(N__3052),
            .I(N__3049));
    Odrv12 I__314 (
            .O(N__3049),
            .I(A_c_28));
    CascadeMux I__313 (
            .O(N__3046),
            .I(\U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_7_cascade_ ));
    CascadeMux I__312 (
            .O(N__3043),
            .I(N__3040));
    InMux I__311 (
            .O(N__3040),
            .I(N__3031));
    InMux I__310 (
            .O(N__3039),
            .I(N__3031));
    InMux I__309 (
            .O(N__3038),
            .I(N__3031));
    LocalMux I__308 (
            .O(N__3031),
            .I(N__3028));
    Sp12to4 I__307 (
            .O(N__3028),
            .I(N__3025));
    Span12Mux_v I__306 (
            .O(N__3025),
            .I(N__3022));
    Odrv12 I__305 (
            .O(N__3022),
            .I(A_c_29));
    InMux I__304 (
            .O(N__3019),
            .I(N__3016));
    LocalMux I__303 (
            .O(N__3016),
            .I(\U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_8 ));
    CascadeMux I__302 (
            .O(N__3013),
            .I(\U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_9_cascade_ ));
    InMux I__301 (
            .O(N__3010),
            .I(N__3007));
    LocalMux I__300 (
            .O(N__3007),
            .I(\U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_10 ));
    IoInMux I__299 (
            .O(N__3004),
            .I(N__3001));
    LocalMux I__298 (
            .O(N__3001),
            .I(N__2998));
    Span4Mux_s3_v I__297 (
            .O(N__2998),
            .I(N__2995));
    Sp12to4 I__296 (
            .O(N__2995),
            .I(N__2992));
    Span12Mux_h I__295 (
            .O(N__2992),
            .I(N__2989));
    Span12Mux_h I__294 (
            .O(N__2989),
            .I(N__2986));
    Odrv12 I__293 (
            .O(N__2986),
            .I(N_31_i));
    InMux I__292 (
            .O(N__2983),
            .I(N__2978));
    InMux I__291 (
            .O(N__2982),
            .I(N__2973));
    InMux I__290 (
            .O(N__2981),
            .I(N__2973));
    LocalMux I__289 (
            .O(N__2978),
            .I(N__2970));
    LocalMux I__288 (
            .O(N__2973),
            .I(N__2967));
    Span4Mux_v I__287 (
            .O(N__2970),
            .I(N__2964));
    Span4Mux_v I__286 (
            .O(N__2967),
            .I(N__2961));
    Span4Mux_v I__285 (
            .O(N__2964),
            .I(N__2958));
    Span4Mux_v I__284 (
            .O(N__2961),
            .I(N__2955));
    Span4Mux_h I__283 (
            .O(N__2958),
            .I(N__2952));
    Span4Mux_h I__282 (
            .O(N__2955),
            .I(N__2949));
    Odrv4 I__281 (
            .O(N__2952),
            .I(A_c_31));
    Odrv4 I__280 (
            .O(N__2949),
            .I(A_c_31));
    CascadeMux I__279 (
            .O(N__2944),
            .I(N__2941));
    InMux I__278 (
            .O(N__2941),
            .I(N__2938));
    LocalMux I__277 (
            .O(N__2938),
            .I(N__2935));
    Span12Mux_v I__276 (
            .O(N__2935),
            .I(N__2932));
    Odrv12 I__275 (
            .O(N__2932),
            .I(TT_c_1));
    CascadeMux I__274 (
            .O(N__2929),
            .I(N__2924));
    InMux I__273 (
            .O(N__2928),
            .I(N__2921));
    InMux I__272 (
            .O(N__2927),
            .I(N__2918));
    InMux I__271 (
            .O(N__2924),
            .I(N__2915));
    LocalMux I__270 (
            .O(N__2921),
            .I(N__2910));
    LocalMux I__269 (
            .O(N__2918),
            .I(N__2910));
    LocalMux I__268 (
            .O(N__2915),
            .I(N__2905));
    Sp12to4 I__267 (
            .O(N__2910),
            .I(N__2905));
    Span12Mux_v I__266 (
            .O(N__2905),
            .I(N__2902));
    Odrv12 I__265 (
            .O(N__2902),
            .I(A_c_30));
    ClkMux I__264 (
            .O(N__2899),
            .I(N__2857));
    ClkMux I__263 (
            .O(N__2898),
            .I(N__2857));
    ClkMux I__262 (
            .O(N__2897),
            .I(N__2857));
    ClkMux I__261 (
            .O(N__2896),
            .I(N__2857));
    ClkMux I__260 (
            .O(N__2895),
            .I(N__2857));
    ClkMux I__259 (
            .O(N__2894),
            .I(N__2857));
    ClkMux I__258 (
            .O(N__2893),
            .I(N__2857));
    ClkMux I__257 (
            .O(N__2892),
            .I(N__2857));
    ClkMux I__256 (
            .O(N__2891),
            .I(N__2857));
    ClkMux I__255 (
            .O(N__2890),
            .I(N__2857));
    ClkMux I__254 (
            .O(N__2889),
            .I(N__2857));
    ClkMux I__253 (
            .O(N__2888),
            .I(N__2857));
    ClkMux I__252 (
            .O(N__2887),
            .I(N__2857));
    ClkMux I__251 (
            .O(N__2886),
            .I(N__2857));
    GlobalMux I__250 (
            .O(N__2857),
            .I(CLK80_OUT));
    INV \INVU409_TRANSFER_ACK.LASTCLK_0C  (
            .O(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .I(N__2892));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .I(N__2897));
    INV \INVU409_TRANSFER_ACK.CIA_ENABLED_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .I(N__2890));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_1C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .I(N__2888));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net ),
            .I(N__2886));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net ),
            .I(N__2899));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ),
            .I(N__2898));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ),
            .I(N__2896));
    INV \INVU409_TRANSFER_ACK.TACK_EN_iC  (
            .O(\INVU409_TRANSFER_ACK.TACK_EN_iC_net ),
            .I(N__2894));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .I(N__2891));
    INV \INVU409_TRANSFER_ACK.CIA_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .I(N__2889));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net ),
            .I(N__2887));
    INV \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC  (
            .O(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .I(N__2895));
    INV \INVU409_TRANSFER_ACK.IRQ_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net ),
            .I(N__2893));
    defparam IN_MUX_bfv_14_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_8_0_));
    defparam IN_MUX_bfv_14_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_9_0_ (
            .carryinitin(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .carryinitout(bfn_14_9_0_));
    defparam IN_MUX_bfv_15_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_3_0_));
    defparam IN_MUX_bfv_15_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_4_0_ (
            .carryinitin(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .carryinitout(bfn_15_4_0_));
    defparam IN_MUX_bfv_15_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_6_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_0_LC_1_11_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_0_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_0_LC_1_11_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_0_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__3149),
            .in2(_gnd_net_),
            .in3(N__3114),
            .lcout(N_105),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_7_LC_1_14_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_7_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_7_LC_1_14_0 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_7_LC_1_14_0  (
            .in0(N__3074),
            .in1(_gnd_net_),
            .in2(N__3043),
            .in3(N__3390),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_a2_4_LC_1_14_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_a2_4_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_a2_4_LC_1_14_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_a2_4_LC_1_14_4  (
            .in0(N__3039),
            .in1(N__2982),
            .in2(N__3076),
            .in3(N__2927),
            .lcout(U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_a2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_a4_7_LC_1_14_6 .C_ON=1'b0;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_a4_7_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_a4_7_LC_1_14_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_DATA_BUFFERS.un1_BUFENn_i_a4_7_LC_1_14_6  (
            .in0(N__3186),
            .in1(N__4207),
            .in2(N__3075),
            .in3(N__2981),
            .lcout(),
            .ltout(\U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_a4_10_LC_1_14_7 .C_ON=1'b0;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_a4_10_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_a4_10_LC_1_14_7 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U409_DATA_BUFFERS.un1_BUFENn_i_a4_10_LC_1_14_7  (
            .in0(N__3345),
            .in1(_gnd_net_),
            .in2(N__3046),
            .in3(N__3038),
            .lcout(\U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_a4_8_LC_2_13_1 .C_ON=1'b0;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_a4_8_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_a4_8_LC_2_13_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_DATA_BUFFERS.un1_BUFENn_i_a4_8_LC_2_13_1  (
            .in0(N__3445),
            .in1(N__3577),
            .in2(N__2929),
            .in3(N__5340),
            .lcout(\U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_a4_9_LC_2_14_0 .C_ON=1'b0;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_a4_9_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_a4_9_LC_2_14_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_DATA_BUFFERS.un1_BUFENn_i_a4_9_LC_2_14_0  (
            .in0(N__3999),
            .in1(N__3386),
            .in2(N__3280),
            .in3(N__3320),
            .lcout(),
            .ltout(\U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_DATA_BUFFERS.N_31_i_LC_2_14_1 .C_ON=1'b0;
    defparam \U409_DATA_BUFFERS.N_31_i_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \U409_DATA_BUFFERS.N_31_i_LC_2_14_1 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \U409_DATA_BUFFERS.N_31_i_LC_2_14_1  (
            .in0(N__4033),
            .in1(N__3019),
            .in2(N__3013),
            .in3(N__3010),
            .lcout(N_31_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_10_LC_2_14_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_10_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_10_LC_2_14_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_10_LC_2_14_4  (
            .in0(N__2983),
            .in1(N__3902),
            .in2(N__2944),
            .in3(N__2928),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_3_13_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_3_13_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_3_13_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_3_13_2  (
            .in0(N__3608),
            .in1(N__3627),
            .in2(_gnd_net_),
            .in3(N__5339),
            .lcout(U409_ADDRESS_DECODE_Z2_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_a2_5_LC_3_14_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_a2_5_LC_3_14_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_a2_5_LC_3_14_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_a2_5_LC_3_14_0  (
            .in0(N__3391),
            .in1(N__3351),
            .in2(N__3321),
            .in3(N__3278),
            .lcout(U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_a2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_8_LC_3_14_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_8_LC_3_14_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_8_LC_3_14_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_8_LC_3_14_4  (
            .in0(N__3535),
            .in1(N__3352),
            .in2(N__3322),
            .in3(N__3279),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_LC_3_14_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_LC_3_14_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_LC_3_14_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_LC_3_14_5  (
            .in0(N__3244),
            .in1(N__3472),
            .in2(N__3235),
            .in3(N__3232),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.N_69_i_LC_5_9_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.N_69_i_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.N_69_i_LC_5_9_0 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \U409_ADDRESS_DECODE.N_69_i_LC_5_9_0  (
            .in0(N__3513),
            .in1(N__3113),
            .in2(N__3169),
            .in3(N__3739),
            .lcout(N_69_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_LC_5_11_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_LC_5_11_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_LC_5_11_1  (
            .in0(N__3457),
            .in1(N__4015),
            .in2(_gnd_net_),
            .in3(N__3578),
            .lcout(N_101),
            .ltout(N_101_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_tz_tz_LC_5_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_tz_tz_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_tz_tz_LC_5_11_2 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_tz_tz_LC_5_11_2  (
            .in0(N__3738),
            .in1(N__3202),
            .in2(N__3190),
            .in3(N__3187),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a4_LC_5_12_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a4_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a4_LC_5_12_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a4_LC_5_12_2  (
            .in0(N__3120),
            .in1(N__3729),
            .in2(N__3512),
            .in3(N__3164),
            .lcout(\U409_ADDRESS_DECODE.N_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_1_LC_5_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_1_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_1_LC_5_12_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_1_LC_5_12_3  (
            .in0(N__3165),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3121),
            .lcout(N_74_1),
            .ltout(N_74_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_o2_LC_5_12_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_o2_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_o2_LC_5_12_4 .LUT_INIT=16'b1011001100110011;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_o2_LC_5_12_4  (
            .in0(N__3458),
            .in1(N__4000),
            .in2(N__3652),
            .in3(N__3579),
            .lcout(N_33),
            .ltout(N_33_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_a4_LC_5_12_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_a4_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_a4_LC_5_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_a4_LC_5_12_5  (
            .in0(N__3646),
            .in1(N__3640),
            .in2(N__3649),
            .in3(N__3613),
            .lcout(\U409_TRANSFER_ACK.N_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_a2_0_LC_5_13_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_a2_0_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_a2_0_LC_5_13_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_a2_0_LC_5_13_0  (
            .in0(N__3922),
            .in1(N__3399),
            .in2(N__3805),
            .in3(N__3763),
            .lcout(N_99),
            .ltout(N_99_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_LC_5_13_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_LC_5_13_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_LC_5_13_1  (
            .in0(N__3639),
            .in1(N__5335),
            .in2(N__3616),
            .in3(N__3609),
            .lcout(N_107),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_1_LC_5_13_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_1_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_1_LC_5_13_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_1_LC_5_13_2  (
            .in0(N__3580),
            .in1(N__3459),
            .in2(N__3531),
            .in3(N__3868),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_9_LC_5_13_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_9_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_9_LC_5_13_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_9_LC_5_13_3  (
            .in0(N__3400),
            .in1(N__3514),
            .in2(N__5341),
            .in3(N__3487),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.HIROM_1_LC_5_13_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.HIROM_1_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.HIROM_1_LC_5_13_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_ADDRESS_DECODE.HIROM_1_LC_5_13_4  (
            .in0(N__3831),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4014),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.HIROMZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.HIROM_LC_5_13_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.HIROM_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.HIROM_LC_5_13_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.HIROM_LC_5_13_5  (
            .in0(N__3460),
            .in1(N__3870),
            .in2(N__3403),
            .in3(N__3921),
            .lcout(U409_ADDRESS_DECODE_HIROM),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_LC_5_13_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_LC_5_13_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_LC_5_13_6  (
            .in0(N__3832),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3869),
            .lcout(\U409_TRANSFER_ACK.N_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_0_LC_5_14_7 .C_ON=1'b0;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_0_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_i_0_LC_5_14_7 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \U409_DATA_BUFFERS.un1_BUFENn_i_0_LC_5_14_7  (
            .in0(N__3730),
            .in1(N__3696),
            .in2(_gnd_net_),
            .in3(N__4144),
            .lcout(\U409_DATA_BUFFERS.un1_BUFENn_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_6_13_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_6_13_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_6_13_0  (
            .in0(N__3802),
            .in1(N__3923),
            .in2(N__4024),
            .in3(N__3764),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_6_13_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_6_13_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_LC_6_13_1  (
            .in0(N__4057),
            .in1(N__4007),
            .in2(N__3961),
            .in3(N__3833),
            .lcout(CIA_SPACE),
            .ltout(CIA_SPACE_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_6_13_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_6_13_2 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_6_13_2  (
            .in0(N__3692),
            .in1(N__3728),
            .in2(N__3958),
            .in3(N__3955),
            .lcout(PORTSIZE_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un5_RAMSPACEn_0_a2_LC_6_13_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un5_RAMSPACEn_0_a2_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un5_RAMSPACEn_0_a2_LC_6_13_3 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \U409_ADDRESS_DECODE.un5_RAMSPACEn_0_a2_LC_6_13_3  (
            .in0(N__3925),
            .in1(_gnd_net_),
            .in2(N__3883),
            .in3(N__3835),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.un5_RAMSPACEn_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a2_LC_6_13_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a2_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a2_LC_6_13_4 .LUT_INIT=16'b0101000010100000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a2_LC_6_13_4  (
            .in0(N__3803),
            .in1(_gnd_net_),
            .in2(N__3928),
            .in3(N__3765),
            .lcout(N_100),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.LOWROM_LC_6_13_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.LOWROM_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.LOWROM_LC_6_13_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U409_ADDRESS_DECODE.LOWROM_LC_6_13_5  (
            .in0(N__3924),
            .in1(N__4180),
            .in2(N__3882),
            .in3(N__3834),
            .lcout(),
            .ltout(U409_ADDRESS_DECODE_LOWROM_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_1_LC_6_13_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_1_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_1_LC_6_13_6 .LUT_INIT=16'b0101010010101000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_1_LC_6_13_6  (
            .in0(N__3804),
            .in1(N__3775),
            .in2(N__3769),
            .in3(N__3766),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER15Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.N_68_i_LC_6_14_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.N_68_i_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.N_68_i_LC_6_14_5 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U409_ADDRESS_DECODE.N_68_i_LC_6_14_5  (
            .in0(N__3734),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3697),
            .lcout(N_68_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_8_12_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_8_12_0 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_8_12_0  (
            .in0(N__4137),
            .in1(N__4264),
            .in2(N__4255),
            .in3(N__5328),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.N_67_i_LC_8_13_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.N_67_i_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.N_67_i_LC_8_13_0 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \U409_ADDRESS_DECODE.N_67_i_LC_8_13_0  (
            .in0(N__4172),
            .in1(N__4061),
            .in2(_gnd_net_),
            .in3(N__4199),
            .lcout(N_67_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a4_LC_8_13_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a4_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a4_LC_8_13_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a4_LC_8_13_3  (
            .in0(N__4062),
            .in1(N__4200),
            .in2(_gnd_net_),
            .in3(N__4173),
            .lcout(N_67),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_1_LC_10_5_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_1_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_1_LC_10_5_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_1_LC_10_5_0  (
            .in0(_gnd_net_),
            .in1(N__4314),
            .in2(_gnd_net_),
            .in3(N__4290),
            .lcout(\U409_TRANSFER_ACK.CO1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_10_7_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_10_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_10_7_1 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_10_7_1  (
            .in0(N__4084),
            .in1(N__4095),
            .in2(N__4126),
            .in3(N__4564),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net ),
            .ce(),
            .sr(N__5650));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_8_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_8_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_8_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_8_3  (
            .in0(N__4942),
            .in1(N__4096),
            .in2(N__4122),
            .in3(N__4878),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_10_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_10_9_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_10_9_5  (
            .in0(_gnd_net_),
            .in1(N__4938),
            .in2(_gnd_net_),
            .in3(N__4871),
            .lcout(\U409_TRANSFER_ACK.N_106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_10_13_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_10_13_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_10_13_5  (
            .in0(N__4075),
            .in1(N__4063),
            .in2(N__4918),
            .in3(N__4859),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_0_3_LC_11_5_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_0_3_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_0_3_LC_11_5_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_0_3_LC_11_5_2  (
            .in0(N__4287),
            .in1(N__4717),
            .in2(N__4696),
            .in3(N__4311),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20 ),
            .ltout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIERIJ7_3_LC_11_5_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIERIJ7_3_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIERIJ7_3_LC_11_5_3 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIERIJ7_3_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(N__4401),
            .in2(N__4411),
            .in3(N__4359),
            .lcout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0 ),
            .ltout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_11_5_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_11_5_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_11_5_4 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_11_5_4  (
            .in0(N__4288),
            .in1(_gnd_net_),
            .in2(N__4408),
            .in3(N__4313),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__5640));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_3_LC_11_5_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_3_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_3_LC_11_5_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_3_LC_11_5_5  (
            .in0(N__4312),
            .in1(N__4689),
            .in2(N__4720),
            .in3(N__4286),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_11_5_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_11_5_6 .LUT_INIT=16'b1111101001010101;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_11_5_6  (
            .in0(N__4289),
            .in1(_gnd_net_),
            .in2(N__4405),
            .in3(N__4371),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__5640));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_6_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_6_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_6_0 .LUT_INIT=16'b0100111001001100;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_6_0  (
            .in0(N__5123),
            .in1(N__4552),
            .in2(N__5152),
            .in3(N__4651),
            .lcout(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(N__5649));
    defparam \U409_TRANSFER_ACK.ROMENn_LC_11_6_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_11_6_1 .SEQ_MODE=4'b1001;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_11_6_1 .LUT_INIT=16'b1111101101110000;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_LC_11_6_1  (
            .in0(N__4400),
            .in1(N__4372),
            .in2(N__4332),
            .in3(N__4360),
            .lcout(ROMENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(N__5649));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_11_6_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_11_6_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_11_6_2  (
            .in0(_gnd_net_),
            .in1(N__4740),
            .in2(_gnd_net_),
            .in3(N__4694),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(N__5649));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_11_6_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_11_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_11_6_6 .LUT_INIT=16'b1011101000101010;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_LC_11_6_6  (
            .in0(N__4539),
            .in1(N__4315),
            .in2(N__4666),
            .in3(N__4291),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(N__5649));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_11_7_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_11_7_0 .LUT_INIT=16'b0000011111110111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_11_7_0  (
            .in0(N__5074),
            .in1(N__5094),
            .in2(N__5128),
            .in3(N__4650),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_7_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_7_1 .LUT_INIT=16'b0000001010001010;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_7_1  (
            .in0(N__5276),
            .in1(N__5151),
            .in2(N__4567),
            .in3(N__4657),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_7_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_7_2 .LUT_INIT=16'b0100000001000100;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_7_2  (
            .in0(N__4461),
            .in1(N__5277),
            .in2(N__4492),
            .in3(N__4440),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNINULI_LC_11_7_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNINULI_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNINULI_LC_11_7_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNINULI_LC_11_7_3  (
            .in0(N__4563),
            .in1(N__4551),
            .in2(N__4540),
            .in3(N__4639),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER6 ),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_11_7_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_11_7_4 .LUT_INIT=16'b1011101100110111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_11_7_4  (
            .in0(N__4459),
            .in1(N__5279),
            .in2(N__4525),
            .in3(N__4482),
            .lcout(\U409_TRANSFER_ACK.TACK_OUTn_0_sqmuxa_0_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_7_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_7_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_7_5  (
            .in0(N__5278),
            .in1(N__4486),
            .in2(_gnd_net_),
            .in3(N__4460),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_7_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_7_6 .LUT_INIT=16'b0010001100100111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_7_6  (
            .in0(N__4458),
            .in1(N__4505),
            .in2(N__4491),
            .in3(N__4439),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_11_7_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_11_7_7 .LUT_INIT=16'b0000111110101010;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_LC_11_7_7  (
            .in0(N__4506),
            .in1(_gnd_net_),
            .in2(N__4522),
            .in3(N__5291),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_11_8_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_11_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_11_8_0 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_i_LC_11_8_0  (
            .in0(N__4490),
            .in1(N__4462),
            .in2(N__5312),
            .in3(N__4441),
            .lcout(TACK_EN_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_EN_iC_net ),
            .ce(N__4426),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_10_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_10_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_10_1 .LUT_INIT=16'b0010001011111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_10_1  (
            .in0(N__4638),
            .in1(N__4788),
            .in2(_gnd_net_),
            .in3(N__4615),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ),
            .ce(),
            .sr(N__5466));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_7_LC_11_11_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_7_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_7_LC_11_11_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_7_LC_11_11_0  (
            .in0(N__4594),
            .in1(N__4577),
            .in2(N__5023),
            .in3(N__5044),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_11_11_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_11_11_1 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_11_11_1  (
            .in0(N__5516),
            .in1(N__4986),
            .in2(N__4624),
            .in3(N__5055),
            .lcout(\U409_TRANSFER_ACK.N_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_0_7_LC_11_11_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_0_7_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_0_7_LC_11_11_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_0_7_LC_11_11_3  (
            .in0(N__4578),
            .in1(N__5019),
            .in2(N__4600),
            .in3(N__5045),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a4_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_3_LC_11_11_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_3_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_3_LC_11_11_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_3_LC_11_11_4  (
            .in0(N__5056),
            .in1(N__4985),
            .in2(N__4621),
            .in3(N__5515),
            .lcout(\U409_TRANSFER_ACK.N_70 ),
            .ltout(\U409_TRANSFER_ACK.N_70_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_3_LC_11_11_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_3_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_3_LC_11_11_5 .LUT_INIT=16'b0010000011111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_3_LC_11_11_5  (
            .in0(N__4861),
            .in1(N__4931),
            .in2(N__4618),
            .in3(N__4614),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_11_6 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_11_6 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(N__4599),
            .in2(N__4603),
            .in3(N__4950),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ),
            .ce(),
            .sr(N__5467));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_11_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_11_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_11_7 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_11_7  (
            .in0(N__4579),
            .in1(N__4595),
            .in2(N__4954),
            .in3(N__5573),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ),
            .ce(),
            .sr(N__5467));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_12_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_12_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_12_2 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_12_2  (
            .in0(N__4776),
            .in1(N__4991),
            .in2(_gnd_net_),
            .in3(N__5568),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net ),
            .ce(),
            .sr(N__5452));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_12_3 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_12_3 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_12_3  (
            .in0(N__4992),
            .in1(N__4777),
            .in2(N__5575),
            .in3(N__5022),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net ),
            .ce(),
            .sr(N__5452));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_11_12_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_11_12_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_11_12_5  (
            .in0(N__5518),
            .in1(N__5487),
            .in2(_gnd_net_),
            .in3(N__5545),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_12_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_12_6 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_12_6 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_12_6  (
            .in0(N__4765),
            .in1(N__5047),
            .in2(N__4768),
            .in3(N__5569),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net ),
            .ce(),
            .sr(N__5452));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_11_13_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_11_13_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__4990),
            .in2(_gnd_net_),
            .in3(N__5021),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_1_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_1_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_1_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_1_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_12_5_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_12_5_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_12_5_6 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_12_5_6  (
            .in0(N__4719),
            .in1(N__4695),
            .in2(N__4744),
            .in3(N__4726),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net ),
            .ce(),
            .sr(N__5624));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_12_6_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_12_6_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_12_6_3  (
            .in0(_gnd_net_),
            .in1(N__4718),
            .in2(_gnd_net_),
            .in3(N__4693),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_EN_e_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_12_7_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_12_7_0 .LUT_INIT=16'b0001111100010000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_12_7_0  (
            .in0(N__5073),
            .in1(N__5092),
            .in2(N__5124),
            .in3(N__5161),
            .lcout(\U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIA48I_1_LC_12_7_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIA48I_1_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIA48I_1_LC_12_7_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_RNIA48I_1_LC_12_7_3  (
            .in0(N__4840),
            .in1(N__5170),
            .in2(_gnd_net_),
            .in3(N__5184),
            .lcout(\U409_TRANSFER_ACK.N_17_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_12_7_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_12_7_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_12_7_5  (
            .in0(_gnd_net_),
            .in1(N__5169),
            .in2(_gnd_net_),
            .in3(N__5183),
            .lcout(\U409_TRANSFER_ACK.N_3_0 ),
            .ltout(\U409_TRANSFER_ACK.N_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_7_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_7_6 .LUT_INIT=16'b0000010100100111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_7_6  (
            .in0(N__5115),
            .in1(N__5093),
            .in2(N__5155),
            .in3(N__5072),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.N_6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_7_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_7_7 .LUT_INIT=16'b0010101000001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_7_7  (
            .in0(N__5269),
            .in1(N__5150),
            .in2(N__5131),
            .in3(N__5119),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_8_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_8_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_8_1  (
            .in0(N__5249),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6795),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .ce(),
            .sr(N__5645));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_8_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5095),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .ce(),
            .sr(N__5645));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_12_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_12_11_2 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5548),
            .in3(N__5485),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_12_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_12_11_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_12_11_6  (
            .in0(N__5046),
            .in1(N__5020),
            .in2(N__4993),
            .in3(N__5486),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_12_11_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_12_11_7 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(N__5517),
            .in2(N__4957),
            .in3(N__5544),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_12_12_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_12_12_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_12_12_0 .LUT_INIT=16'b1101110000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_12_12_0  (
            .in0(N__4930),
            .in1(N__5519),
            .in2(N__4860),
            .in3(N__4789),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5462));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_12_12_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_12_12_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_12_12_1 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_12_12_1  (
            .in0(N__5520),
            .in1(N__5546),
            .in2(_gnd_net_),
            .in3(N__5574),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5462));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_12_12_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_12_12_4 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_12_12_4 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_12_12_4  (
            .in0(N__5547),
            .in1(N__5521),
            .in2(_gnd_net_),
            .in3(N__5488),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5462));
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_13_3_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_13_3_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_13_3_0 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_13_3_0  (
            .in0(_gnd_net_),
            .in1(N__5428),
            .in2(_gnd_net_),
            .in3(N__5350),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS1n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_13_3_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_13_3_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_13_3_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_13_3_5  (
            .in0(N__5349),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5389),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS0n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNI692L_0_LC_13_4_0 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNI692L_0_LC_13_4_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNI692L_0_LC_13_4_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_CIA.VMA_RNI692L_0_LC_13_4_0  (
            .in0(N__5267),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6796),
            .lcout(CIA_ENABLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_13_5_4.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_13_5_4.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_13_5_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_13_5_4 (
            .in0(N__5268),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_13_7_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_13_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_13_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_0_LC_13_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6843),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .ce(),
            .sr(N__5641));
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_13_7_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_13_7_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_13_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_1_LC_13_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5185),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .ce(),
            .sr(N__5641));
    defparam \U409_TICK.COUNTER60_9_LC_13_8_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_9_LC_13_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_9_LC_13_8_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_9_LC_13_8_0  (
            .in0(N__5699),
            .in1(N__5733),
            .in2(N__5776),
            .in3(N__6238),
            .lcout(\U409_TICK.COUNTER60Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6460),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_13_8_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_13_8_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_TICK.COUNTER60_RNIHJU51_4_LC_13_8_1  (
            .in0(N__6007),
            .in1(N__6031),
            .in2(_gnd_net_),
            .in3(N__6085),
            .lcout(),
            .ltout(\U409_TICK.TICK603_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_13_8_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_13_8_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_TICK.COUNTER60_RNI335G2_11_LC_13_8_2  (
            .in0(N__6214),
            .in1(N__5587),
            .in2(N__5593),
            .in3(N__6046),
            .lcout(\U409_TICK.TICK603_14 ),
            .ltout(\U409_TICK.TICK603_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_4_LC_13_8_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_4_LC_13_8_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_4_LC_13_8_3 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \U409_TICK.COUNTER60_4_LC_13_8_3  (
            .in0(N__6019),
            .in1(N__5700),
            .in2(N__5590),
            .in3(N__5774),
            .lcout(\U409_TICK.COUNTER60Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6460),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_14_LC_13_8_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_14_LC_13_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_14_LC_13_8_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_14_LC_13_8_4  (
            .in0(N__5698),
            .in1(N__5732),
            .in2(N__5775),
            .in3(N__6157),
            .lcout(\U409_TICK.COUNTER60Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6460),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_13_8_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_13_8_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER60_RNIDB4S_16_LC_13_8_5  (
            .in0(N__6199),
            .in1(N__6061),
            .in2(N__6112),
            .in3(N__6123),
            .lcout(\U409_TICK.TICK603_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_13_8_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_13_8_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_TICK.COUNTER60_RNI2USG_10_LC_13_8_6  (
            .in0(N__6184),
            .in1(N__6229),
            .in2(N__5965),
            .in3(N__6148),
            .lcout(\U409_TICK.TICK603_10 ),
            .ltout(\U409_TICK.TICK603_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_15_LC_13_8_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_15_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_15_LC_13_8_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_15_LC_13_8_7  (
            .in0(N__5731),
            .in1(N__5773),
            .in2(N__5581),
            .in3(N__6136),
            .lcout(\U409_TICK.COUNTER60Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6460),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_14_3_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_14_3_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_14_3_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U409_TICK.COUNTER50_RNII24V_14_LC_14_3_0  (
            .in0(N__6526),
            .in1(N__6499),
            .in2(N__6355),
            .in3(N__6280),
            .lcout(\U409_TICK.TICK503_10 ),
            .ltout(\U409_TICK.TICK503_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_15_LC_14_3_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_15_LC_14_3_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_15_LC_14_3_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_15_LC_14_3_1  (
            .in0(N__5845),
            .in1(N__5908),
            .in2(N__5578),
            .in3(N__6487),
            .lcout(\U409_TICK.COUNTER50Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6456),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_5_LC_14_3_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_5_LC_14_3_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_5_LC_14_3_2 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_5_LC_14_3_2  (
            .in0(N__5909),
            .in1(N__5874),
            .in2(N__6322),
            .in3(N__5849),
            .lcout(\U409_TICK.COUNTER50Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6456),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_1_LC_14_3_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_1_LC_14_3_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_1_LC_14_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_TICK.COUNTER50_1_LC_14_3_3  (
            .in0(_gnd_net_),
            .in1(N__6432),
            .in2(_gnd_net_),
            .in3(N__6413),
            .lcout(\U409_TICK.COUNTER50Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6456),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_3_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_3_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_3_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_3_4  (
            .in0(N__6265),
            .in1(N__6385),
            .in2(N__6433),
            .in3(N__6474),
            .lcout(\U409_TICK.TICK503_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK50_LC_14_3_5 .C_ON=1'b0;
    defparam \U409_TICK.TICK50_LC_14_3_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK50_LC_14_3_5 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \U409_TICK.TICK50_LC_14_3_5  (
            .in0(N__5876),
            .in1(N__5664),
            .in2(N__5851),
            .in3(N__5911),
            .lcout(TICK50_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6456),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_6_LC_14_3_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_6_LC_14_3_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_6_LC_14_3_6 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_6_LC_14_3_6  (
            .in0(N__5910),
            .in1(N__5875),
            .in2(N__6295),
            .in3(N__5850),
            .lcout(\U409_TICK.COUNTER50Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6456),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_11_LC_14_4_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_11_LC_14_4_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_11_LC_14_4_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_11_LC_14_4_0  (
            .in0(N__5878),
            .in1(N__5905),
            .in2(N__5843),
            .in3(N__6571),
            .lcout(\U409_TICK.COUNTER50Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6457),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_14_4_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_14_4_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_14_4_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNIH14V_11_LC_14_4_1  (
            .in0(N__6583),
            .in1(N__6619),
            .in2(N__6310),
            .in3(N__6547),
            .lcout(\U409_TICK.TICK503_9 ),
            .ltout(\U409_TICK.TICK503_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_0_LC_14_4_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_0_LC_14_4_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_0_LC_14_4_2 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \U409_TICK.COUNTER50_0_LC_14_4_2  (
            .in0(N__5877),
            .in1(N__6415),
            .in2(N__5653),
            .in3(N__5904),
            .lcout(\U409_TICK.COUNTER50Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6457),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_14_4_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_14_4_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_14_4_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_TICK.COUNTER50_RNID6CP_3_LC_14_4_3  (
            .in0(N__6370),
            .in1(N__6336),
            .in2(_gnd_net_),
            .in3(N__6409),
            .lcout(),
            .ltout(\U409_TICK.TICK503_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_14_4_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_14_4_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_14_4_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER50_RNITU182_10_LC_14_4_4  (
            .in0(N__5923),
            .in1(N__6562),
            .in2(N__5917),
            .in3(N__6598),
            .lcout(\U409_TICK.TICK503_14 ),
            .ltout(\U409_TICK.TICK503_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_9_LC_14_4_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_9_LC_14_4_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_9_LC_14_4_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_9_LC_14_4_5  (
            .in0(N__5842),
            .in1(N__5881),
            .in2(N__5914),
            .in3(N__6607),
            .lcout(\U409_TICK.COUNTER50Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6457),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_13_LC_14_4_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_13_LC_14_4_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_13_LC_14_4_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_13_LC_14_4_6  (
            .in0(N__5879),
            .in1(N__5906),
            .in2(N__5844),
            .in3(N__6535),
            .lcout(\U409_TICK.COUNTER50Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6457),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_14_LC_14_4_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_14_LC_14_4_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_14_LC_14_4_7 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_14_LC_14_4_7  (
            .in0(N__5907),
            .in1(N__5880),
            .in2(N__6514),
            .in3(N__5832),
            .lcout(\U409_TICK.COUNTER50Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6457),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_8_LC_14_7_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_8_LC_14_7_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_8_LC_14_7_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_8_LC_14_7_0  (
            .in0(N__5734),
            .in1(N__5766),
            .in2(N__5707),
            .in3(N__5932),
            .lcout(\U409_TICK.COUNTER60Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6461),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK60_LC_14_7_1 .C_ON=1'b0;
    defparam \U409_TICK.TICK60_LC_14_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK60_LC_14_7_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \U409_TICK.TICK60_LC_14_7_1  (
            .in0(N__5765),
            .in1(N__5790),
            .in2(N__5743),
            .in3(N__5702),
            .lcout(TICK60_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6461),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_14_7_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_14_7_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER60_RNICDC71_14_LC_14_7_2  (
            .in0(N__6250),
            .in1(N__5944),
            .in2(N__5992),
            .in3(N__6169),
            .lcout(\U409_TICK.TICK603_9 ),
            .ltout(\U409_TICK.TICK603_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_6_LC_14_7_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_6_LC_14_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_6_LC_14_7_3 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \U409_TICK.COUNTER60_6_LC_14_7_3  (
            .in0(N__5974),
            .in1(N__5701),
            .in2(N__5779),
            .in3(N__5736),
            .lcout(\U409_TICK.COUNTER60Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6461),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_0_LC_14_7_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_0_LC_14_7_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_0_LC_14_7_5 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U409_TICK.COUNTER60_0_LC_14_7_5  (
            .in0(N__5764),
            .in1(N__5735),
            .in2(N__6091),
            .in3(N__5706),
            .lcout(\U409_TICK.COUNTER60Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6461),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_1_LC_14_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_1_LC_14_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_1_LC_14_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_TICK.COUNTER60_1_LC_14_7_7  (
            .in0(_gnd_net_),
            .in1(N__6086),
            .in2(_gnd_net_),
            .in3(N__6111),
            .lcout(\U409_TICK.COUNTER60Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6461),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_14_8_0 .C_ON=1'b1;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_14_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(N__6107),
            .in2(N__6090),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_8_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_2_LC_14_8_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_2_LC_14_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_2_LC_14_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_2_LC_14_8_1  (
            .in0(_gnd_net_),
            .in1(N__6060),
            .in2(_gnd_net_),
            .in3(N__6049),
            .lcout(\U409_TICK.COUNTER60Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .clk(N__6462),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_3_LC_14_8_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_3_LC_14_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_3_LC_14_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_3_LC_14_8_2  (
            .in0(_gnd_net_),
            .in1(N__6045),
            .in2(_gnd_net_),
            .in3(N__6034),
            .lcout(\U409_TICK.COUNTER60Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .clk(N__6462),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_14_8_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_14_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_4_LC_14_8_3  (
            .in0(_gnd_net_),
            .in1(N__6030),
            .in2(_gnd_net_),
            .in3(N__6010),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_5_LC_14_8_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_5_LC_14_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_5_LC_14_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_5_LC_14_8_4  (
            .in0(_gnd_net_),
            .in1(N__6006),
            .in2(_gnd_net_),
            .in3(N__5995),
            .lcout(\U409_TICK.COUNTER60Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .clk(N__6462),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_14_8_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_14_8_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_6_LC_14_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5991),
            .in3(N__5968),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_7_LC_14_8_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_7_LC_14_8_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_7_LC_14_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_7_LC_14_8_6  (
            .in0(_gnd_net_),
            .in1(N__5958),
            .in2(_gnd_net_),
            .in3(N__5947),
            .lcout(\U409_TICK.COUNTER60Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .clk(N__6462),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_14_8_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_14_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_8_LC_14_8_7  (
            .in0(_gnd_net_),
            .in1(N__5943),
            .in2(_gnd_net_),
            .in3(N__5926),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_14_9_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_14_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_9_LC_14_9_0  (
            .in0(_gnd_net_),
            .in1(N__6249),
            .in2(_gnd_net_),
            .in3(N__6232),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_14_9_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_10_LC_14_9_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_10_LC_14_9_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_10_LC_14_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_10_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(N__6228),
            .in2(_gnd_net_),
            .in3(N__6217),
            .lcout(\U409_TICK.COUNTER60Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .clk(N__6463),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_11_LC_14_9_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_11_LC_14_9_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_11_LC_14_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_11_LC_14_9_2  (
            .in0(_gnd_net_),
            .in1(N__6213),
            .in2(_gnd_net_),
            .in3(N__6202),
            .lcout(\U409_TICK.COUNTER60Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .clk(N__6463),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_12_LC_14_9_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_12_LC_14_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_12_LC_14_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_12_LC_14_9_3  (
            .in0(_gnd_net_),
            .in1(N__6198),
            .in2(_gnd_net_),
            .in3(N__6187),
            .lcout(\U409_TICK.COUNTER60Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .clk(N__6463),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_13_LC_14_9_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_13_LC_14_9_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_13_LC_14_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_13_LC_14_9_4  (
            .in0(_gnd_net_),
            .in1(N__6183),
            .in2(_gnd_net_),
            .in3(N__6172),
            .lcout(\U409_TICK.COUNTER60Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .clk(N__6463),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_14_9_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_14_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_14_LC_14_9_5  (
            .in0(_gnd_net_),
            .in1(N__6168),
            .in2(_gnd_net_),
            .in3(N__6151),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_14_9_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_14_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_15_LC_14_9_6  (
            .in0(_gnd_net_),
            .in1(N__6147),
            .in2(_gnd_net_),
            .in3(N__6130),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_16_LC_14_9_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_16_LC_14_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_16_LC_14_9_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER60_16_LC_14_9_7  (
            .in0(_gnd_net_),
            .in1(N__6124),
            .in2(_gnd_net_),
            .in3(N__6127),
            .lcout(\U409_TICK.COUNTER60Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6463),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_15_3_0 .C_ON=1'b1;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_15_3_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_15_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_15_3_0  (
            .in0(_gnd_net_),
            .in1(N__6428),
            .in2(N__6414),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_3_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_2_LC_15_3_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_2_LC_15_3_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_2_LC_15_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_2_LC_15_3_1  (
            .in0(_gnd_net_),
            .in1(N__6384),
            .in2(_gnd_net_),
            .in3(N__6373),
            .lcout(\U409_TICK.COUNTER50Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .clk(N__6458),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_3_LC_15_3_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_3_LC_15_3_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_3_LC_15_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_3_LC_15_3_2  (
            .in0(_gnd_net_),
            .in1(N__6369),
            .in2(_gnd_net_),
            .in3(N__6358),
            .lcout(\U409_TICK.COUNTER50Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .clk(N__6458),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_4_LC_15_3_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_4_LC_15_3_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_4_LC_15_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_4_LC_15_3_3  (
            .in0(_gnd_net_),
            .in1(N__6351),
            .in2(_gnd_net_),
            .in3(N__6340),
            .lcout(\U409_TICK.COUNTER50Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .clk(N__6458),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_15_3_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_15_3_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_15_3_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_5_LC_15_3_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6337),
            .in3(N__6313),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_15_3_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_15_3_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_15_3_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_6_LC_15_3_5  (
            .in0(_gnd_net_),
            .in1(N__6306),
            .in2(_gnd_net_),
            .in3(N__6283),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_7_LC_15_3_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_7_LC_15_3_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_7_LC_15_3_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_7_LC_15_3_6  (
            .in0(_gnd_net_),
            .in1(N__6279),
            .in2(_gnd_net_),
            .in3(N__6268),
            .lcout(\U409_TICK.COUNTER50Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .clk(N__6458),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_8_LC_15_3_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_8_LC_15_3_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_8_LC_15_3_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_8_LC_15_3_7  (
            .in0(_gnd_net_),
            .in1(N__6264),
            .in2(_gnd_net_),
            .in3(N__6253),
            .lcout(\U409_TICK.COUNTER50Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .clk(N__6458),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_15_4_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_15_4_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_15_4_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_9_LC_15_4_0  (
            .in0(_gnd_net_),
            .in1(N__6618),
            .in2(_gnd_net_),
            .in3(N__6601),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_15_4_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_10_LC_15_4_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_10_LC_15_4_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_10_LC_15_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_10_LC_15_4_1  (
            .in0(_gnd_net_),
            .in1(N__6597),
            .in2(_gnd_net_),
            .in3(N__6586),
            .lcout(\U409_TICK.COUNTER50Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .clk(N__6459),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_15_4_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_15_4_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_15_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_11_LC_15_4_2  (
            .in0(_gnd_net_),
            .in1(N__6582),
            .in2(_gnd_net_),
            .in3(N__6565),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_12_LC_15_4_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_12_LC_15_4_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_12_LC_15_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_12_LC_15_4_3  (
            .in0(_gnd_net_),
            .in1(N__6561),
            .in2(_gnd_net_),
            .in3(N__6550),
            .lcout(\U409_TICK.COUNTER50Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .clk(N__6459),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_15_4_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_15_4_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_15_4_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_13_LC_15_4_4  (
            .in0(_gnd_net_),
            .in1(N__6546),
            .in2(_gnd_net_),
            .in3(N__6529),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_15_4_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_15_4_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_15_4_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_14_LC_15_4_5  (
            .in0(_gnd_net_),
            .in1(N__6525),
            .in2(_gnd_net_),
            .in3(N__6502),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_15_4_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_15_4_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_15_4_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_15_LC_15_4_6  (
            .in0(_gnd_net_),
            .in1(N__6498),
            .in2(_gnd_net_),
            .in3(N__6481),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_16_LC_15_4_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_16_LC_15_4_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_16_LC_15_4_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER50_16_LC_15_4_7  (
            .in0(_gnd_net_),
            .in1(N__6475),
            .in2(_gnd_net_),
            .in3(N__6478),
            .lcout(\U409_TICK.COUNTER50Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6459),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_15_6_0 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_15_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_15_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_15_6_0  (
            .in0(_gnd_net_),
            .in1(N__6969),
            .in2(N__7003),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_6_0_),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_15_6_1 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_15_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_15_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_2_LC_15_6_1  (
            .in0(_gnd_net_),
            .in1(N__6753),
            .in2(_gnd_net_),
            .in3(N__6655),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .clk(N__6940),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_15_6_2 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_15_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_15_6_2 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_3_LC_15_6_2  (
            .in0(N__6765),
            .in1(_gnd_net_),
            .in2(N__6637),
            .in3(N__6652),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .clk(N__6940),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_15_6_3 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_15_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_15_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_4_LC_15_6_3  (
            .in0(_gnd_net_),
            .in1(N__6702),
            .in2(_gnd_net_),
            .in3(N__6649),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .clk(N__6940),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_15_6_4 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_15_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_15_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_5_LC_15_6_4  (
            .in0(N__6766),
            .in1(N__6730),
            .in2(_gnd_net_),
            .in3(N__6646),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .clk(N__6940),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_15_6_5 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_15_6_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_15_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_6_LC_15_6_5  (
            .in0(_gnd_net_),
            .in1(N__6873),
            .in2(_gnd_net_),
            .in3(N__6643),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ),
            .clk(N__6940),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_15_6_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_15_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_15_6_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_7_LC_15_6_6  (
            .in0(_gnd_net_),
            .in1(N__6891),
            .in2(_gnd_net_),
            .in3(N__6640),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6940),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIMC921_7_LC_15_6_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIMC921_7_LC_15_6_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIMC921_7_LC_15_6_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIMC921_7_LC_15_6_7  (
            .in0(N__6890),
            .in1(N__6872),
            .in2(_gnd_net_),
            .in3(N__6632),
            .lcout(\U409_CIA.N_104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_2_LC_15_7_0 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_2_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_2_LC_15_7_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_2_LC_15_7_0  (
            .in0(N__6994),
            .in1(N__6700),
            .in2(_gnd_net_),
            .in3(N__6636),
            .lcout(),
            .ltout(\U409_CIA.un1_CIA_CLK_COUNT_2_0_a4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_15_7_1 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_15_7_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_15_7_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_1_LC_15_7_1  (
            .in0(N__6709),
            .in1(N__6892),
            .in2(N__6877),
            .in3(N__6874),
            .lcout(),
            .ltout(\U409_CIA.CLK_CIA_RNOZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_LC_15_7_2 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_LC_15_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CLK_CIA_LC_15_7_2 .LUT_INIT=16'b0011001100110000;
    LogicCell40 \U409_CIA.CLK_CIA_LC_15_7_2  (
            .in0(_gnd_net_),
            .in1(N__6661),
            .in2(N__6859),
            .in3(N__6836),
            .lcout(CLK_CIA_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6938),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_1_LC_15_7_3 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_1_LC_15_7_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_1_LC_15_7_3 .LUT_INIT=16'b0101000010100000;
    LogicCell40 \U409_CIA.VMA_RNO_1_LC_15_7_3  (
            .in0(N__6701),
            .in1(_gnd_net_),
            .in2(N__6970),
            .in3(N__6995),
            .lcout(),
            .ltout(\U409_CIA.un1_CIA_CLK_COUNT_3_0_a4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_0_LC_15_7_4 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_0_LC_15_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_0_LC_15_7_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_CIA.VMA_RNO_0_LC_15_7_4  (
            .in0(N__6675),
            .in1(N__6757),
            .in2(N__6820),
            .in3(N__6728),
            .lcout(),
            .ltout(\U409_CIA.VMA_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_LC_15_7_5 .C_ON=1'b0;
    defparam \U409_CIA.VMA_LC_15_7_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.VMA_LC_15_7_5 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \U409_CIA.VMA_LC_15_7_5  (
            .in0(N__6817),
            .in1(N__6782),
            .in2(N__6799),
            .in3(N__6997),
            .lcout(\U409_CIA.VMAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6938),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_2_LC_15_7_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_2_LC_15_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_2_LC_15_7_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIH7921_2_LC_15_7_6  (
            .in0(N__6752),
            .in1(N__6727),
            .in2(_gnd_net_),
            .in3(N__6699),
            .lcout(),
            .ltout(\U409_CIA.CIA_CLK_COUNT11_0_a4_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNICTDR2_0_LC_15_7_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNICTDR2_0_LC_15_7_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNICTDR2_0_LC_15_7_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNICTDR2_0_LC_15_7_7  (
            .in0(N__6968),
            .in1(N__6996),
            .in2(N__6769),
            .in3(N__6674),
            .lcout(\U409_CIA.CIA_CLK_COUNT11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNID3921_2_LC_16_6_0 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNID3921_2_LC_16_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNID3921_2_LC_16_6_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNID3921_2_LC_16_6_0  (
            .in0(N__6962),
            .in1(N__6751),
            .in2(_gnd_net_),
            .in3(N__6729),
            .lcout(\U409_CIA.CLK_CIA6_1 ),
            .ltout(\U409_CIA.CLK_CIA6_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_16_6_1 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_16_6_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_16_6_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_0_LC_16_6_1  (
            .in0(N__7001),
            .in1(N__6703),
            .in2(N__6679),
            .in3(N__6676),
            .lcout(\U409_CIA.CLK_CIA6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_16_6_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_16_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_16_6_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_1_LC_16_6_4  (
            .in0(N__6964),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7002),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6939),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_16_6_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_16_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_16_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_0_LC_16_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6963),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6939),
            .ce(),
            .sr(_gnd_net_));
    defparam TACKn_iobuf_RNO_LC_16_13_3.C_ON=1'b0;
    defparam TACKn_iobuf_RNO_LC_16_13_3.SEQ_MODE=4'b0000;
    defparam TACKn_iobuf_RNO_LC_16_13_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 TACKn_iobuf_RNO_LC_16_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6925),
            .lcout(N_465_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U409_TOP

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Sep 14 2025 12:26:09

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U409_TOP" view "INTERFACE"

module U409_TOP (
    ROM_DELAY,
    TM,
    TT,
    A,
    D,
    RESETn,
    OVL,
    CONFIGENn,
    PPIO,
    PORTSIZE,
    TICK60,
    PCS1,
    CIACS0n,
    SCS0,
    CPUCONFn,
    CLK6,
    AGNUS_CLK,
    CLK_CIA,
    BUFENn,
    AUTOBOOT,
    RnW,
    XCLK,
    CIACS1n,
    PPIO_J,
    TICK50,
    TCIn,
    TBIn,
    RAMSPACEn,
    PCS0,
    CLK40_IN,
    CLK28_IN,
    XCLK_ENn,
    SCS1,
    REGSPACEn,
    F_ENn,
    TSn,
    SPIO_J,
    SPIO,
    RTC_ENn,
    ATA_ENn,
    TACKn,
    ROMENn);

    input [1:0] ROM_DELAY;
    input [2:0] TM;
    input [1:0] TT;
    input [31:1] A;
    inout [7:4] D;
    input RESETn;
    input OVL;
    output CONFIGENn;
    output PPIO;
    output PORTSIZE;
    output TICK60;
    output PCS1;
    output CIACS0n;
    output SCS0;
    input CPUCONFn;
    input CLK6;
    output AGNUS_CLK;
    output CLK_CIA;
    output BUFENn;
    input AUTOBOOT;
    input RnW;
    input XCLK;
    output CIACS1n;
    input PPIO_J;
    output TICK50;
    output TCIn;
    output TBIn;
    output RAMSPACEn;
    output PCS0;
    input CLK40_IN;
    input CLK28_IN;
    input XCLK_ENn;
    output SCS1;
    output REGSPACEn;
    output F_ENn;
    input TSn;
    input SPIO_J;
    output SPIO;
    output RTC_ENn;
    output ATA_ENn;
    inout TACKn;
    output ROMENn;

    wire N__11848;
    wire N__11847;
    wire N__11846;
    wire N__11838;
    wire N__11837;
    wire N__11836;
    wire N__11828;
    wire N__11827;
    wire N__11826;
    wire N__11817;
    wire N__11816;
    wire N__11815;
    wire N__11808;
    wire N__11807;
    wire N__11806;
    wire N__11799;
    wire N__11798;
    wire N__11797;
    wire N__11790;
    wire N__11789;
    wire N__11788;
    wire N__11781;
    wire N__11780;
    wire N__11779;
    wire N__11772;
    wire N__11771;
    wire N__11770;
    wire N__11763;
    wire N__11762;
    wire N__11761;
    wire N__11754;
    wire N__11753;
    wire N__11752;
    wire N__11745;
    wire N__11744;
    wire N__11743;
    wire N__11736;
    wire N__11735;
    wire N__11734;
    wire N__11727;
    wire N__11726;
    wire N__11725;
    wire N__11718;
    wire N__11717;
    wire N__11716;
    wire N__11709;
    wire N__11708;
    wire N__11707;
    wire N__11700;
    wire N__11699;
    wire N__11698;
    wire N__11691;
    wire N__11690;
    wire N__11689;
    wire N__11682;
    wire N__11681;
    wire N__11680;
    wire N__11673;
    wire N__11672;
    wire N__11671;
    wire N__11664;
    wire N__11663;
    wire N__11662;
    wire N__11655;
    wire N__11654;
    wire N__11653;
    wire N__11646;
    wire N__11645;
    wire N__11644;
    wire N__11637;
    wire N__11636;
    wire N__11635;
    wire N__11628;
    wire N__11627;
    wire N__11626;
    wire N__11619;
    wire N__11618;
    wire N__11617;
    wire N__11610;
    wire N__11609;
    wire N__11608;
    wire N__11601;
    wire N__11600;
    wire N__11599;
    wire N__11592;
    wire N__11591;
    wire N__11590;
    wire N__11583;
    wire N__11582;
    wire N__11581;
    wire N__11574;
    wire N__11573;
    wire N__11572;
    wire N__11565;
    wire N__11564;
    wire N__11563;
    wire N__11556;
    wire N__11555;
    wire N__11554;
    wire N__11547;
    wire N__11546;
    wire N__11545;
    wire N__11538;
    wire N__11537;
    wire N__11536;
    wire N__11529;
    wire N__11528;
    wire N__11527;
    wire N__11520;
    wire N__11519;
    wire N__11518;
    wire N__11511;
    wire N__11510;
    wire N__11509;
    wire N__11502;
    wire N__11501;
    wire N__11500;
    wire N__11493;
    wire N__11492;
    wire N__11491;
    wire N__11484;
    wire N__11483;
    wire N__11482;
    wire N__11475;
    wire N__11474;
    wire N__11473;
    wire N__11466;
    wire N__11465;
    wire N__11464;
    wire N__11457;
    wire N__11456;
    wire N__11455;
    wire N__11448;
    wire N__11447;
    wire N__11446;
    wire N__11439;
    wire N__11438;
    wire N__11437;
    wire N__11430;
    wire N__11429;
    wire N__11428;
    wire N__11421;
    wire N__11420;
    wire N__11419;
    wire N__11412;
    wire N__11411;
    wire N__11410;
    wire N__11403;
    wire N__11402;
    wire N__11401;
    wire N__11394;
    wire N__11393;
    wire N__11392;
    wire N__11385;
    wire N__11384;
    wire N__11383;
    wire N__11376;
    wire N__11375;
    wire N__11374;
    wire N__11367;
    wire N__11366;
    wire N__11365;
    wire N__11358;
    wire N__11357;
    wire N__11356;
    wire N__11349;
    wire N__11348;
    wire N__11347;
    wire N__11340;
    wire N__11339;
    wire N__11338;
    wire N__11331;
    wire N__11330;
    wire N__11329;
    wire N__11322;
    wire N__11321;
    wire N__11320;
    wire N__11313;
    wire N__11312;
    wire N__11311;
    wire N__11304;
    wire N__11303;
    wire N__11302;
    wire N__11295;
    wire N__11294;
    wire N__11293;
    wire N__11286;
    wire N__11285;
    wire N__11284;
    wire N__11277;
    wire N__11276;
    wire N__11275;
    wire N__11268;
    wire N__11267;
    wire N__11266;
    wire N__11259;
    wire N__11258;
    wire N__11257;
    wire N__11250;
    wire N__11249;
    wire N__11248;
    wire N__11241;
    wire N__11240;
    wire N__11239;
    wire N__11232;
    wire N__11231;
    wire N__11230;
    wire N__11223;
    wire N__11222;
    wire N__11221;
    wire N__11214;
    wire N__11213;
    wire N__11212;
    wire N__11205;
    wire N__11204;
    wire N__11203;
    wire N__11186;
    wire N__11183;
    wire N__11180;
    wire N__11177;
    wire N__11176;
    wire N__11173;
    wire N__11170;
    wire N__11167;
    wire N__11164;
    wire N__11161;
    wire N__11158;
    wire N__11153;
    wire N__11150;
    wire N__11149;
    wire N__11148;
    wire N__11147;
    wire N__11146;
    wire N__11143;
    wire N__11132;
    wire N__11129;
    wire N__11126;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11114;
    wire N__11111;
    wire N__11108;
    wire N__11105;
    wire N__11102;
    wire N__11099;
    wire N__11096;
    wire N__11093;
    wire N__11090;
    wire N__11089;
    wire N__11086;
    wire N__11083;
    wire N__11078;
    wire N__11075;
    wire N__11072;
    wire N__11069;
    wire N__11068;
    wire N__11065;
    wire N__11062;
    wire N__11057;
    wire N__11054;
    wire N__11051;
    wire N__11048;
    wire N__11045;
    wire N__11044;
    wire N__11041;
    wire N__11038;
    wire N__11033;
    wire N__11032;
    wire N__11031;
    wire N__11030;
    wire N__11029;
    wire N__11028;
    wire N__11025;
    wire N__11024;
    wire N__11023;
    wire N__11018;
    wire N__11015;
    wire N__11012;
    wire N__11003;
    wire N__10994;
    wire N__10993;
    wire N__10990;
    wire N__10989;
    wire N__10988;
    wire N__10987;
    wire N__10984;
    wire N__10983;
    wire N__10982;
    wire N__10981;
    wire N__10978;
    wire N__10975;
    wire N__10972;
    wire N__10969;
    wire N__10966;
    wire N__10959;
    wire N__10946;
    wire N__10945;
    wire N__10942;
    wire N__10941;
    wire N__10936;
    wire N__10933;
    wire N__10932;
    wire N__10931;
    wire N__10930;
    wire N__10929;
    wire N__10928;
    wire N__10925;
    wire N__10922;
    wire N__10911;
    wire N__10908;
    wire N__10901;
    wire N__10898;
    wire N__10895;
    wire N__10892;
    wire N__10891;
    wire N__10888;
    wire N__10885;
    wire N__10882;
    wire N__10877;
    wire N__10876;
    wire N__10875;
    wire N__10874;
    wire N__10873;
    wire N__10872;
    wire N__10871;
    wire N__10870;
    wire N__10869;
    wire N__10868;
    wire N__10847;
    wire N__10844;
    wire N__10841;
    wire N__10838;
    wire N__10835;
    wire N__10832;
    wire N__10829;
    wire N__10826;
    wire N__10823;
    wire N__10820;
    wire N__10817;
    wire N__10814;
    wire N__10811;
    wire N__10808;
    wire N__10805;
    wire N__10804;
    wire N__10801;
    wire N__10798;
    wire N__10793;
    wire N__10790;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10772;
    wire N__10769;
    wire N__10768;
    wire N__10767;
    wire N__10766;
    wire N__10763;
    wire N__10760;
    wire N__10757;
    wire N__10754;
    wire N__10749;
    wire N__10744;
    wire N__10741;
    wire N__10738;
    wire N__10735;
    wire N__10732;
    wire N__10727;
    wire N__10724;
    wire N__10721;
    wire N__10720;
    wire N__10717;
    wire N__10714;
    wire N__10709;
    wire N__10706;
    wire N__10703;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10691;
    wire N__10688;
    wire N__10685;
    wire N__10682;
    wire N__10681;
    wire N__10678;
    wire N__10675;
    wire N__10670;
    wire N__10667;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10655;
    wire N__10654;
    wire N__10651;
    wire N__10648;
    wire N__10643;
    wire N__10640;
    wire N__10639;
    wire N__10636;
    wire N__10633;
    wire N__10628;
    wire N__10625;
    wire N__10622;
    wire N__10619;
    wire N__10618;
    wire N__10615;
    wire N__10612;
    wire N__10607;
    wire N__10604;
    wire N__10601;
    wire N__10598;
    wire N__10595;
    wire N__10594;
    wire N__10591;
    wire N__10588;
    wire N__10583;
    wire N__10580;
    wire N__10577;
    wire N__10574;
    wire N__10573;
    wire N__10570;
    wire N__10567;
    wire N__10562;
    wire N__10559;
    wire N__10558;
    wire N__10555;
    wire N__10552;
    wire N__10547;
    wire N__10544;
    wire N__10541;
    wire N__10540;
    wire N__10537;
    wire N__10534;
    wire N__10529;
    wire N__10526;
    wire N__10523;
    wire N__10520;
    wire N__10519;
    wire N__10516;
    wire N__10513;
    wire N__10508;
    wire N__10507;
    wire N__10504;
    wire N__10501;
    wire N__10496;
    wire N__10493;
    wire N__10492;
    wire N__10489;
    wire N__10486;
    wire N__10481;
    wire N__10480;
    wire N__10477;
    wire N__10474;
    wire N__10469;
    wire N__10466;
    wire N__10463;
    wire N__10460;
    wire N__10459;
    wire N__10456;
    wire N__10453;
    wire N__10448;
    wire N__10447;
    wire N__10444;
    wire N__10443;
    wire N__10438;
    wire N__10435;
    wire N__10430;
    wire N__10429;
    wire N__10426;
    wire N__10425;
    wire N__10424;
    wire N__10421;
    wire N__10416;
    wire N__10413;
    wire N__10410;
    wire N__10403;
    wire N__10402;
    wire N__10399;
    wire N__10396;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10384;
    wire N__10381;
    wire N__10378;
    wire N__10373;
    wire N__10370;
    wire N__10367;
    wire N__10366;
    wire N__10363;
    wire N__10360;
    wire N__10357;
    wire N__10352;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10337;
    wire N__10336;
    wire N__10333;
    wire N__10330;
    wire N__10325;
    wire N__10322;
    wire N__10321;
    wire N__10320;
    wire N__10319;
    wire N__10318;
    wire N__10317;
    wire N__10314;
    wire N__10311;
    wire N__10310;
    wire N__10303;
    wire N__10294;
    wire N__10289;
    wire N__10288;
    wire N__10287;
    wire N__10286;
    wire N__10285;
    wire N__10284;
    wire N__10283;
    wire N__10272;
    wire N__10267;
    wire N__10262;
    wire N__10259;
    wire N__10258;
    wire N__10257;
    wire N__10256;
    wire N__10255;
    wire N__10254;
    wire N__10253;
    wire N__10250;
    wire N__10247;
    wire N__10236;
    wire N__10229;
    wire N__10226;
    wire N__10225;
    wire N__10222;
    wire N__10219;
    wire N__10214;
    wire N__10211;
    wire N__10208;
    wire N__10205;
    wire N__10204;
    wire N__10201;
    wire N__10198;
    wire N__10193;
    wire N__10190;
    wire N__10189;
    wire N__10186;
    wire N__10183;
    wire N__10178;
    wire N__10175;
    wire N__10172;
    wire N__10169;
    wire N__10166;
    wire N__10165;
    wire N__10164;
    wire N__10161;
    wire N__10158;
    wire N__10157;
    wire N__10154;
    wire N__10151;
    wire N__10146;
    wire N__10143;
    wire N__10136;
    wire N__10133;
    wire N__10130;
    wire N__10129;
    wire N__10126;
    wire N__10123;
    wire N__10118;
    wire N__10117;
    wire N__10114;
    wire N__10111;
    wire N__10106;
    wire N__10103;
    wire N__10102;
    wire N__10099;
    wire N__10096;
    wire N__10091;
    wire N__10088;
    wire N__10085;
    wire N__10082;
    wire N__10081;
    wire N__10080;
    wire N__10077;
    wire N__10072;
    wire N__10067;
    wire N__10064;
    wire N__10063;
    wire N__10062;
    wire N__10059;
    wire N__10058;
    wire N__10053;
    wire N__10050;
    wire N__10047;
    wire N__10044;
    wire N__10037;
    wire N__10036;
    wire N__10035;
    wire N__10034;
    wire N__10027;
    wire N__10024;
    wire N__10023;
    wire N__10020;
    wire N__10017;
    wire N__10016;
    wire N__10015;
    wire N__10012;
    wire N__10011;
    wire N__10006;
    wire N__10003;
    wire N__10000;
    wire N__9995;
    wire N__9986;
    wire N__9983;
    wire N__9982;
    wire N__9979;
    wire N__9976;
    wire N__9973;
    wire N__9970;
    wire N__9965;
    wire N__9962;
    wire N__9959;
    wire N__9958;
    wire N__9957;
    wire N__9956;
    wire N__9953;
    wire N__9950;
    wire N__9949;
    wire N__9940;
    wire N__9937;
    wire N__9936;
    wire N__9935;
    wire N__9934;
    wire N__9933;
    wire N__9932;
    wire N__9927;
    wire N__9924;
    wire N__9921;
    wire N__9918;
    wire N__9913;
    wire N__9910;
    wire N__9899;
    wire N__9896;
    wire N__9893;
    wire N__9890;
    wire N__9887;
    wire N__9884;
    wire N__9883;
    wire N__9880;
    wire N__9877;
    wire N__9872;
    wire N__9871;
    wire N__9870;
    wire N__9869;
    wire N__9866;
    wire N__9865;
    wire N__9864;
    wire N__9861;
    wire N__9858;
    wire N__9855;
    wire N__9852;
    wire N__9847;
    wire N__9846;
    wire N__9843;
    wire N__9842;
    wire N__9841;
    wire N__9840;
    wire N__9839;
    wire N__9838;
    wire N__9837;
    wire N__9834;
    wire N__9833;
    wire N__9832;
    wire N__9831;
    wire N__9830;
    wire N__9827;
    wire N__9826;
    wire N__9825;
    wire N__9824;
    wire N__9823;
    wire N__9822;
    wire N__9821;
    wire N__9820;
    wire N__9819;
    wire N__9818;
    wire N__9815;
    wire N__9812;
    wire N__9761;
    wire N__9758;
    wire N__9755;
    wire N__9752;
    wire N__9751;
    wire N__9750;
    wire N__9749;
    wire N__9748;
    wire N__9747;
    wire N__9746;
    wire N__9745;
    wire N__9744;
    wire N__9743;
    wire N__9740;
    wire N__9739;
    wire N__9738;
    wire N__9737;
    wire N__9736;
    wire N__9735;
    wire N__9734;
    wire N__9733;
    wire N__9732;
    wire N__9731;
    wire N__9692;
    wire N__9689;
    wire N__9686;
    wire N__9683;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9671;
    wire N__9668;
    wire N__9665;
    wire N__9662;
    wire N__9659;
    wire N__9656;
    wire N__9655;
    wire N__9652;
    wire N__9649;
    wire N__9646;
    wire N__9641;
    wire N__9638;
    wire N__9635;
    wire N__9632;
    wire N__9629;
    wire N__9628;
    wire N__9627;
    wire N__9624;
    wire N__9621;
    wire N__9620;
    wire N__9617;
    wire N__9614;
    wire N__9611;
    wire N__9606;
    wire N__9599;
    wire N__9598;
    wire N__9597;
    wire N__9594;
    wire N__9589;
    wire N__9584;
    wire N__9583;
    wire N__9582;
    wire N__9579;
    wire N__9576;
    wire N__9573;
    wire N__9566;
    wire N__9565;
    wire N__9562;
    wire N__9559;
    wire N__9554;
    wire N__9551;
    wire N__9548;
    wire N__9545;
    wire N__9542;
    wire N__9539;
    wire N__9536;
    wire N__9533;
    wire N__9530;
    wire N__9527;
    wire N__9524;
    wire N__9523;
    wire N__9520;
    wire N__9517;
    wire N__9512;
    wire N__9509;
    wire N__9508;
    wire N__9505;
    wire N__9500;
    wire N__9497;
    wire N__9494;
    wire N__9491;
    wire N__9488;
    wire N__9485;
    wire N__9482;
    wire N__9481;
    wire N__9480;
    wire N__9475;
    wire N__9472;
    wire N__9467;
    wire N__9464;
    wire N__9463;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9436;
    wire N__9435;
    wire N__9432;
    wire N__9427;
    wire N__9424;
    wire N__9419;
    wire N__9416;
    wire N__9413;
    wire N__9410;
    wire N__9407;
    wire N__9404;
    wire N__9401;
    wire N__9398;
    wire N__9397;
    wire N__9394;
    wire N__9391;
    wire N__9386;
    wire N__9383;
    wire N__9380;
    wire N__9377;
    wire N__9374;
    wire N__9371;
    wire N__9370;
    wire N__9367;
    wire N__9364;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9350;
    wire N__9347;
    wire N__9344;
    wire N__9341;
    wire N__9338;
    wire N__9335;
    wire N__9332;
    wire N__9331;
    wire N__9330;
    wire N__9329;
    wire N__9326;
    wire N__9323;
    wire N__9318;
    wire N__9311;
    wire N__9310;
    wire N__9309;
    wire N__9306;
    wire N__9301;
    wire N__9296;
    wire N__9293;
    wire N__9292;
    wire N__9291;
    wire N__9290;
    wire N__9287;
    wire N__9284;
    wire N__9279;
    wire N__9272;
    wire N__9269;
    wire N__9266;
    wire N__9265;
    wire N__9260;
    wire N__9257;
    wire N__9256;
    wire N__9253;
    wire N__9250;
    wire N__9245;
    wire N__9244;
    wire N__9241;
    wire N__9238;
    wire N__9233;
    wire N__9230;
    wire N__9227;
    wire N__9224;
    wire N__9221;
    wire N__9218;
    wire N__9215;
    wire N__9212;
    wire N__9211;
    wire N__9208;
    wire N__9205;
    wire N__9200;
    wire N__9197;
    wire N__9194;
    wire N__9193;
    wire N__9192;
    wire N__9189;
    wire N__9186;
    wire N__9185;
    wire N__9182;
    wire N__9179;
    wire N__9174;
    wire N__9171;
    wire N__9166;
    wire N__9161;
    wire N__9160;
    wire N__9159;
    wire N__9158;
    wire N__9157;
    wire N__9156;
    wire N__9155;
    wire N__9154;
    wire N__9153;
    wire N__9134;
    wire N__9131;
    wire N__9128;
    wire N__9125;
    wire N__9122;
    wire N__9121;
    wire N__9118;
    wire N__9115;
    wire N__9112;
    wire N__9109;
    wire N__9108;
    wire N__9103;
    wire N__9100;
    wire N__9097;
    wire N__9096;
    wire N__9093;
    wire N__9090;
    wire N__9087;
    wire N__9082;
    wire N__9079;
    wire N__9078;
    wire N__9075;
    wire N__9072;
    wire N__9069;
    wire N__9062;
    wire N__9059;
    wire N__9058;
    wire N__9055;
    wire N__9052;
    wire N__9049;
    wire N__9048;
    wire N__9047;
    wire N__9046;
    wire N__9045;
    wire N__9042;
    wire N__9041;
    wire N__9040;
    wire N__9037;
    wire N__9036;
    wire N__9035;
    wire N__9034;
    wire N__9031;
    wire N__9028;
    wire N__9027;
    wire N__9026;
    wire N__9025;
    wire N__9024;
    wire N__9023;
    wire N__9022;
    wire N__9021;
    wire N__9016;
    wire N__9013;
    wire N__9008;
    wire N__9007;
    wire N__9004;
    wire N__9001;
    wire N__8998;
    wire N__8985;
    wire N__8984;
    wire N__8983;
    wire N__8980;
    wire N__8977;
    wire N__8976;
    wire N__8973;
    wire N__8970;
    wire N__8969;
    wire N__8966;
    wire N__8961;
    wire N__8958;
    wire N__8949;
    wire N__8948;
    wire N__8945;
    wire N__8940;
    wire N__8937;
    wire N__8934;
    wire N__8929;
    wire N__8928;
    wire N__8925;
    wire N__8918;
    wire N__8915;
    wire N__8912;
    wire N__8901;
    wire N__8898;
    wire N__8895;
    wire N__8892;
    wire N__8887;
    wire N__8882;
    wire N__8879;
    wire N__8876;
    wire N__8871;
    wire N__8868;
    wire N__8865;
    wire N__8862;
    wire N__8857;
    wire N__8854;
    wire N__8849;
    wire N__8846;
    wire N__8843;
    wire N__8840;
    wire N__8837;
    wire N__8834;
    wire N__8833;
    wire N__8832;
    wire N__8829;
    wire N__8828;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8807;
    wire N__8806;
    wire N__8803;
    wire N__8802;
    wire N__8801;
    wire N__8800;
    wire N__8799;
    wire N__8796;
    wire N__8793;
    wire N__8788;
    wire N__8783;
    wire N__8780;
    wire N__8771;
    wire N__8768;
    wire N__8767;
    wire N__8764;
    wire N__8763;
    wire N__8762;
    wire N__8759;
    wire N__8756;
    wire N__8753;
    wire N__8750;
    wire N__8741;
    wire N__8738;
    wire N__8737;
    wire N__8736;
    wire N__8735;
    wire N__8734;
    wire N__8731;
    wire N__8730;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8705;
    wire N__8702;
    wire N__8701;
    wire N__8700;
    wire N__8697;
    wire N__8696;
    wire N__8695;
    wire N__8692;
    wire N__8689;
    wire N__8686;
    wire N__8683;
    wire N__8678;
    wire N__8675;
    wire N__8666;
    wire N__8665;
    wire N__8662;
    wire N__8661;
    wire N__8658;
    wire N__8657;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8636;
    wire N__8633;
    wire N__8632;
    wire N__8631;
    wire N__8630;
    wire N__8629;
    wire N__8626;
    wire N__8623;
    wire N__8620;
    wire N__8615;
    wire N__8606;
    wire N__8603;
    wire N__8602;
    wire N__8601;
    wire N__8600;
    wire N__8597;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8572;
    wire N__8569;
    wire N__8568;
    wire N__8565;
    wire N__8562;
    wire N__8559;
    wire N__8556;
    wire N__8549;
    wire N__8546;
    wire N__8545;
    wire N__8544;
    wire N__8541;
    wire N__8538;
    wire N__8535;
    wire N__8528;
    wire N__8525;
    wire N__8522;
    wire N__8519;
    wire N__8516;
    wire N__8513;
    wire N__8510;
    wire N__8507;
    wire N__8506;
    wire N__8503;
    wire N__8500;
    wire N__8495;
    wire N__8494;
    wire N__8491;
    wire N__8488;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8476;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8455;
    wire N__8452;
    wire N__8451;
    wire N__8448;
    wire N__8445;
    wire N__8442;
    wire N__8439;
    wire N__8436;
    wire N__8431;
    wire N__8428;
    wire N__8425;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire N__8402;
    wire N__8399;
    wire N__8396;
    wire N__8395;
    wire N__8392;
    wire N__8389;
    wire N__8384;
    wire N__8383;
    wire N__8380;
    wire N__8379;
    wire N__8376;
    wire N__8373;
    wire N__8370;
    wire N__8367;
    wire N__8364;
    wire N__8359;
    wire N__8356;
    wire N__8353;
    wire N__8350;
    wire N__8347;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8333;
    wire N__8330;
    wire N__8327;
    wire N__8324;
    wire N__8321;
    wire N__8318;
    wire N__8315;
    wire N__8314;
    wire N__8313;
    wire N__8312;
    wire N__8311;
    wire N__8304;
    wire N__8301;
    wire N__8298;
    wire N__8291;
    wire N__8290;
    wire N__8289;
    wire N__8288;
    wire N__8285;
    wire N__8282;
    wire N__8277;
    wire N__8270;
    wire N__8269;
    wire N__8268;
    wire N__8267;
    wire N__8264;
    wire N__8261;
    wire N__8258;
    wire N__8253;
    wire N__8246;
    wire N__8245;
    wire N__8244;
    wire N__8241;
    wire N__8236;
    wire N__8231;
    wire N__8230;
    wire N__8229;
    wire N__8228;
    wire N__8225;
    wire N__8220;
    wire N__8215;
    wire N__8210;
    wire N__8207;
    wire N__8206;
    wire N__8205;
    wire N__8204;
    wire N__8203;
    wire N__8200;
    wire N__8191;
    wire N__8186;
    wire N__8185;
    wire N__8184;
    wire N__8181;
    wire N__8180;
    wire N__8177;
    wire N__8170;
    wire N__8165;
    wire N__8164;
    wire N__8159;
    wire N__8156;
    wire N__8155;
    wire N__8152;
    wire N__8149;
    wire N__8146;
    wire N__8141;
    wire N__8140;
    wire N__8139;
    wire N__8134;
    wire N__8131;
    wire N__8126;
    wire N__8125;
    wire N__8124;
    wire N__8121;
    wire N__8120;
    wire N__8119;
    wire N__8118;
    wire N__8117;
    wire N__8114;
    wire N__8111;
    wire N__8108;
    wire N__8099;
    wire N__8090;
    wire N__8087;
    wire N__8086;
    wire N__8085;
    wire N__8082;
    wire N__8079;
    wire N__8076;
    wire N__8073;
    wire N__8070;
    wire N__8067;
    wire N__8062;
    wire N__8059;
    wire N__8054;
    wire N__8051;
    wire N__8048;
    wire N__8047;
    wire N__8044;
    wire N__8041;
    wire N__8036;
    wire N__8033;
    wire N__8030;
    wire N__8027;
    wire N__8024;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8012;
    wire N__8009;
    wire N__8008;
    wire N__8007;
    wire N__8004;
    wire N__8001;
    wire N__7998;
    wire N__7997;
    wire N__7994;
    wire N__7991;
    wire N__7988;
    wire N__7987;
    wire N__7984;
    wire N__7981;
    wire N__7976;
    wire N__7973;
    wire N__7964;
    wire N__7961;
    wire N__7958;
    wire N__7955;
    wire N__7952;
    wire N__7949;
    wire N__7948;
    wire N__7947;
    wire N__7946;
    wire N__7943;
    wire N__7938;
    wire N__7935;
    wire N__7928;
    wire N__7925;
    wire N__7922;
    wire N__7919;
    wire N__7916;
    wire N__7913;
    wire N__7910;
    wire N__7907;
    wire N__7904;
    wire N__7901;
    wire N__7898;
    wire N__7895;
    wire N__7892;
    wire N__7889;
    wire N__7886;
    wire N__7883;
    wire N__7880;
    wire N__7877;
    wire N__7876;
    wire N__7873;
    wire N__7870;
    wire N__7865;
    wire N__7862;
    wire N__7861;
    wire N__7860;
    wire N__7853;
    wire N__7850;
    wire N__7849;
    wire N__7848;
    wire N__7847;
    wire N__7844;
    wire N__7843;
    wire N__7840;
    wire N__7833;
    wire N__7830;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7814;
    wire N__7811;
    wire N__7808;
    wire N__7805;
    wire N__7802;
    wire N__7799;
    wire N__7796;
    wire N__7793;
    wire N__7790;
    wire N__7787;
    wire N__7786;
    wire N__7783;
    wire N__7780;
    wire N__7775;
    wire N__7772;
    wire N__7769;
    wire N__7766;
    wire N__7763;
    wire N__7760;
    wire N__7757;
    wire N__7754;
    wire N__7753;
    wire N__7752;
    wire N__7751;
    wire N__7748;
    wire N__7743;
    wire N__7740;
    wire N__7733;
    wire N__7732;
    wire N__7731;
    wire N__7728;
    wire N__7721;
    wire N__7718;
    wire N__7717;
    wire N__7714;
    wire N__7711;
    wire N__7710;
    wire N__7705;
    wire N__7704;
    wire N__7703;
    wire N__7700;
    wire N__7697;
    wire N__7694;
    wire N__7691;
    wire N__7690;
    wire N__7687;
    wire N__7680;
    wire N__7677;
    wire N__7674;
    wire N__7671;
    wire N__7668;
    wire N__7665;
    wire N__7662;
    wire N__7659;
    wire N__7656;
    wire N__7653;
    wire N__7646;
    wire N__7645;
    wire N__7642;
    wire N__7639;
    wire N__7636;
    wire N__7631;
    wire N__7628;
    wire N__7625;
    wire N__7622;
    wire N__7619;
    wire N__7616;
    wire N__7615;
    wire N__7612;
    wire N__7609;
    wire N__7606;
    wire N__7605;
    wire N__7602;
    wire N__7599;
    wire N__7596;
    wire N__7593;
    wire N__7590;
    wire N__7587;
    wire N__7586;
    wire N__7583;
    wire N__7580;
    wire N__7577;
    wire N__7574;
    wire N__7565;
    wire N__7562;
    wire N__7561;
    wire N__7558;
    wire N__7555;
    wire N__7552;
    wire N__7549;
    wire N__7544;
    wire N__7541;
    wire N__7538;
    wire N__7535;
    wire N__7532;
    wire N__7529;
    wire N__7526;
    wire N__7523;
    wire N__7520;
    wire N__7517;
    wire N__7514;
    wire N__7511;
    wire N__7508;
    wire N__7505;
    wire N__7502;
    wire N__7499;
    wire N__7496;
    wire N__7493;
    wire N__7490;
    wire N__7487;
    wire N__7486;
    wire N__7481;
    wire N__7478;
    wire N__7477;
    wire N__7474;
    wire N__7471;
    wire N__7466;
    wire N__7465;
    wire N__7460;
    wire N__7457;
    wire N__7454;
    wire N__7451;
    wire N__7448;
    wire N__7445;
    wire N__7442;
    wire N__7439;
    wire N__7436;
    wire N__7433;
    wire N__7430;
    wire N__7427;
    wire N__7424;
    wire N__7421;
    wire N__7418;
    wire N__7415;
    wire N__7412;
    wire N__7411;
    wire N__7408;
    wire N__7407;
    wire N__7406;
    wire N__7403;
    wire N__7400;
    wire N__7397;
    wire N__7394;
    wire N__7391;
    wire N__7390;
    wire N__7385;
    wire N__7382;
    wire N__7379;
    wire N__7376;
    wire N__7371;
    wire N__7368;
    wire N__7365;
    wire N__7362;
    wire N__7355;
    wire N__7352;
    wire N__7351;
    wire N__7348;
    wire N__7345;
    wire N__7340;
    wire N__7339;
    wire N__7338;
    wire N__7337;
    wire N__7334;
    wire N__7333;
    wire N__7332;
    wire N__7329;
    wire N__7326;
    wire N__7325;
    wire N__7324;
    wire N__7323;
    wire N__7322;
    wire N__7321;
    wire N__7320;
    wire N__7317;
    wire N__7316;
    wire N__7315;
    wire N__7314;
    wire N__7313;
    wire N__7308;
    wire N__7305;
    wire N__7300;
    wire N__7297;
    wire N__7294;
    wire N__7291;
    wire N__7288;
    wire N__7285;
    wire N__7282;
    wire N__7275;
    wire N__7272;
    wire N__7269;
    wire N__7266;
    wire N__7263;
    wire N__7250;
    wire N__7247;
    wire N__7240;
    wire N__7235;
    wire N__7232;
    wire N__7227;
    wire N__7220;
    wire N__7217;
    wire N__7214;
    wire N__7211;
    wire N__7208;
    wire N__7205;
    wire N__7202;
    wire N__7199;
    wire N__7196;
    wire N__7193;
    wire N__7190;
    wire N__7187;
    wire N__7184;
    wire N__7183;
    wire N__7180;
    wire N__7175;
    wire N__7174;
    wire N__7171;
    wire N__7168;
    wire N__7163;
    wire N__7160;
    wire N__7157;
    wire N__7154;
    wire N__7151;
    wire N__7148;
    wire N__7145;
    wire N__7142;
    wire N__7139;
    wire N__7138;
    wire N__7137;
    wire N__7134;
    wire N__7129;
    wire N__7124;
    wire N__7121;
    wire N__7118;
    wire N__7117;
    wire N__7114;
    wire N__7111;
    wire N__7108;
    wire N__7105;
    wire N__7100;
    wire N__7099;
    wire N__7096;
    wire N__7095;
    wire N__7094;
    wire N__7093;
    wire N__7090;
    wire N__7089;
    wire N__7088;
    wire N__7085;
    wire N__7082;
    wire N__7077;
    wire N__7074;
    wire N__7069;
    wire N__7064;
    wire N__7055;
    wire N__7052;
    wire N__7049;
    wire N__7046;
    wire N__7045;
    wire N__7044;
    wire N__7041;
    wire N__7040;
    wire N__7037;
    wire N__7032;
    wire N__7029;
    wire N__7022;
    wire N__7019;
    wire N__7016;
    wire N__7013;
    wire N__7010;
    wire N__7007;
    wire N__7004;
    wire N__7001;
    wire N__6998;
    wire N__6995;
    wire N__6994;
    wire N__6991;
    wire N__6988;
    wire N__6987;
    wire N__6986;
    wire N__6985;
    wire N__6984;
    wire N__6983;
    wire N__6982;
    wire N__6981;
    wire N__6976;
    wire N__6971;
    wire N__6966;
    wire N__6963;
    wire N__6958;
    wire N__6947;
    wire N__6944;
    wire N__6941;
    wire N__6940;
    wire N__6939;
    wire N__6938;
    wire N__6937;
    wire N__6936;
    wire N__6935;
    wire N__6932;
    wire N__6929;
    wire N__6928;
    wire N__6925;
    wire N__6924;
    wire N__6921;
    wire N__6916;
    wire N__6913;
    wire N__6906;
    wire N__6903;
    wire N__6902;
    wire N__6899;
    wire N__6896;
    wire N__6893;
    wire N__6890;
    wire N__6885;
    wire N__6880;
    wire N__6879;
    wire N__6876;
    wire N__6871;
    wire N__6866;
    wire N__6863;
    wire N__6854;
    wire N__6853;
    wire N__6852;
    wire N__6849;
    wire N__6848;
    wire N__6847;
    wire N__6846;
    wire N__6843;
    wire N__6842;
    wire N__6839;
    wire N__6836;
    wire N__6831;
    wire N__6828;
    wire N__6825;
    wire N__6822;
    wire N__6809;
    wire N__6808;
    wire N__6805;
    wire N__6802;
    wire N__6797;
    wire N__6794;
    wire N__6791;
    wire N__6788;
    wire N__6785;
    wire N__6782;
    wire N__6779;
    wire N__6776;
    wire N__6773;
    wire N__6770;
    wire N__6767;
    wire N__6764;
    wire N__6761;
    wire N__6758;
    wire N__6755;
    wire N__6752;
    wire N__6751;
    wire N__6748;
    wire N__6743;
    wire N__6740;
    wire N__6737;
    wire N__6734;
    wire N__6731;
    wire N__6728;
    wire N__6725;
    wire N__6722;
    wire N__6719;
    wire N__6718;
    wire N__6713;
    wire N__6712;
    wire N__6709;
    wire N__6706;
    wire N__6705;
    wire N__6704;
    wire N__6701;
    wire N__6698;
    wire N__6693;
    wire N__6686;
    wire N__6685;
    wire N__6684;
    wire N__6679;
    wire N__6676;
    wire N__6675;
    wire N__6674;
    wire N__6673;
    wire N__6672;
    wire N__6671;
    wire N__6670;
    wire N__6665;
    wire N__6660;
    wire N__6657;
    wire N__6656;
    wire N__6655;
    wire N__6652;
    wire N__6649;
    wire N__6646;
    wire N__6641;
    wire N__6636;
    wire N__6633;
    wire N__6632;
    wire N__6627;
    wire N__6620;
    wire N__6617;
    wire N__6614;
    wire N__6611;
    wire N__6604;
    wire N__6601;
    wire N__6598;
    wire N__6593;
    wire N__6590;
    wire N__6587;
    wire N__6584;
    wire N__6581;
    wire N__6578;
    wire N__6575;
    wire N__6572;
    wire N__6569;
    wire N__6566;
    wire N__6563;
    wire N__6560;
    wire N__6557;
    wire N__6554;
    wire N__6553;
    wire N__6550;
    wire N__6547;
    wire N__6544;
    wire N__6541;
    wire N__6536;
    wire N__6533;
    wire N__6532;
    wire N__6527;
    wire N__6524;
    wire N__6521;
    wire N__6520;
    wire N__6515;
    wire N__6514;
    wire N__6513;
    wire N__6512;
    wire N__6511;
    wire N__6508;
    wire N__6505;
    wire N__6502;
    wire N__6497;
    wire N__6496;
    wire N__6495;
    wire N__6492;
    wire N__6489;
    wire N__6486;
    wire N__6483;
    wire N__6480;
    wire N__6477;
    wire N__6464;
    wire N__6463;
    wire N__6462;
    wire N__6461;
    wire N__6458;
    wire N__6457;
    wire N__6456;
    wire N__6455;
    wire N__6452;
    wire N__6451;
    wire N__6450;
    wire N__6449;
    wire N__6446;
    wire N__6445;
    wire N__6442;
    wire N__6439;
    wire N__6436;
    wire N__6433;
    wire N__6428;
    wire N__6425;
    wire N__6422;
    wire N__6417;
    wire N__6412;
    wire N__6411;
    wire N__6410;
    wire N__6401;
    wire N__6396;
    wire N__6391;
    wire N__6386;
    wire N__6383;
    wire N__6380;
    wire N__6375;
    wire N__6372;
    wire N__6369;
    wire N__6362;
    wire N__6359;
    wire N__6356;
    wire N__6353;
    wire N__6350;
    wire N__6347;
    wire N__6344;
    wire N__6341;
    wire N__6338;
    wire N__6335;
    wire N__6332;
    wire N__6329;
    wire N__6326;
    wire N__6323;
    wire N__6320;
    wire N__6317;
    wire N__6314;
    wire N__6311;
    wire N__6308;
    wire N__6307;
    wire N__6302;
    wire N__6299;
    wire N__6296;
    wire N__6293;
    wire N__6290;
    wire N__6287;
    wire N__6284;
    wire N__6283;
    wire N__6280;
    wire N__6277;
    wire N__6272;
    wire N__6269;
    wire N__6268;
    wire N__6267;
    wire N__6266;
    wire N__6263;
    wire N__6260;
    wire N__6257;
    wire N__6254;
    wire N__6253;
    wire N__6248;
    wire N__6247;
    wire N__6246;
    wire N__6245;
    wire N__6244;
    wire N__6239;
    wire N__6238;
    wire N__6235;
    wire N__6232;
    wire N__6225;
    wire N__6222;
    wire N__6219;
    wire N__6216;
    wire N__6203;
    wire N__6200;
    wire N__6197;
    wire N__6194;
    wire N__6191;
    wire N__6188;
    wire N__6185;
    wire N__6184;
    wire N__6183;
    wire N__6180;
    wire N__6177;
    wire N__6174;
    wire N__6171;
    wire N__6166;
    wire N__6163;
    wire N__6160;
    wire N__6157;
    wire N__6152;
    wire N__6149;
    wire N__6146;
    wire N__6143;
    wire N__6140;
    wire N__6139;
    wire N__6138;
    wire N__6137;
    wire N__6136;
    wire N__6135;
    wire N__6132;
    wire N__6131;
    wire N__6128;
    wire N__6121;
    wire N__6118;
    wire N__6117;
    wire N__6114;
    wire N__6111;
    wire N__6106;
    wire N__6101;
    wire N__6098;
    wire N__6095;
    wire N__6090;
    wire N__6085;
    wire N__6082;
    wire N__6079;
    wire N__6076;
    wire N__6071;
    wire N__6068;
    wire N__6065;
    wire N__6062;
    wire N__6059;
    wire N__6056;
    wire N__6053;
    wire N__6050;
    wire N__6049;
    wire N__6048;
    wire N__6047;
    wire N__6044;
    wire N__6043;
    wire N__6042;
    wire N__6039;
    wire N__6036;
    wire N__6033;
    wire N__6030;
    wire N__6025;
    wire N__6022;
    wire N__6011;
    wire N__6010;
    wire N__6009;
    wire N__6002;
    wire N__6001;
    wire N__6000;
    wire N__5999;
    wire N__5996;
    wire N__5993;
    wire N__5990;
    wire N__5989;
    wire N__5986;
    wire N__5985;
    wire N__5984;
    wire N__5983;
    wire N__5982;
    wire N__5981;
    wire N__5976;
    wire N__5971;
    wire N__5968;
    wire N__5965;
    wire N__5962;
    wire N__5959;
    wire N__5954;
    wire N__5949;
    wire N__5938;
    wire N__5935;
    wire N__5932;
    wire N__5929;
    wire N__5926;
    wire N__5923;
    wire N__5920;
    wire N__5915;
    wire N__5912;
    wire N__5909;
    wire N__5906;
    wire N__5905;
    wire N__5902;
    wire N__5899;
    wire N__5894;
    wire N__5891;
    wire N__5888;
    wire N__5885;
    wire N__5882;
    wire N__5879;
    wire N__5876;
    wire N__5873;
    wire N__5870;
    wire N__5867;
    wire N__5864;
    wire N__5861;
    wire N__5860;
    wire N__5857;
    wire N__5854;
    wire N__5849;
    wire N__5846;
    wire N__5843;
    wire N__5840;
    wire N__5837;
    wire N__5834;
    wire N__5831;
    wire N__5828;
    wire N__5825;
    wire N__5822;
    wire N__5821;
    wire N__5818;
    wire N__5815;
    wire N__5810;
    wire N__5807;
    wire N__5804;
    wire N__5801;
    wire N__5798;
    wire N__5797;
    wire N__5792;
    wire N__5789;
    wire N__5786;
    wire N__5783;
    wire N__5782;
    wire N__5781;
    wire N__5780;
    wire N__5779;
    wire N__5776;
    wire N__5773;
    wire N__5770;
    wire N__5769;
    wire N__5766;
    wire N__5763;
    wire N__5762;
    wire N__5757;
    wire N__5750;
    wire N__5749;
    wire N__5746;
    wire N__5743;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5729;
    wire N__5720;
    wire N__5719;
    wire N__5718;
    wire N__5713;
    wire N__5712;
    wire N__5711;
    wire N__5710;
    wire N__5709;
    wire N__5706;
    wire N__5703;
    wire N__5698;
    wire N__5697;
    wire N__5694;
    wire N__5691;
    wire N__5684;
    wire N__5681;
    wire N__5672;
    wire N__5669;
    wire N__5668;
    wire N__5667;
    wire N__5666;
    wire N__5665;
    wire N__5658;
    wire N__5655;
    wire N__5652;
    wire N__5649;
    wire N__5642;
    wire N__5639;
    wire N__5636;
    wire N__5633;
    wire N__5632;
    wire N__5631;
    wire N__5628;
    wire N__5625;
    wire N__5624;
    wire N__5623;
    wire N__5620;
    wire N__5619;
    wire N__5618;
    wire N__5617;
    wire N__5614;
    wire N__5609;
    wire N__5604;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5594;
    wire N__5587;
    wire N__5584;
    wire N__5583;
    wire N__5576;
    wire N__5571;
    wire N__5568;
    wire N__5565;
    wire N__5560;
    wire N__5557;
    wire N__5554;
    wire N__5549;
    wire N__5546;
    wire N__5545;
    wire N__5542;
    wire N__5541;
    wire N__5540;
    wire N__5537;
    wire N__5536;
    wire N__5533;
    wire N__5530;
    wire N__5527;
    wire N__5524;
    wire N__5521;
    wire N__5520;
    wire N__5519;
    wire N__5512;
    wire N__5507;
    wire N__5504;
    wire N__5501;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5489;
    wire N__5482;
    wire N__5479;
    wire N__5474;
    wire N__5471;
    wire N__5468;
    wire N__5465;
    wire N__5462;
    wire N__5459;
    wire N__5456;
    wire N__5453;
    wire N__5450;
    wire N__5447;
    wire N__5444;
    wire N__5441;
    wire N__5438;
    wire N__5435;
    wire N__5434;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5411;
    wire N__5410;
    wire N__5409;
    wire N__5408;
    wire N__5407;
    wire N__5404;
    wire N__5399;
    wire N__5396;
    wire N__5393;
    wire N__5384;
    wire N__5381;
    wire N__5378;
    wire N__5375;
    wire N__5372;
    wire N__5371;
    wire N__5370;
    wire N__5369;
    wire N__5368;
    wire N__5365;
    wire N__5360;
    wire N__5359;
    wire N__5356;
    wire N__5353;
    wire N__5348;
    wire N__5345;
    wire N__5340;
    wire N__5337;
    wire N__5334;
    wire N__5331;
    wire N__5324;
    wire N__5321;
    wire N__5318;
    wire N__5315;
    wire N__5314;
    wire N__5309;
    wire N__5306;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5294;
    wire N__5291;
    wire N__5290;
    wire N__5287;
    wire N__5284;
    wire N__5281;
    wire N__5278;
    wire N__5273;
    wire N__5270;
    wire N__5267;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5255;
    wire N__5252;
    wire N__5249;
    wire N__5246;
    wire N__5243;
    wire N__5240;
    wire N__5237;
    wire N__5234;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5222;
    wire N__5219;
    wire N__5216;
    wire N__5213;
    wire N__5210;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5198;
    wire N__5195;
    wire N__5192;
    wire N__5191;
    wire N__5188;
    wire N__5187;
    wire N__5186;
    wire N__5183;
    wire N__5180;
    wire N__5177;
    wire N__5174;
    wire N__5169;
    wire N__5164;
    wire N__5161;
    wire N__5156;
    wire N__5153;
    wire N__5150;
    wire N__5149;
    wire N__5146;
    wire N__5143;
    wire N__5138;
    wire N__5137;
    wire N__5134;
    wire N__5131;
    wire N__5128;
    wire N__5127;
    wire N__5126;
    wire N__5125;
    wire N__5122;
    wire N__5119;
    wire N__5116;
    wire N__5113;
    wire N__5110;
    wire N__5107;
    wire N__5100;
    wire N__5093;
    wire N__5090;
    wire N__5087;
    wire N__5086;
    wire N__5083;
    wire N__5080;
    wire N__5075;
    wire N__5072;
    wire N__5069;
    wire N__5066;
    wire N__5063;
    wire N__5060;
    wire N__5059;
    wire N__5058;
    wire N__5051;
    wire N__5048;
    wire N__5045;
    wire N__5044;
    wire N__5043;
    wire N__5036;
    wire N__5033;
    wire N__5030;
    wire N__5029;
    wire N__5028;
    wire N__5025;
    wire N__5024;
    wire N__5021;
    wire N__5018;
    wire N__5015;
    wire N__5012;
    wire N__5007;
    wire N__5004;
    wire N__5001;
    wire N__4994;
    wire N__4991;
    wire N__4990;
    wire N__4987;
    wire N__4984;
    wire N__4981;
    wire N__4978;
    wire N__4977;
    wire N__4976;
    wire N__4975;
    wire N__4974;
    wire N__4973;
    wire N__4968;
    wire N__4961;
    wire N__4956;
    wire N__4949;
    wire N__4946;
    wire N__4945;
    wire N__4942;
    wire N__4939;
    wire N__4938;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4928;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4916;
    wire N__4907;
    wire N__4904;
    wire N__4903;
    wire N__4902;
    wire N__4901;
    wire N__4900;
    wire N__4899;
    wire N__4894;
    wire N__4889;
    wire N__4884;
    wire N__4879;
    wire N__4876;
    wire N__4873;
    wire N__4870;
    wire N__4867;
    wire N__4864;
    wire N__4859;
    wire N__4858;
    wire N__4857;
    wire N__4854;
    wire N__4849;
    wire N__4844;
    wire N__4841;
    wire N__4838;
    wire N__4835;
    wire N__4832;
    wire N__4831;
    wire N__4828;
    wire N__4825;
    wire N__4822;
    wire N__4819;
    wire N__4816;
    wire N__4815;
    wire N__4814;
    wire N__4811;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4799;
    wire N__4792;
    wire N__4789;
    wire N__4786;
    wire N__4781;
    wire N__4778;
    wire N__4777;
    wire N__4774;
    wire N__4771;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4753;
    wire N__4752;
    wire N__4749;
    wire N__4746;
    wire N__4743;
    wire N__4742;
    wire N__4739;
    wire N__4734;
    wire N__4731;
    wire N__4728;
    wire N__4725;
    wire N__4722;
    wire N__4717;
    wire N__4714;
    wire N__4709;
    wire N__4706;
    wire N__4703;
    wire N__4700;
    wire N__4697;
    wire N__4694;
    wire N__4693;
    wire N__4690;
    wire N__4687;
    wire N__4682;
    wire N__4681;
    wire N__4678;
    wire N__4675;
    wire N__4670;
    wire N__4667;
    wire N__4664;
    wire N__4661;
    wire N__4658;
    wire N__4655;
    wire N__4652;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4642;
    wire N__4637;
    wire N__4634;
    wire N__4631;
    wire N__4628;
    wire N__4625;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4613;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4603;
    wire N__4602;
    wire N__4601;
    wire N__4600;
    wire N__4597;
    wire N__4594;
    wire N__4589;
    wire N__4586;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4565;
    wire N__4562;
    wire N__4559;
    wire N__4556;
    wire N__4553;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4541;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4523;
    wire N__4520;
    wire N__4517;
    wire N__4514;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4502;
    wire N__4499;
    wire N__4498;
    wire N__4495;
    wire N__4492;
    wire N__4487;
    wire N__4484;
    wire N__4483;
    wire N__4480;
    wire N__4477;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4463;
    wire N__4460;
    wire N__4457;
    wire N__4456;
    wire N__4453;
    wire N__4450;
    wire N__4445;
    wire N__4442;
    wire N__4439;
    wire N__4436;
    wire N__4433;
    wire N__4430;
    wire N__4429;
    wire N__4424;
    wire N__4421;
    wire N__4418;
    wire N__4415;
    wire N__4412;
    wire N__4411;
    wire N__4406;
    wire N__4403;
    wire N__4400;
    wire N__4397;
    wire N__4394;
    wire N__4393;
    wire N__4390;
    wire N__4385;
    wire N__4382;
    wire N__4379;
    wire N__4376;
    wire N__4373;
    wire N__4372;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4346;
    wire N__4343;
    wire N__4340;
    wire N__4337;
    wire N__4334;
    wire N__4331;
    wire N__4328;
    wire N__4325;
    wire N__4322;
    wire N__4319;
    wire N__4316;
    wire N__4313;
    wire N__4310;
    wire N__4307;
    wire N__4304;
    wire N__4301;
    wire N__4298;
    wire N__4297;
    wire N__4294;
    wire N__4291;
    wire N__4286;
    wire N__4283;
    wire N__4280;
    wire N__4277;
    wire N__4274;
    wire N__4273;
    wire N__4270;
    wire N__4267;
    wire N__4262;
    wire N__4259;
    wire N__4256;
    wire N__4253;
    wire N__4250;
    wire N__4247;
    wire N__4244;
    wire N__4241;
    wire N__4238;
    wire N__4235;
    wire PPIO_c;
    wire GNDG0;
    wire SPIO_c;
    wire VCCG0;
    wire A_c_26;
    wire A_c_27;
    wire \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_5_cascade_ ;
    wire A_c_25;
    wire A_c_24;
    wire \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4 ;
    wire A_c_29;
    wire A_c_31;
    wire A_c_30;
    wire A_c_28;
    wire U409_ADDRESS_DECODE_un1_RTC_ENn_i;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0 ;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0_cascade_ ;
    wire \U409_ADDRESS_DECODE.HIROMZ0Z_0_cascade_ ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0Z0Z_0 ;
    wire \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7 ;
    wire TT_c_1;
    wire TT_c_0;
    wire \INVU409_AUTOCONFIG.LIDE_BASE_3C_net ;
    wire LIDE_BASE_6;
    wire \U409_AUTOCONFIG.N_99_cascade_ ;
    wire LIDE_BASE_5;
    wire \INVU409_AUTOCONFIG.LIDE_BASE_5C_net ;
    wire D_in_4;
    wire \U409_AUTOCONFIG.N_101 ;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2_cascade_ ;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4 ;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2 ;
    wire U409_ADDRESS_DECODE_un1_REGSPACEn_i;
    wire \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_5 ;
    wire \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_0Z0Z_3_cascade_ ;
    wire \U409_ADDRESS_DECODE.HIROMZ0Z_0 ;
    wire \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_0 ;
    wire \U409_AUTOCONFIG.N_121_cascade_ ;
    wire A_c_7;
    wire A_c_6;
    wire A_c_5;
    wire A_c_3;
    wire \U409_AUTOCONFIG.N_121 ;
    wire \U409_AUTOCONFIG.N_123 ;
    wire A_c_16;
    wire A_c_15;
    wire D_1_i;
    wire \U409_AUTOCONFIG.N_103 ;
    wire LIDE_BASE_4;
    wire LIDE_BASE_3;
    wire \INVU409_AUTOCONFIG.LIDE_BASE_1C_net ;
    wire D_in_7;
    wire \U409_ADDRESS_DECODE.PORTSIZEZ0Z_1 ;
    wire \U409_ADDRESS_DECODE.PORTSIZEZ0Z_0_cascade_ ;
    wire PORTSIZE_0_i;
    wire BUFENn_c;
    wire U409_ADDRESS_DECODE_un1_ATA_ENn_i;
    wire A_c_18;
    wire LIDE_BASE_2;
    wire A_c_17;
    wire LIDE_BASE_1;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3 ;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1_cascade_ ;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2 ;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0 ;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_ ;
    wire \U409_ADDRESS_DECODE.ATA_ENZ0 ;
    wire \U409_AUTOCONFIG.PR_OUT_cnst_i_i_0_0_2 ;
    wire \INVU409_AUTOCONFIG.PR_OUT_2C_net ;
    wire \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_1_cascade_ ;
    wire A_c_19;
    wire \U409_AUTOCONFIG.N_84 ;
    wire \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net ;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ;
    wire \U409_ADDRESS_DECODE.LOWROMZ0Z_3 ;
    wire A_c_21;
    wire A_c_20;
    wire \U409_AUTOCONFIG.PR_OUTZ0Z_2 ;
    wire D_OUT_2;
    wire \U409_AUTOCONFIG.N_97 ;
    wire \U409_AUTOCONFIG.STATE_d_2_cascade_ ;
    wire D_in_6;
    wire \U409_AUTOCONFIG.N_105 ;
    wire \U409_AUTOCONFIG.N_49 ;
    wire D_in_5;
    wire \U409_AUTOCONFIG.N_49_cascade_ ;
    wire \U409_AUTOCONFIG.N_107 ;
    wire \U409_AUTOCONFIG.N_95 ;
    wire \U409_AUTOCONFIG.N_48_cascade_ ;
    wire \U409_AUTOCONFIG.un1_A_13 ;
    wire \U409_AUTOCONFIG.STATE_d_2 ;
    wire \INVU409_AUTOCONFIG.LIDE_BASE_7C_net ;
    wire LIDE_BASE_7;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_4 ;
    wire \U409_AUTOCONFIG.un1_STATE_6_0 ;
    wire \U409_AUTOCONFIG.N_48 ;
    wire \U409_AUTOCONFIG.LIDE_CONFZ0 ;
    wire \INVU409_AUTOCONFIG.STATE_0C_net ;
    wire \U409_AUTOCONFIG.STATE_ns_1_cascade_ ;
    wire A_c_22;
    wire \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_1 ;
    wire OVL_c;
    wire A_c_23;
    wire U409_ADDRESS_DECODE_un1_RAMSPACEn_i;
    wire \U409_AUTOCONFIG.STATEZ0Z_1 ;
    wire RnW_c;
    wire CPUCONFn_c;
    wire \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_a3_1_cascade_ ;
    wire \U409_AUTOCONFIG.N_227_3_cascade_ ;
    wire \INVU409_AUTOCONFIG.LIDE_OUT_2C_net ;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2 ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ;
    wire \U409_AUTOCONFIG.LIDE_OUT_RNI9FMPZ0Z_2 ;
    wire \U409_AUTOCONFIG.N_129 ;
    wire \U409_AUTOCONFIG.N_133_cascade_ ;
    wire \U409_AUTOCONFIG.N_127 ;
    wire \U409_AUTOCONFIG.N_110 ;
    wire A_c_4;
    wire D_OUT_1;
    wire \U409_AUTOCONFIG.LIDE_OUT_RNIBHMPZ0Z_3 ;
    wire D_OUT_3;
    wire \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa ;
    wire CONFIGENn_c;
    wire \INVU409_AUTOCONFIG.CONFIGUREDC_net ;
    wire \U409_AUTOCONFIG.N_4 ;
    wire D_OUT_0;
    wire \U409_AUTOCONFIG.LIDE_OUT_RNI7DMPZ0Z_1 ;
    wire \U409_AUTOCONFIG.BRIDGE_CONFZ0 ;
    wire \U409_AUTOCONFIG.LIDE_OUT_RNI5BMPZ0Z_0 ;
    wire AUTOCONFIG_SPACE;
    wire CONFIGURED;
    wire \U409_AUTOCONFIG.AC_STARTZ0 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0 ;
    wire \U409_AUTOCONFIG.N_82 ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ;
    wire \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_0Z0Z_3 ;
    wire \U409_AUTOCONFIG.PR_OUTZ0Z_3 ;
    wire \U409_AUTOCONFIG.N_131 ;
    wire \U409_AUTOCONFIG.N_93 ;
    wire \U409_AUTOCONFIG.PR_OUTZ0Z_1 ;
    wire \U409_AUTOCONFIG.N_116 ;
    wire A_c_2;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1 ;
    wire \U409_AUTOCONFIG.N_78 ;
    wire \U409_AUTOCONFIG.N_92 ;
    wire \U409_AUTOCONFIG.PR_OUTZ0Z_0 ;
    wire \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ;
    wire \U409_AUTOCONFIG.LIDE_OUT_7_i_a3_1_0 ;
    wire \U409_AUTOCONFIG.LIDE_OUT_7_i_a3_0_0 ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_0 ;
    wire \INVU409_AUTOCONFIG.LIDE_OUT_0C_net ;
    wire \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i ;
    wire \U409_AUTOCONFIG.N_133 ;
    wire A_c_1;
    wire AUTOBOOT_c;
    wire \U409_AUTOCONFIG.N_126 ;
    wire \U409_AUTOCONFIG.LIDE_OUT_7_i_1_0 ;
    wire TACKn_in;
    wire U409_ADDRESS_DECODE_un1_REGSPACEn;
    wire U409_ADDRESS_DECODE_un1_RAMSPACEn;
    wire \U409_AUTOCONFIG.STATEZ0Z_0 ;
    wire \INVU409_AUTOCONFIG.AC_TACK_nesrC_net ;
    wire \U409_AUTOCONFIG.STATE_ns_0_0_1 ;
    wire \U409_CIA.CIA_CLK_COUNT11_2_0_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ;
    wire \U409_TRANSFER_ACK.TACK_EN8 ;
    wire \U409_TRANSFER_ACK.TACK_STATE_ns_1_0 ;
    wire \U409_TRANSFER_ACK.TACK_STATEZ0Z_0 ;
    wire \U409_TRANSFER_ACK.TACK_STATEZ0Z_1 ;
    wire U409_ADDRESS_DECODE_Z2_SPACE;
    wire U409_ADDRESS_DECODE_HIROM;
    wire TACK_OUT;
    wire U409_ADDRESS_DECODE_LOWROM;
    wire U409_TRANSFER_ACK_un1_TACK_OUT_0_i;
    wire GB_BUFFER_CLK40_IN_c_g_THRU_CO;
    wire bfn_12_6_0_;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_1 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_3 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_5 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_6 ;
    wire \U409_CIA.CIA_CLK_COUNT11_2_0 ;
    wire \U409_CIA.CIA_CLK_COUNT11_3 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ;
    wire \U409_CIA.CLK_CIA6_4 ;
    wire \U409_CIA.un1_CIA_CLK_COUNT_3_2_cascade_ ;
    wire CIA_SPACE;
    wire \U409_CIA.VMA_RNOZ0Z_0_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ;
    wire U409_ADDRESS_DECODE_un1_RTC_ENn;
    wire U409_ADDRESS_DECODE_AUTOVECTOR_10;
    wire TSn_c;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_2_cascade_ ;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_5 ;
    wire \U409_ADDRESS_DECODE.AUTOVECTOR_4Z0Z_0 ;
    wire \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8 ;
    wire U409_ADDRESS_DECODE_AUTOVECTOR_11;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_2 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_cascade_ ;
    wire \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ;
    wire RESETn_c_i;
    wire A_c_12;
    wire U409_ADDRESS_DECODE_un1_CIACS0n_i;
    wire CIA_ENABLE;
    wire A_c_13;
    wire U409_ADDRESS_DECODE_un1_CIACS1n_i;
    wire \U409_TRANSFER_ACK.N_5_0 ;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_1C_net ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ;
    wire \U409_CIA.VMAZ0 ;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_0C_net ;
    wire bfn_13_8_0_;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_0 ;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_1 ;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_2 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_2 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_1 ;
    wire \U409_TRANSFER_ACK.CIA_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_3 ;
    wire AC_TACK;
    wire \U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.TACK_START_2_1 ;
    wire \U409_TRANSFER_ACK.TACK_STARTZ0 ;
    wire CLK80_OUT;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_0 ;
    wire TACK_EN;
    wire RESETn_c;
    wire \U409_TRANSFER_ACK.TACK_RST_0_i ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_6 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_0 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_7 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_1 ;
    wire \U409_CIA.CLK_CIA6_3_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_5 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_4 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_3 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_2 ;
    wire \U409_CIA.CLK_CIA_r_1_0 ;
    wire \U409_TRANSFER_ACK.N_17_mux ;
    wire \U409_TRANSFER_ACK.N_17_mux_cascade_ ;
    wire \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0 ;
    wire \U409_TRANSFER_ACK.N_3_0 ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ;
    wire \U409_TRANSFER_ACK.N_3_0_cascade_ ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0 ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.LASTCLK_1C_net ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.N_7_cascade_ ;
    wire ROM_DELAY_c_0;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ;
    wire ROM_DELAY_c_1;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.N_19_mux ;
    wire TICK60_c;
    wire \U409_TICK.TICK603_9_cascade_ ;
    wire TICK50_c;
    wire \U409_TICK.TICK603_8_cascade_ ;
    wire \U409_TICK.TICK603_14_cascade_ ;
    wire \U409_TICK.COUNTER50Z0Z_1 ;
    wire bfn_15_6_0_;
    wire \U409_TICK.COUNTER50Z0Z_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_1 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_3 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_4 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_6 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_5 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_6 ;
    wire \U409_TICK.COUNTER50Z0Z_8 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_8 ;
    wire bfn_15_7_0_;
    wire \U409_TICK.un2_COUNTER50_1_cry_9 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_10 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_11 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_12 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_13 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_15 ;
    wire \U409_TICK.COUNTER50Z0Z_16 ;
    wire CLK_CIA_c;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_0 ;
    wire \INVU409_TRANSFER_ACK.LASTCLK_0C_net ;
    wire \U409_TRANSFER_ACK.N_11 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_1 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z5 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_0 ;
    wire ROMENn_c;
    wire CLK40_IN_c_g;
    wire RESETn_c_i_g;
    wire \U409_TICK.TICK603_11 ;
    wire \U409_TICK.TICK603_10 ;
    wire \U409_TICK.TICK603_14 ;
    wire \U409_TICK.TICK603_9 ;
    wire \U409_TICK.TICK603_10_cascade_ ;
    wire \U409_TICK.COUNTER50Z0Z_3 ;
    wire \U409_TICK.TICK503_11 ;
    wire \U409_TICK.COUNTER50Z0Z_12 ;
    wire \U409_TICK.TICK503_8_cascade_ ;
    wire \U409_TICK.COUNTER50Z0Z_10 ;
    wire \U409_TICK.TICK503_14_cascade_ ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_9 ;
    wire \U409_TICK.COUNTER50Z0Z_0 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_11 ;
    wire \U409_TICK.COUNTER50Z0Z_11 ;
    wire \U409_TICK.COUNTER50Z0Z_9 ;
    wire \U409_TICK.COUNTER50Z0Z_6 ;
    wire \U409_TICK.TICK503_9_cascade_ ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_14 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_5 ;
    wire \U409_TICK.COUNTER50Z0Z_5 ;
    wire \U409_TICK.COUNTER50Z0Z_7 ;
    wire \U409_TICK.COUNTER50Z0Z_4 ;
    wire \U409_TICK.COUNTER50Z0Z_14 ;
    wire \U409_TICK.TICK503_10_cascade_ ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_15 ;
    wire \U409_TICK.COUNTER50Z0Z_15 ;
    wire \U409_TICK.COUNTER60Z0Z_1 ;
    wire \U409_TICK.COUNTER60Z0Z_0 ;
    wire bfn_17_5_0_;
    wire \U409_TICK.COUNTER60Z0Z_2 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_1 ;
    wire \U409_TICK.COUNTER60Z0Z_3 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_2 ;
    wire \U409_TICK.COUNTER60Z0Z_4 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_4 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_3 ;
    wire \U409_TICK.COUNTER60Z0Z_5 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_4 ;
    wire \U409_TICK.COUNTER60Z0Z_6 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_6 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_5 ;
    wire \U409_TICK.COUNTER60Z0Z_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_6 ;
    wire \U409_TICK.COUNTER60Z0Z_8 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_8 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_8 ;
    wire \U409_TICK.COUNTER60Z0Z_9 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_9 ;
    wire bfn_17_6_0_;
    wire \U409_TICK.COUNTER60Z0Z_10 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_9 ;
    wire \U409_TICK.COUNTER60Z0Z_11 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_10 ;
    wire \U409_TICK.COUNTER60Z0Z_12 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_11 ;
    wire \U409_TICK.COUNTER60Z0Z_13 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_12 ;
    wire \U409_TICK.COUNTER60Z0Z_14 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_13 ;
    wire \U409_TICK.COUNTER60Z0Z_15 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_15 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_15 ;
    wire \U409_TICK.COUNTER60Z0Z_16 ;
    wire \U409_TICK.TICK503_9 ;
    wire \U409_TICK.TICK503_14 ;
    wire \U409_TICK.TICK503_10 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_13 ;
    wire \U409_TICK.COUNTER50Z0Z_13 ;
    wire CLK6_c_g;
    wire PCS1_c;
    wire SCS0_c;
    wire \U409_ADDRESS_DECODE.CSZ0Z0 ;
    wire PCS0_c;
    wire A_c_14;
    wire \U409_ADDRESS_DECODE.CSZ0Z1 ;
    wire SCS1_c;
    wire CONSTANT_ONE_NET;
    wire CLK28_IN_c_g;
    wire XCLK_c;
    wire XCLK_ENn_c;
    wire AGNUS_CLK_c;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="SIMPLE";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0001111;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE pll (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__7523),
            .RESETB(N__11186),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(CLK80_OUT));
    PRE_IO_GBUF CLK6_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__11846),
            .GLOBALBUFFEROUTPUT(CLK6_c_g));
    IO_PAD CLK6_ibuf_gb_io_iopad (
            .OE(N__11848),
            .DIN(N__11847),
            .DOUT(N__11846),
            .PACKAGEPIN(CLK6));
    defparam CLK6_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK6_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK6_ibuf_gb_io_preio (
            .PADOEN(N__11848),
            .PADOUT(N__11847),
            .PADIN(N__11846),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK40_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__11836),
            .GLOBALBUFFEROUTPUT(CLK40_IN_c_g));
    IO_PAD CLK40_IN_ibuf_gb_io_iopad (
            .OE(N__11838),
            .DIN(N__11837),
            .DOUT(N__11836),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_gb_io_preio (
            .PADOEN(N__11838),
            .PADOUT(N__11837),
            .PADIN(N__11836),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK28_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__11826),
            .GLOBALBUFFEROUTPUT(CLK28_IN_c_g));
    IO_PAD CLK28_IN_ibuf_gb_io_iopad (
            .OE(N__11828),
            .DIN(N__11827),
            .DOUT(N__11826),
            .PACKAGEPIN(CLK28_IN));
    defparam CLK28_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK28_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK28_IN_ibuf_gb_io_preio (
            .PADOEN(N__11828),
            .PADOUT(N__11827),
            .PADIN(N__11826),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__11817),
            .DIN(N__11816),
            .DOUT(N__11815),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__11817),
            .PADOUT(N__11816),
            .PADIN(N__11815),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_0_iopad (
            .OE(N__11808),
            .DIN(N__11807),
            .DOUT(N__11806),
            .PACKAGEPIN(TT[0]));
    defparam TT_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_0_preio (
            .PADOEN(N__11808),
            .PADOUT(N__11807),
            .PADIN(N__11806),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ROM_DELAY_ibuf_1_iopad.PULLUP=1'b1;
    IO_PAD ROM_DELAY_ibuf_1_iopad (
            .OE(N__11799),
            .DIN(N__11798),
            .DOUT(N__11797),
            .PACKAGEPIN(ROM_DELAY[1]));
    defparam ROM_DELAY_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam ROM_DELAY_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ROM_DELAY_ibuf_1_preio (
            .PADOEN(N__11799),
            .PADOUT(N__11798),
            .PADIN(N__11797),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ROM_DELAY_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_7_iopad (
            .OE(N__11790),
            .DIN(N__11789),
            .DOUT(N__11788),
            .PACKAGEPIN(D[7]));
    defparam D_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_7_preio (
            .PADOEN(N__11790),
            .PADOUT(N__11789),
            .PADIN(N__11788),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4757),
            .DIN0(D_in_7),
            .DOUT0(N__6326),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__11781),
            .DIN(N__11780),
            .DOUT(N__11779),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__11781),
            .PADOUT(N__11780),
            .PADIN(N__11779),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CPUCONFn_ibuf_iopad (
            .OE(N__11772),
            .DIN(N__11771),
            .DOUT(N__11770),
            .PACKAGEPIN(CPUCONFn));
    defparam CPUCONFn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CPUCONFn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CPUCONFn_ibuf_preio (
            .PADOEN(N__11772),
            .PADOUT(N__11771),
            .PADIN(N__11770),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CPUCONFn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RTC_ENn_obuf_iopad (
            .OE(N__11763),
            .DIN(N__11762),
            .DOUT(N__11761),
            .PACKAGEPIN(RTC_ENn));
    defparam RTC_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RTC_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RTC_ENn_obuf_preio (
            .PADOEN(N__11763),
            .PADOUT(N__11762),
            .PADIN(N__11761),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4352),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_24_iopad (
            .OE(N__11754),
            .DIN(N__11753),
            .DOUT(N__11752),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__11754),
            .PADOUT(N__11753),
            .PADIN(N__11752),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SPIO_J_ibuf_iopad.PULLUP=1'b1;
    IO_PAD SPIO_J_ibuf_iopad (
            .OE(N__11745),
            .DIN(N__11744),
            .DOUT(N__11743),
            .PACKAGEPIN(SPIO_J));
    defparam SPIO_J_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam SPIO_J_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO SPIO_J_ibuf_preio (
            .PADOEN(N__11745),
            .PADOUT(N__11744),
            .PADIN(N__11743),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SPIO_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_4_iopad (
            .OE(N__11736),
            .DIN(N__11735),
            .DOUT(N__11734),
            .PACKAGEPIN(D[4]));
    defparam D_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_4_preio (
            .PADOEN(N__11736),
            .PADOUT(N__11735),
            .PADIN(N__11734),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4742),
            .DIN0(D_in_4),
            .DOUT0(N__7022),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PPIO_obuf_iopad (
            .OE(N__11727),
            .DIN(N__11726),
            .DOUT(N__11725),
            .PACKAGEPIN(PPIO));
    defparam PPIO_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PPIO_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PPIO_obuf_preio (
            .PADOEN(N__11727),
            .PADOUT(N__11726),
            .PADIN(N__11725),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4253),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__11718),
            .DIN(N__11717),
            .DOUT(N__11716),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__11718),
            .PADOUT(N__11717),
            .PADIN(N__11716),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_21_iopad (
            .OE(N__11709),
            .DIN(N__11708),
            .DOUT(N__11707),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__11709),
            .PADOUT(N__11708),
            .PADIN(N__11707),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam PPIO_J_ibuf_iopad.PULLUP=1'b1;
    IO_PAD PPIO_J_ibuf_iopad (
            .OE(N__11700),
            .DIN(N__11699),
            .DOUT(N__11698),
            .PACKAGEPIN(PPIO_J));
    defparam PPIO_J_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam PPIO_J_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO PPIO_J_ibuf_preio (
            .PADOEN(N__11700),
            .PADOUT(N__11699),
            .PADIN(N__11698),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(PPIO_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_obuf_iopad (
            .OE(N__11691),
            .DIN(N__11690),
            .DOUT(N__11689),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMSPACEn_obuf_preio (
            .PADOEN(N__11691),
            .PADOUT(N__11690),
            .PADIN(N__11689),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6068),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__11682),
            .DIN(N__11681),
            .DOUT(N__11680),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__11682),
            .PADOUT(N__11681),
            .PADIN(N__11680),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ROMENn_obuf_iopad (
            .OE(N__11673),
            .DIN(N__11672),
            .DOUT(N__11671),
            .PACKAGEPIN(ROMENn));
    defparam ROMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ROMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ROMENn_obuf_preio (
            .PADOEN(N__11673),
            .PADOUT(N__11672),
            .PADIN(N__11671),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9899),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_obuft_iopad (
            .OE(N__11664),
            .DIN(N__11663),
            .DOUT(N__11662),
            .PACKAGEPIN(TBIn));
    defparam TBIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TBIn_obuft_preio (
            .PADOEN(N__11664),
            .PADOUT(N__11663),
            .PADIN(N__11662),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9108),
            .DIN0(),
            .DOUT0(N__7615),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam AUTOBOOT_ibuf_iopad.PULLUP=1'b1;
    IO_PAD AUTOBOOT_ibuf_iopad (
            .OE(N__11655),
            .DIN(N__11654),
            .DOUT(N__11653),
            .PACKAGEPIN(AUTOBOOT));
    defparam AUTOBOOT_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AUTOBOOT_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AUTOBOOT_ibuf_preio (
            .PADOEN(N__11655),
            .PADOUT(N__11654),
            .PADIN(N__11653),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AUTOBOOT_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__11646),
            .DIN(N__11645),
            .DOUT(N__11644),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__11646),
            .PADOUT(N__11645),
            .PADIN(N__11644),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PORTSIZE_obuf_iopad (
            .OE(N__11637),
            .DIN(N__11636),
            .DOUT(N__11635),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PORTSIZE_obuf_preio (
            .PADOEN(N__11637),
            .PADOUT(N__11636),
            .PADIN(N__11635),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5255),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD F_ENn_obuf_iopad (
            .OE(N__11628),
            .DIN(N__11627),
            .DOUT(N__11626),
            .PACKAGEPIN(F_ENn));
    defparam F_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam F_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO F_ENn_obuf_preio (
            .PADOEN(N__11628),
            .PADOUT(N__11627),
            .PADIN(N__11626),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11176),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__11619),
            .DIN(N__11618),
            .DOUT(N__11617),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__11619),
            .PADOUT(N__11618),
            .PADIN(N__11617),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_22_iopad (
            .OE(N__11610),
            .DIN(N__11609),
            .DOUT(N__11608),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__11610),
            .PADOUT(N__11609),
            .PADIN(N__11608),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__11601),
            .DIN(N__11600),
            .DOUT(N__11599),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__11601),
            .PADOUT(N__11600),
            .PADIN(N__11599),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__11592),
            .DIN(N__11591),
            .DOUT(N__11590),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__11592),
            .PADOUT(N__11591),
            .PADIN(N__11590),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__11583),
            .DIN(N__11582),
            .DOUT(N__11581),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__11583),
            .PADOUT(N__11582),
            .PADIN(N__11581),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ROM_DELAY_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD ROM_DELAY_ibuf_0_iopad (
            .OE(N__11574),
            .DIN(N__11573),
            .DOUT(N__11572),
            .PACKAGEPIN(ROM_DELAY[0]));
    defparam ROM_DELAY_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam ROM_DELAY_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO ROM_DELAY_ibuf_0_preio (
            .PADOEN(N__11574),
            .PADOUT(N__11573),
            .PADIN(N__11572),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ROM_DELAY_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SCS1_obuf_iopad (
            .OE(N__11565),
            .DIN(N__11564),
            .DOUT(N__11563),
            .PACKAGEPIN(SCS1));
    defparam SCS1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam SCS1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO SCS1_obuf_preio (
            .PADOEN(N__11565),
            .PADOUT(N__11564),
            .PADIN(N__11563),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10703),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_CLK_obuf_iopad (
            .OE(N__11556),
            .DIN(N__11555),
            .DOUT(N__11554),
            .PACKAGEPIN(AGNUS_CLK));
    defparam AGNUS_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO AGNUS_CLK_obuf_preio (
            .PADOEN(N__11556),
            .PADOUT(N__11555),
            .PADIN(N__11554),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11102),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_25_iopad (
            .OE(N__11547),
            .DIN(N__11546),
            .DOUT(N__11545),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__11547),
            .PADOUT(N__11546),
            .PADIN(N__11545),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS0n_obuf_iopad (
            .OE(N__11538),
            .DIN(N__11537),
            .DOUT(N__11536),
            .PACKAGEPIN(CIACS0n));
    defparam CIACS0n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS0n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS0n_obuf_preio (
            .PADOEN(N__11538),
            .PADOUT(N__11537),
            .PADIN(N__11536),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8417),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK50_obuf_iopad (
            .OE(N__11529),
            .DIN(N__11528),
            .DOUT(N__11527),
            .PACKAGEPIN(TICK50));
    defparam TICK50_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK50_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK50_obuf_preio (
            .PADOEN(N__11529),
            .PADOUT(N__11528),
            .PADIN(N__11527),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9383),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__11520),
            .DIN(N__11519),
            .DOUT(N__11518),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__11520),
            .PADOUT(N__11519),
            .PADIN(N__11518),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_28_iopad (
            .OE(N__11511),
            .DIN(N__11510),
            .DOUT(N__11509),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__11511),
            .PADOUT(N__11510),
            .PADIN(N__11509),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_30_iopad (
            .OE(N__11502),
            .DIN(N__11501),
            .DOUT(N__11500),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__11502),
            .PADOUT(N__11501),
            .PADIN(N__11500),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD OVL_ibuf_iopad (
            .OE(N__11493),
            .DIN(N__11492),
            .DOUT(N__11491),
            .PACKAGEPIN(OVL));
    defparam OVL_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam OVL_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO OVL_ibuf_preio (
            .PADOEN(N__11493),
            .PADOUT(N__11492),
            .PADIN(N__11491),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(OVL_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_obuft_iopad (
            .OE(N__11484),
            .DIN(N__11483),
            .DOUT(N__11482),
            .PACKAGEPIN(TCIn));
    defparam TCIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TCIn_obuft_preio (
            .PADOEN(N__11484),
            .PADOUT(N__11483),
            .PADIN(N__11482),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9122),
            .DIN0(),
            .DOUT0(N__7544),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_5_iopad (
            .OE(N__11475),
            .DIN(N__11474),
            .DOUT(N__11473),
            .PACKAGEPIN(D[5]));
    defparam D_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_5_preio (
            .PADOEN(N__11475),
            .PADOUT(N__11474),
            .PADIN(N__11473),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4752),
            .DIN0(D_in_5),
            .DOUT0(N__6359),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD XCLK_ENn_ibuf_iopad (
            .OE(N__11466),
            .DIN(N__11465),
            .DOUT(N__11464),
            .PACKAGEPIN(XCLK_ENn));
    defparam XCLK_ENn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam XCLK_ENn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO XCLK_ENn_ibuf_preio (
            .PADOEN(N__11466),
            .PADOUT(N__11465),
            .PADIN(N__11464),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(XCLK_ENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__11457),
            .DIN(N__11456),
            .DOUT(N__11455),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__11457),
            .PADOUT(N__11456),
            .PADIN(N__11455),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__11448),
            .DIN(N__11447),
            .DOUT(N__11446),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__11448),
            .PADOUT(N__11447),
            .PADIN(N__11446),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__11439),
            .DIN(N__11438),
            .DOUT(N__11437),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__11439),
            .PADOUT(N__11438),
            .PADIN(N__11437),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CONFIGENn_obuf_iopad (
            .OE(N__11430),
            .DIN(N__11429),
            .DOUT(N__11428),
            .PACKAGEPIN(CONFIGENn));
    defparam CONFIGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CONFIGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CONFIGENn_obuf_preio (
            .PADOEN(N__11430),
            .PADOUT(N__11429),
            .PADIN(N__11428),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6299),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SPIO_obuf_iopad (
            .OE(N__11421),
            .DIN(N__11420),
            .DOUT(N__11419),
            .PACKAGEPIN(SPIO));
    defparam SPIO_obuf_preio.NEG_TRIGGER=1'b0;
    defparam SPIO_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO SPIO_obuf_preio (
            .PADOEN(N__11421),
            .PADOUT(N__11420),
            .PADIN(N__11419),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4316),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK60_obuf_iopad (
            .OE(N__11412),
            .DIN(N__11411),
            .DOUT(N__11410),
            .PACKAGEPIN(TICK60));
    defparam TICK60_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK60_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK60_obuf_preio (
            .PADOEN(N__11412),
            .PADOUT(N__11411),
            .PADIN(N__11410),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9413),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_26_iopad (
            .OE(N__11403),
            .DIN(N__11402),
            .DOUT(N__11401),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__11403),
            .PADOUT(N__11402),
            .PADIN(N__11401),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_23_iopad (
            .OE(N__11394),
            .DIN(N__11393),
            .DOUT(N__11392),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__11394),
            .PADOUT(N__11393),
            .PADIN(N__11392),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__11385),
            .DIN(N__11384),
            .DOUT(N__11383),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__11385),
            .PADOUT(N__11384),
            .PADIN(N__11383),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ATA_ENn_obuf_iopad (
            .OE(N__11376),
            .DIN(N__11375),
            .DOUT(N__11374),
            .PACKAGEPIN(ATA_ENn));
    defparam ATA_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ATA_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ATA_ENn_obuf_preio (
            .PADOEN(N__11376),
            .PADOUT(N__11375),
            .PADIN(N__11374),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5213),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_31_iopad (
            .OE(N__11367),
            .DIN(N__11366),
            .DOUT(N__11365),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__11367),
            .PADOUT(N__11366),
            .PADIN(N__11365),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS1n_obuf_iopad (
            .OE(N__11358),
            .DIN(N__11357),
            .DOUT(N__11356),
            .PACKAGEPIN(CIACS1n));
    defparam CIACS1n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS1n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS1n_obuf_preio (
            .PADOEN(N__11358),
            .PADOUT(N__11357),
            .PADIN(N__11356),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8342),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_obuf_iopad (
            .OE(N__11349),
            .DIN(N__11348),
            .DOUT(N__11347),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGSPACEn_obuf_preio (
            .PADOEN(N__11349),
            .PADOUT(N__11348),
            .PADIN(N__11347),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4571),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PCS0_obuf_iopad (
            .OE(N__11340),
            .DIN(N__11339),
            .DOUT(N__11338),
            .PACKAGEPIN(PCS0));
    defparam PCS0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PCS0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PCS0_obuf_preio (
            .PADOEN(N__11340),
            .PADOUT(N__11339),
            .PADIN(N__11338),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10787),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__11331),
            .DIN(N__11330),
            .DOUT(N__11329),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__11331),
            .PADOUT(N__11330),
            .PADIN(N__11329),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_CIA_obuf_iopad (
            .OE(N__11322),
            .DIN(N__11321),
            .DOUT(N__11320),
            .PACKAGEPIN(CLK_CIA));
    defparam CLK_CIA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_CIA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_CIA_obuf_preio (
            .PADOEN(N__11322),
            .PADOUT(N__11321),
            .PADIN(N__11320),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9641),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__11313),
            .DIN(N__11312),
            .DOUT(N__11311),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__11313),
            .PADOUT(N__11312),
            .PADIN(N__11311),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PCS1_obuf_iopad (
            .OE(N__11304),
            .DIN(N__11303),
            .DOUT(N__11302),
            .PACKAGEPIN(PCS1));
    defparam PCS1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PCS1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PCS1_obuf_preio (
            .PADOEN(N__11304),
            .PADOUT(N__11303),
            .PADIN(N__11302),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10841),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__11295),
            .DIN(N__11294),
            .DOUT(N__11293),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__11295),
            .PADOUT(N__11294),
            .PADIN(N__11293),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9121),
            .DIN0(TACKn_in),
            .DOUT0(N__7622),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_1_iopad (
            .OE(N__11286),
            .DIN(N__11285),
            .DOUT(N__11284),
            .PACKAGEPIN(TT[1]));
    defparam TT_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_1_preio (
            .PADOEN(N__11286),
            .PADOUT(N__11285),
            .PADIN(N__11284),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__11277),
            .DIN(N__11276),
            .DOUT(N__11275),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__11277),
            .PADOUT(N__11276),
            .PADIN(N__11275),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5234),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_29_iopad (
            .OE(N__11268),
            .DIN(N__11267),
            .DOUT(N__11266),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__11268),
            .PADOUT(N__11267),
            .PADIN(N__11266),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_6_iopad (
            .OE(N__11259),
            .DIN(N__11258),
            .DOUT(N__11257),
            .PACKAGEPIN(D[6]));
    defparam D_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_6_preio (
            .PADOEN(N__11259),
            .PADOUT(N__11258),
            .PADIN(N__11257),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4753),
            .DIN0(D_in_6),
            .DOUT0(N__5462),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__11250),
            .DIN(N__11249),
            .DOUT(N__11248),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__11250),
            .PADOUT(N__11249),
            .PADIN(N__11248),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_27_iopad (
            .OE(N__11241),
            .DIN(N__11240),
            .DOUT(N__11239),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__11241),
            .PADOUT(N__11240),
            .PADIN(N__11239),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SCS0_obuf_iopad (
            .OE(N__11232),
            .DIN(N__11231),
            .DOUT(N__11230),
            .PACKAGEPIN(SCS0));
    defparam SCS0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam SCS0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO SCS0_obuf_preio (
            .PADOEN(N__11232),
            .PADOUT(N__11231),
            .PADIN(N__11230),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10823),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD XCLK_ibuf_iopad (
            .OE(N__11223),
            .DIN(N__11222),
            .DOUT(N__11221),
            .PACKAGEPIN(XCLK));
    defparam XCLK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam XCLK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO XCLK_ibuf_preio (
            .PADOEN(N__11223),
            .PADOUT(N__11222),
            .PADIN(N__11221),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(XCLK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__11214),
            .DIN(N__11213),
            .DOUT(N__11212),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__11214),
            .PADOUT(N__11213),
            .PADIN(N__11212),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__11205),
            .DIN(N__11204),
            .DOUT(N__11203),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__11205),
            .PADOUT(N__11204),
            .PADIN(N__11203),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IoInMux I__2688 (
            .O(N__11186),
            .I(N__11183));
    LocalMux I__2687 (
            .O(N__11183),
            .I(N__11180));
    Span4Mux_s2_v I__2686 (
            .O(N__11180),
            .I(N__11177));
    Sp12to4 I__2685 (
            .O(N__11177),
            .I(N__11173));
    IoInMux I__2684 (
            .O(N__11176),
            .I(N__11170));
    Span12Mux_h I__2683 (
            .O(N__11173),
            .I(N__11167));
    LocalMux I__2682 (
            .O(N__11170),
            .I(N__11164));
    Span12Mux_v I__2681 (
            .O(N__11167),
            .I(N__11161));
    Span12Mux_s6_h I__2680 (
            .O(N__11164),
            .I(N__11158));
    Odrv12 I__2679 (
            .O(N__11161),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__2678 (
            .O(N__11158),
            .I(CONSTANT_ONE_NET));
    InMux I__2677 (
            .O(N__11153),
            .I(N__11150));
    LocalMux I__2676 (
            .O(N__11150),
            .I(N__11143));
    ClkMux I__2675 (
            .O(N__11149),
            .I(N__11132));
    ClkMux I__2674 (
            .O(N__11148),
            .I(N__11132));
    ClkMux I__2673 (
            .O(N__11147),
            .I(N__11132));
    ClkMux I__2672 (
            .O(N__11146),
            .I(N__11132));
    Glb2LocalMux I__2671 (
            .O(N__11143),
            .I(N__11132));
    GlobalMux I__2670 (
            .O(N__11132),
            .I(N__11129));
    gio2CtrlBuf I__2669 (
            .O(N__11129),
            .I(CLK28_IN_c_g));
    InMux I__2668 (
            .O(N__11126),
            .I(N__11123));
    LocalMux I__2667 (
            .O(N__11123),
            .I(N__11120));
    Span4Mux_v I__2666 (
            .O(N__11120),
            .I(N__11117));
    Odrv4 I__2665 (
            .O(N__11117),
            .I(XCLK_c));
    InMux I__2664 (
            .O(N__11114),
            .I(N__11111));
    LocalMux I__2663 (
            .O(N__11111),
            .I(N__11108));
    Span12Mux_v I__2662 (
            .O(N__11108),
            .I(N__11105));
    Odrv12 I__2661 (
            .O(N__11105),
            .I(XCLK_ENn_c));
    IoInMux I__2660 (
            .O(N__11102),
            .I(N__11099));
    LocalMux I__2659 (
            .O(N__11099),
            .I(N__11096));
    Span4Mux_s3_h I__2658 (
            .O(N__11096),
            .I(N__11093));
    Odrv4 I__2657 (
            .O(N__11093),
            .I(AGNUS_CLK_c));
    InMux I__2656 (
            .O(N__11090),
            .I(N__11086));
    InMux I__2655 (
            .O(N__11089),
            .I(N__11083));
    LocalMux I__2654 (
            .O(N__11086),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    LocalMux I__2653 (
            .O(N__11083),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    InMux I__2652 (
            .O(N__11078),
            .I(N__11075));
    LocalMux I__2651 (
            .O(N__11075),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ));
    InMux I__2650 (
            .O(N__11072),
            .I(\U409_TICK.un3_COUNTER60_1_cry_13 ));
    InMux I__2649 (
            .O(N__11069),
            .I(N__11065));
    InMux I__2648 (
            .O(N__11068),
            .I(N__11062));
    LocalMux I__2647 (
            .O(N__11065),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    LocalMux I__2646 (
            .O(N__11062),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    InMux I__2645 (
            .O(N__11057),
            .I(N__11054));
    LocalMux I__2644 (
            .O(N__11054),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ));
    InMux I__2643 (
            .O(N__11051),
            .I(\U409_TICK.un3_COUNTER60_1_cry_14 ));
    InMux I__2642 (
            .O(N__11048),
            .I(\U409_TICK.un3_COUNTER60_1_cry_15 ));
    InMux I__2641 (
            .O(N__11045),
            .I(N__11041));
    InMux I__2640 (
            .O(N__11044),
            .I(N__11038));
    LocalMux I__2639 (
            .O(N__11041),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    LocalMux I__2638 (
            .O(N__11038),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    CascadeMux I__2637 (
            .O(N__11033),
            .I(N__11025));
    InMux I__2636 (
            .O(N__11032),
            .I(N__11018));
    InMux I__2635 (
            .O(N__11031),
            .I(N__11018));
    InMux I__2634 (
            .O(N__11030),
            .I(N__11015));
    InMux I__2633 (
            .O(N__11029),
            .I(N__11012));
    InMux I__2632 (
            .O(N__11028),
            .I(N__11003));
    InMux I__2631 (
            .O(N__11025),
            .I(N__11003));
    InMux I__2630 (
            .O(N__11024),
            .I(N__11003));
    InMux I__2629 (
            .O(N__11023),
            .I(N__11003));
    LocalMux I__2628 (
            .O(N__11018),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__2627 (
            .O(N__11015),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__2626 (
            .O(N__11012),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__2625 (
            .O(N__11003),
            .I(\U409_TICK.TICK503_9 ));
    CascadeMux I__2624 (
            .O(N__10994),
            .I(N__10990));
    InMux I__2623 (
            .O(N__10993),
            .I(N__10984));
    InMux I__2622 (
            .O(N__10990),
            .I(N__10978));
    InMux I__2621 (
            .O(N__10989),
            .I(N__10975));
    InMux I__2620 (
            .O(N__10988),
            .I(N__10972));
    InMux I__2619 (
            .O(N__10987),
            .I(N__10969));
    LocalMux I__2618 (
            .O(N__10984),
            .I(N__10966));
    InMux I__2617 (
            .O(N__10983),
            .I(N__10959));
    InMux I__2616 (
            .O(N__10982),
            .I(N__10959));
    InMux I__2615 (
            .O(N__10981),
            .I(N__10959));
    LocalMux I__2614 (
            .O(N__10978),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__2613 (
            .O(N__10975),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__2612 (
            .O(N__10972),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__2611 (
            .O(N__10969),
            .I(\U409_TICK.TICK503_14 ));
    Odrv4 I__2610 (
            .O(N__10966),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__2609 (
            .O(N__10959),
            .I(\U409_TICK.TICK503_14 ));
    CascadeMux I__2608 (
            .O(N__10946),
            .I(N__10942));
    InMux I__2607 (
            .O(N__10945),
            .I(N__10936));
    InMux I__2606 (
            .O(N__10942),
            .I(N__10936));
    CascadeMux I__2605 (
            .O(N__10941),
            .I(N__10933));
    LocalMux I__2604 (
            .O(N__10936),
            .I(N__10925));
    InMux I__2603 (
            .O(N__10933),
            .I(N__10922));
    InMux I__2602 (
            .O(N__10932),
            .I(N__10911));
    InMux I__2601 (
            .O(N__10931),
            .I(N__10911));
    InMux I__2600 (
            .O(N__10930),
            .I(N__10911));
    InMux I__2599 (
            .O(N__10929),
            .I(N__10911));
    InMux I__2598 (
            .O(N__10928),
            .I(N__10911));
    Span4Mux_h I__2597 (
            .O(N__10925),
            .I(N__10908));
    LocalMux I__2596 (
            .O(N__10922),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__2595 (
            .O(N__10911),
            .I(\U409_TICK.TICK503_10 ));
    Odrv4 I__2594 (
            .O(N__10908),
            .I(\U409_TICK.TICK503_10 ));
    InMux I__2593 (
            .O(N__10901),
            .I(N__10898));
    LocalMux I__2592 (
            .O(N__10898),
            .I(N__10895));
    Odrv4 I__2591 (
            .O(N__10895),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ));
    InMux I__2590 (
            .O(N__10892),
            .I(N__10888));
    InMux I__2589 (
            .O(N__10891),
            .I(N__10885));
    LocalMux I__2588 (
            .O(N__10888),
            .I(N__10882));
    LocalMux I__2587 (
            .O(N__10885),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    Odrv12 I__2586 (
            .O(N__10882),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    ClkMux I__2585 (
            .O(N__10877),
            .I(N__10847));
    ClkMux I__2584 (
            .O(N__10876),
            .I(N__10847));
    ClkMux I__2583 (
            .O(N__10875),
            .I(N__10847));
    ClkMux I__2582 (
            .O(N__10874),
            .I(N__10847));
    ClkMux I__2581 (
            .O(N__10873),
            .I(N__10847));
    ClkMux I__2580 (
            .O(N__10872),
            .I(N__10847));
    ClkMux I__2579 (
            .O(N__10871),
            .I(N__10847));
    ClkMux I__2578 (
            .O(N__10870),
            .I(N__10847));
    ClkMux I__2577 (
            .O(N__10869),
            .I(N__10847));
    ClkMux I__2576 (
            .O(N__10868),
            .I(N__10847));
    GlobalMux I__2575 (
            .O(N__10847),
            .I(N__10844));
    gio2CtrlBuf I__2574 (
            .O(N__10844),
            .I(CLK6_c_g));
    IoInMux I__2573 (
            .O(N__10841),
            .I(N__10838));
    LocalMux I__2572 (
            .O(N__10838),
            .I(N__10835));
    Span4Mux_s3_h I__2571 (
            .O(N__10835),
            .I(N__10832));
    Span4Mux_v I__2570 (
            .O(N__10832),
            .I(N__10829));
    Span4Mux_h I__2569 (
            .O(N__10829),
            .I(N__10826));
    Odrv4 I__2568 (
            .O(N__10826),
            .I(PCS1_c));
    IoInMux I__2567 (
            .O(N__10823),
            .I(N__10820));
    LocalMux I__2566 (
            .O(N__10820),
            .I(N__10817));
    IoSpan4Mux I__2565 (
            .O(N__10817),
            .I(N__10814));
    Span4Mux_s3_h I__2564 (
            .O(N__10814),
            .I(N__10811));
    Span4Mux_h I__2563 (
            .O(N__10811),
            .I(N__10808));
    Odrv4 I__2562 (
            .O(N__10808),
            .I(SCS0_c));
    InMux I__2561 (
            .O(N__10805),
            .I(N__10801));
    InMux I__2560 (
            .O(N__10804),
            .I(N__10798));
    LocalMux I__2559 (
            .O(N__10801),
            .I(N__10793));
    LocalMux I__2558 (
            .O(N__10798),
            .I(N__10793));
    Span12Mux_s10_h I__2557 (
            .O(N__10793),
            .I(N__10790));
    Odrv12 I__2556 (
            .O(N__10790),
            .I(\U409_ADDRESS_DECODE.CSZ0Z0 ));
    IoInMux I__2555 (
            .O(N__10787),
            .I(N__10784));
    LocalMux I__2554 (
            .O(N__10784),
            .I(N__10781));
    IoSpan4Mux I__2553 (
            .O(N__10781),
            .I(N__10778));
    Span4Mux_s3_v I__2552 (
            .O(N__10778),
            .I(N__10775));
    Span4Mux_v I__2551 (
            .O(N__10775),
            .I(N__10772));
    Odrv4 I__2550 (
            .O(N__10772),
            .I(PCS0_c));
    InMux I__2549 (
            .O(N__10769),
            .I(N__10763));
    InMux I__2548 (
            .O(N__10768),
            .I(N__10760));
    InMux I__2547 (
            .O(N__10767),
            .I(N__10757));
    InMux I__2546 (
            .O(N__10766),
            .I(N__10754));
    LocalMux I__2545 (
            .O(N__10763),
            .I(N__10749));
    LocalMux I__2544 (
            .O(N__10760),
            .I(N__10749));
    LocalMux I__2543 (
            .O(N__10757),
            .I(N__10744));
    LocalMux I__2542 (
            .O(N__10754),
            .I(N__10744));
    Span4Mux_v I__2541 (
            .O(N__10749),
            .I(N__10741));
    Span4Mux_v I__2540 (
            .O(N__10744),
            .I(N__10738));
    Sp12to4 I__2539 (
            .O(N__10741),
            .I(N__10735));
    Span4Mux_h I__2538 (
            .O(N__10738),
            .I(N__10732));
    Span12Mux_h I__2537 (
            .O(N__10735),
            .I(N__10727));
    Sp12to4 I__2536 (
            .O(N__10732),
            .I(N__10727));
    Span12Mux_h I__2535 (
            .O(N__10727),
            .I(N__10724));
    Odrv12 I__2534 (
            .O(N__10724),
            .I(A_c_14));
    InMux I__2533 (
            .O(N__10721),
            .I(N__10717));
    InMux I__2532 (
            .O(N__10720),
            .I(N__10714));
    LocalMux I__2531 (
            .O(N__10717),
            .I(N__10709));
    LocalMux I__2530 (
            .O(N__10714),
            .I(N__10709));
    Span12Mux_h I__2529 (
            .O(N__10709),
            .I(N__10706));
    Odrv12 I__2528 (
            .O(N__10706),
            .I(\U409_ADDRESS_DECODE.CSZ0Z1 ));
    IoInMux I__2527 (
            .O(N__10703),
            .I(N__10700));
    LocalMux I__2526 (
            .O(N__10700),
            .I(N__10697));
    IoSpan4Mux I__2525 (
            .O(N__10697),
            .I(N__10694));
    IoSpan4Mux I__2524 (
            .O(N__10694),
            .I(N__10691));
    Span4Mux_s3_h I__2523 (
            .O(N__10691),
            .I(N__10688));
    Odrv4 I__2522 (
            .O(N__10688),
            .I(SCS1_c));
    CascadeMux I__2521 (
            .O(N__10685),
            .I(N__10682));
    InMux I__2520 (
            .O(N__10682),
            .I(N__10678));
    InMux I__2519 (
            .O(N__10681),
            .I(N__10675));
    LocalMux I__2518 (
            .O(N__10678),
            .I(N__10670));
    LocalMux I__2517 (
            .O(N__10675),
            .I(N__10670));
    Odrv4 I__2516 (
            .O(N__10670),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    InMux I__2515 (
            .O(N__10667),
            .I(N__10664));
    LocalMux I__2514 (
            .O(N__10664),
            .I(N__10661));
    Odrv4 I__2513 (
            .O(N__10661),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ));
    InMux I__2512 (
            .O(N__10658),
            .I(\U409_TICK.un3_COUNTER60_1_cry_5 ));
    InMux I__2511 (
            .O(N__10655),
            .I(N__10651));
    InMux I__2510 (
            .O(N__10654),
            .I(N__10648));
    LocalMux I__2509 (
            .O(N__10651),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    LocalMux I__2508 (
            .O(N__10648),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    InMux I__2507 (
            .O(N__10643),
            .I(\U409_TICK.un3_COUNTER60_1_cry_6 ));
    InMux I__2506 (
            .O(N__10640),
            .I(N__10636));
    InMux I__2505 (
            .O(N__10639),
            .I(N__10633));
    LocalMux I__2504 (
            .O(N__10636),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    LocalMux I__2503 (
            .O(N__10633),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    InMux I__2502 (
            .O(N__10628),
            .I(N__10625));
    LocalMux I__2501 (
            .O(N__10625),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ));
    InMux I__2500 (
            .O(N__10622),
            .I(\U409_TICK.un3_COUNTER60_1_cry_7 ));
    InMux I__2499 (
            .O(N__10619),
            .I(N__10615));
    InMux I__2498 (
            .O(N__10618),
            .I(N__10612));
    LocalMux I__2497 (
            .O(N__10615),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    LocalMux I__2496 (
            .O(N__10612),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    CascadeMux I__2495 (
            .O(N__10607),
            .I(N__10604));
    InMux I__2494 (
            .O(N__10604),
            .I(N__10601));
    LocalMux I__2493 (
            .O(N__10601),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ));
    InMux I__2492 (
            .O(N__10598),
            .I(bfn_17_6_0_));
    InMux I__2491 (
            .O(N__10595),
            .I(N__10591));
    InMux I__2490 (
            .O(N__10594),
            .I(N__10588));
    LocalMux I__2489 (
            .O(N__10591),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    LocalMux I__2488 (
            .O(N__10588),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    InMux I__2487 (
            .O(N__10583),
            .I(\U409_TICK.un3_COUNTER60_1_cry_9 ));
    InMux I__2486 (
            .O(N__10580),
            .I(N__10577));
    LocalMux I__2485 (
            .O(N__10577),
            .I(N__10574));
    Span4Mux_h I__2484 (
            .O(N__10574),
            .I(N__10570));
    InMux I__2483 (
            .O(N__10573),
            .I(N__10567));
    Odrv4 I__2482 (
            .O(N__10570),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    LocalMux I__2481 (
            .O(N__10567),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    InMux I__2480 (
            .O(N__10562),
            .I(\U409_TICK.un3_COUNTER60_1_cry_10 ));
    InMux I__2479 (
            .O(N__10559),
            .I(N__10555));
    InMux I__2478 (
            .O(N__10558),
            .I(N__10552));
    LocalMux I__2477 (
            .O(N__10555),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    LocalMux I__2476 (
            .O(N__10552),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    InMux I__2475 (
            .O(N__10547),
            .I(\U409_TICK.un3_COUNTER60_1_cry_11 ));
    CascadeMux I__2474 (
            .O(N__10544),
            .I(N__10541));
    InMux I__2473 (
            .O(N__10541),
            .I(N__10537));
    InMux I__2472 (
            .O(N__10540),
            .I(N__10534));
    LocalMux I__2471 (
            .O(N__10537),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    LocalMux I__2470 (
            .O(N__10534),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    InMux I__2469 (
            .O(N__10529),
            .I(\U409_TICK.un3_COUNTER60_1_cry_12 ));
    InMux I__2468 (
            .O(N__10526),
            .I(N__10523));
    LocalMux I__2467 (
            .O(N__10523),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ));
    InMux I__2466 (
            .O(N__10520),
            .I(N__10516));
    InMux I__2465 (
            .O(N__10519),
            .I(N__10513));
    LocalMux I__2464 (
            .O(N__10516),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    LocalMux I__2463 (
            .O(N__10513),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    InMux I__2462 (
            .O(N__10508),
            .I(N__10504));
    InMux I__2461 (
            .O(N__10507),
            .I(N__10501));
    LocalMux I__2460 (
            .O(N__10504),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    LocalMux I__2459 (
            .O(N__10501),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    CascadeMux I__2458 (
            .O(N__10496),
            .I(N__10493));
    InMux I__2457 (
            .O(N__10493),
            .I(N__10489));
    InMux I__2456 (
            .O(N__10492),
            .I(N__10486));
    LocalMux I__2455 (
            .O(N__10489),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    LocalMux I__2454 (
            .O(N__10486),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    InMux I__2453 (
            .O(N__10481),
            .I(N__10477));
    InMux I__2452 (
            .O(N__10480),
            .I(N__10474));
    LocalMux I__2451 (
            .O(N__10477),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    LocalMux I__2450 (
            .O(N__10474),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    CascadeMux I__2449 (
            .O(N__10469),
            .I(\U409_TICK.TICK503_10_cascade_ ));
    InMux I__2448 (
            .O(N__10466),
            .I(N__10463));
    LocalMux I__2447 (
            .O(N__10463),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ));
    InMux I__2446 (
            .O(N__10460),
            .I(N__10456));
    InMux I__2445 (
            .O(N__10459),
            .I(N__10453));
    LocalMux I__2444 (
            .O(N__10456),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    LocalMux I__2443 (
            .O(N__10453),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    CascadeMux I__2442 (
            .O(N__10448),
            .I(N__10444));
    InMux I__2441 (
            .O(N__10447),
            .I(N__10438));
    InMux I__2440 (
            .O(N__10444),
            .I(N__10438));
    InMux I__2439 (
            .O(N__10443),
            .I(N__10435));
    LocalMux I__2438 (
            .O(N__10438),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__2437 (
            .O(N__10435),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    CascadeMux I__2436 (
            .O(N__10430),
            .I(N__10426));
    CascadeMux I__2435 (
            .O(N__10429),
            .I(N__10421));
    InMux I__2434 (
            .O(N__10426),
            .I(N__10416));
    InMux I__2433 (
            .O(N__10425),
            .I(N__10416));
    InMux I__2432 (
            .O(N__10424),
            .I(N__10413));
    InMux I__2431 (
            .O(N__10421),
            .I(N__10410));
    LocalMux I__2430 (
            .O(N__10416),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__2429 (
            .O(N__10413),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__2428 (
            .O(N__10410),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    InMux I__2427 (
            .O(N__10403),
            .I(N__10399));
    InMux I__2426 (
            .O(N__10402),
            .I(N__10396));
    LocalMux I__2425 (
            .O(N__10399),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    LocalMux I__2424 (
            .O(N__10396),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    InMux I__2423 (
            .O(N__10391),
            .I(\U409_TICK.un3_COUNTER60_1_cry_1 ));
    InMux I__2422 (
            .O(N__10388),
            .I(N__10385));
    LocalMux I__2421 (
            .O(N__10385),
            .I(N__10381));
    InMux I__2420 (
            .O(N__10384),
            .I(N__10378));
    Odrv4 I__2419 (
            .O(N__10381),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    LocalMux I__2418 (
            .O(N__10378),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    InMux I__2417 (
            .O(N__10373),
            .I(\U409_TICK.un3_COUNTER60_1_cry_2 ));
    CascadeMux I__2416 (
            .O(N__10370),
            .I(N__10367));
    InMux I__2415 (
            .O(N__10367),
            .I(N__10363));
    InMux I__2414 (
            .O(N__10366),
            .I(N__10360));
    LocalMux I__2413 (
            .O(N__10363),
            .I(N__10357));
    LocalMux I__2412 (
            .O(N__10360),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    Odrv12 I__2411 (
            .O(N__10357),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    InMux I__2410 (
            .O(N__10352),
            .I(N__10349));
    LocalMux I__2409 (
            .O(N__10349),
            .I(N__10346));
    Odrv4 I__2408 (
            .O(N__10346),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ));
    InMux I__2407 (
            .O(N__10343),
            .I(\U409_TICK.un3_COUNTER60_1_cry_3 ));
    InMux I__2406 (
            .O(N__10340),
            .I(N__10337));
    LocalMux I__2405 (
            .O(N__10337),
            .I(N__10333));
    InMux I__2404 (
            .O(N__10336),
            .I(N__10330));
    Odrv4 I__2403 (
            .O(N__10333),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    LocalMux I__2402 (
            .O(N__10330),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    InMux I__2401 (
            .O(N__10325),
            .I(\U409_TICK.un3_COUNTER60_1_cry_4 ));
    CascadeMux I__2400 (
            .O(N__10322),
            .I(N__10314));
    CascadeMux I__2399 (
            .O(N__10321),
            .I(N__10311));
    InMux I__2398 (
            .O(N__10320),
            .I(N__10303));
    InMux I__2397 (
            .O(N__10319),
            .I(N__10303));
    InMux I__2396 (
            .O(N__10318),
            .I(N__10303));
    InMux I__2395 (
            .O(N__10317),
            .I(N__10294));
    InMux I__2394 (
            .O(N__10314),
            .I(N__10294));
    InMux I__2393 (
            .O(N__10311),
            .I(N__10294));
    InMux I__2392 (
            .O(N__10310),
            .I(N__10294));
    LocalMux I__2391 (
            .O(N__10303),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__2390 (
            .O(N__10294),
            .I(\U409_TICK.TICK603_10 ));
    InMux I__2389 (
            .O(N__10289),
            .I(N__10272));
    InMux I__2388 (
            .O(N__10288),
            .I(N__10272));
    InMux I__2387 (
            .O(N__10287),
            .I(N__10272));
    InMux I__2386 (
            .O(N__10286),
            .I(N__10272));
    InMux I__2385 (
            .O(N__10285),
            .I(N__10272));
    InMux I__2384 (
            .O(N__10284),
            .I(N__10267));
    InMux I__2383 (
            .O(N__10283),
            .I(N__10267));
    LocalMux I__2382 (
            .O(N__10272),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__2381 (
            .O(N__10267),
            .I(\U409_TICK.TICK603_14 ));
    CascadeMux I__2380 (
            .O(N__10262),
            .I(N__10259));
    InMux I__2379 (
            .O(N__10259),
            .I(N__10250));
    InMux I__2378 (
            .O(N__10258),
            .I(N__10247));
    InMux I__2377 (
            .O(N__10257),
            .I(N__10236));
    InMux I__2376 (
            .O(N__10256),
            .I(N__10236));
    InMux I__2375 (
            .O(N__10255),
            .I(N__10236));
    InMux I__2374 (
            .O(N__10254),
            .I(N__10236));
    InMux I__2373 (
            .O(N__10253),
            .I(N__10236));
    LocalMux I__2372 (
            .O(N__10250),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__2371 (
            .O(N__10247),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__2370 (
            .O(N__10236),
            .I(\U409_TICK.TICK603_9 ));
    CascadeMux I__2369 (
            .O(N__10229),
            .I(\U409_TICK.TICK603_10_cascade_ ));
    InMux I__2368 (
            .O(N__10226),
            .I(N__10222));
    InMux I__2367 (
            .O(N__10225),
            .I(N__10219));
    LocalMux I__2366 (
            .O(N__10222),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    LocalMux I__2365 (
            .O(N__10219),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    InMux I__2364 (
            .O(N__10214),
            .I(N__10211));
    LocalMux I__2363 (
            .O(N__10211),
            .I(N__10208));
    Odrv12 I__2362 (
            .O(N__10208),
            .I(\U409_TICK.TICK503_11 ));
    InMux I__2361 (
            .O(N__10205),
            .I(N__10201));
    InMux I__2360 (
            .O(N__10204),
            .I(N__10198));
    LocalMux I__2359 (
            .O(N__10201),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    LocalMux I__2358 (
            .O(N__10198),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    CascadeMux I__2357 (
            .O(N__10193),
            .I(\U409_TICK.TICK503_8_cascade_ ));
    InMux I__2356 (
            .O(N__10190),
            .I(N__10186));
    InMux I__2355 (
            .O(N__10189),
            .I(N__10183));
    LocalMux I__2354 (
            .O(N__10186),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    LocalMux I__2353 (
            .O(N__10183),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    CascadeMux I__2352 (
            .O(N__10178),
            .I(\U409_TICK.TICK503_14_cascade_ ));
    InMux I__2351 (
            .O(N__10175),
            .I(N__10172));
    LocalMux I__2350 (
            .O(N__10172),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ));
    InMux I__2349 (
            .O(N__10169),
            .I(N__10166));
    LocalMux I__2348 (
            .O(N__10166),
            .I(N__10161));
    CascadeMux I__2347 (
            .O(N__10165),
            .I(N__10158));
    CascadeMux I__2346 (
            .O(N__10164),
            .I(N__10154));
    Span4Mux_h I__2345 (
            .O(N__10161),
            .I(N__10151));
    InMux I__2344 (
            .O(N__10158),
            .I(N__10146));
    InMux I__2343 (
            .O(N__10157),
            .I(N__10146));
    InMux I__2342 (
            .O(N__10154),
            .I(N__10143));
    Odrv4 I__2341 (
            .O(N__10151),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__2340 (
            .O(N__10146),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__2339 (
            .O(N__10143),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    InMux I__2338 (
            .O(N__10136),
            .I(N__10133));
    LocalMux I__2337 (
            .O(N__10133),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ));
    InMux I__2336 (
            .O(N__10130),
            .I(N__10126));
    InMux I__2335 (
            .O(N__10129),
            .I(N__10123));
    LocalMux I__2334 (
            .O(N__10126),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    LocalMux I__2333 (
            .O(N__10123),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    InMux I__2332 (
            .O(N__10118),
            .I(N__10114));
    InMux I__2331 (
            .O(N__10117),
            .I(N__10111));
    LocalMux I__2330 (
            .O(N__10114),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    LocalMux I__2329 (
            .O(N__10111),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    CascadeMux I__2328 (
            .O(N__10106),
            .I(N__10103));
    InMux I__2327 (
            .O(N__10103),
            .I(N__10099));
    InMux I__2326 (
            .O(N__10102),
            .I(N__10096));
    LocalMux I__2325 (
            .O(N__10099),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    LocalMux I__2324 (
            .O(N__10096),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    CascadeMux I__2323 (
            .O(N__10091),
            .I(\U409_TICK.TICK503_9_cascade_ ));
    InMux I__2322 (
            .O(N__10088),
            .I(N__10085));
    LocalMux I__2321 (
            .O(N__10085),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ));
    InMux I__2320 (
            .O(N__10082),
            .I(N__10077));
    InMux I__2319 (
            .O(N__10081),
            .I(N__10072));
    InMux I__2318 (
            .O(N__10080),
            .I(N__10072));
    LocalMux I__2317 (
            .O(N__10077),
            .I(\U409_TRANSFER_ACK.N_11 ));
    LocalMux I__2316 (
            .O(N__10072),
            .I(\U409_TRANSFER_ACK.N_11 ));
    InMux I__2315 (
            .O(N__10067),
            .I(N__10064));
    LocalMux I__2314 (
            .O(N__10064),
            .I(N__10059));
    InMux I__2313 (
            .O(N__10063),
            .I(N__10053));
    InMux I__2312 (
            .O(N__10062),
            .I(N__10053));
    Span4Mux_h I__2311 (
            .O(N__10059),
            .I(N__10050));
    InMux I__2310 (
            .O(N__10058),
            .I(N__10047));
    LocalMux I__2309 (
            .O(N__10053),
            .I(N__10044));
    Odrv4 I__2308 (
            .O(N__10050),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    LocalMux I__2307 (
            .O(N__10047),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    Odrv12 I__2306 (
            .O(N__10044),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    InMux I__2305 (
            .O(N__10037),
            .I(N__10027));
    InMux I__2304 (
            .O(N__10036),
            .I(N__10027));
    InMux I__2303 (
            .O(N__10035),
            .I(N__10027));
    InMux I__2302 (
            .O(N__10034),
            .I(N__10024));
    LocalMux I__2301 (
            .O(N__10027),
            .I(N__10020));
    LocalMux I__2300 (
            .O(N__10024),
            .I(N__10017));
    CascadeMux I__2299 (
            .O(N__10023),
            .I(N__10012));
    Span4Mux_v I__2298 (
            .O(N__10020),
            .I(N__10006));
    Span4Mux_v I__2297 (
            .O(N__10017),
            .I(N__10006));
    InMux I__2296 (
            .O(N__10016),
            .I(N__10003));
    InMux I__2295 (
            .O(N__10015),
            .I(N__10000));
    InMux I__2294 (
            .O(N__10012),
            .I(N__9995));
    InMux I__2293 (
            .O(N__10011),
            .I(N__9995));
    Odrv4 I__2292 (
            .O(N__10006),
            .I(\U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_1 ));
    LocalMux I__2291 (
            .O(N__10003),
            .I(\U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_1 ));
    LocalMux I__2290 (
            .O(N__10000),
            .I(\U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_1 ));
    LocalMux I__2289 (
            .O(N__9995),
            .I(\U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_1 ));
    CascadeMux I__2288 (
            .O(N__9986),
            .I(N__9983));
    InMux I__2287 (
            .O(N__9983),
            .I(N__9979));
    CascadeMux I__2286 (
            .O(N__9982),
            .I(N__9976));
    LocalMux I__2285 (
            .O(N__9979),
            .I(N__9973));
    InMux I__2284 (
            .O(N__9976),
            .I(N__9970));
    Span4Mux_h I__2283 (
            .O(N__9973),
            .I(N__9965));
    LocalMux I__2282 (
            .O(N__9970),
            .I(N__9965));
    Span4Mux_h I__2281 (
            .O(N__9965),
            .I(N__9962));
    Odrv4 I__2280 (
            .O(N__9962),
            .I(\U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z5 ));
    CascadeMux I__2279 (
            .O(N__9959),
            .I(N__9953));
    CascadeMux I__2278 (
            .O(N__9958),
            .I(N__9950));
    InMux I__2277 (
            .O(N__9957),
            .I(N__9940));
    InMux I__2276 (
            .O(N__9956),
            .I(N__9940));
    InMux I__2275 (
            .O(N__9953),
            .I(N__9940));
    InMux I__2274 (
            .O(N__9950),
            .I(N__9940));
    InMux I__2273 (
            .O(N__9949),
            .I(N__9937));
    LocalMux I__2272 (
            .O(N__9940),
            .I(N__9927));
    LocalMux I__2271 (
            .O(N__9937),
            .I(N__9927));
    InMux I__2270 (
            .O(N__9936),
            .I(N__9924));
    InMux I__2269 (
            .O(N__9935),
            .I(N__9921));
    InMux I__2268 (
            .O(N__9934),
            .I(N__9918));
    InMux I__2267 (
            .O(N__9933),
            .I(N__9913));
    InMux I__2266 (
            .O(N__9932),
            .I(N__9913));
    Span4Mux_h I__2265 (
            .O(N__9927),
            .I(N__9910));
    LocalMux I__2264 (
            .O(N__9924),
            .I(\U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_0 ));
    LocalMux I__2263 (
            .O(N__9921),
            .I(\U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_0 ));
    LocalMux I__2262 (
            .O(N__9918),
            .I(\U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_0 ));
    LocalMux I__2261 (
            .O(N__9913),
            .I(\U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_0 ));
    Odrv4 I__2260 (
            .O(N__9910),
            .I(\U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_0 ));
    IoInMux I__2259 (
            .O(N__9899),
            .I(N__9896));
    LocalMux I__2258 (
            .O(N__9896),
            .I(N__9893));
    Span4Mux_s1_v I__2257 (
            .O(N__9893),
            .I(N__9890));
    Span4Mux_v I__2256 (
            .O(N__9890),
            .I(N__9887));
    Span4Mux_v I__2255 (
            .O(N__9887),
            .I(N__9884));
    Span4Mux_v I__2254 (
            .O(N__9884),
            .I(N__9880));
    InMux I__2253 (
            .O(N__9883),
            .I(N__9877));
    Odrv4 I__2252 (
            .O(N__9880),
            .I(ROMENn_c));
    LocalMux I__2251 (
            .O(N__9877),
            .I(ROMENn_c));
    CascadeMux I__2250 (
            .O(N__9872),
            .I(N__9866));
    InMux I__2249 (
            .O(N__9871),
            .I(N__9861));
    InMux I__2248 (
            .O(N__9870),
            .I(N__9858));
    InMux I__2247 (
            .O(N__9869),
            .I(N__9855));
    InMux I__2246 (
            .O(N__9866),
            .I(N__9852));
    InMux I__2245 (
            .O(N__9865),
            .I(N__9847));
    InMux I__2244 (
            .O(N__9864),
            .I(N__9847));
    LocalMux I__2243 (
            .O(N__9861),
            .I(N__9843));
    LocalMux I__2242 (
            .O(N__9858),
            .I(N__9834));
    LocalMux I__2241 (
            .O(N__9855),
            .I(N__9827));
    LocalMux I__2240 (
            .O(N__9852),
            .I(N__9815));
    LocalMux I__2239 (
            .O(N__9847),
            .I(N__9812));
    ClkMux I__2238 (
            .O(N__9846),
            .I(N__9761));
    Glb2LocalMux I__2237 (
            .O(N__9843),
            .I(N__9761));
    ClkMux I__2236 (
            .O(N__9842),
            .I(N__9761));
    ClkMux I__2235 (
            .O(N__9841),
            .I(N__9761));
    ClkMux I__2234 (
            .O(N__9840),
            .I(N__9761));
    ClkMux I__2233 (
            .O(N__9839),
            .I(N__9761));
    ClkMux I__2232 (
            .O(N__9838),
            .I(N__9761));
    ClkMux I__2231 (
            .O(N__9837),
            .I(N__9761));
    Glb2LocalMux I__2230 (
            .O(N__9834),
            .I(N__9761));
    ClkMux I__2229 (
            .O(N__9833),
            .I(N__9761));
    ClkMux I__2228 (
            .O(N__9832),
            .I(N__9761));
    ClkMux I__2227 (
            .O(N__9831),
            .I(N__9761));
    ClkMux I__2226 (
            .O(N__9830),
            .I(N__9761));
    Glb2LocalMux I__2225 (
            .O(N__9827),
            .I(N__9761));
    ClkMux I__2224 (
            .O(N__9826),
            .I(N__9761));
    ClkMux I__2223 (
            .O(N__9825),
            .I(N__9761));
    ClkMux I__2222 (
            .O(N__9824),
            .I(N__9761));
    ClkMux I__2221 (
            .O(N__9823),
            .I(N__9761));
    ClkMux I__2220 (
            .O(N__9822),
            .I(N__9761));
    ClkMux I__2219 (
            .O(N__9821),
            .I(N__9761));
    ClkMux I__2218 (
            .O(N__9820),
            .I(N__9761));
    ClkMux I__2217 (
            .O(N__9819),
            .I(N__9761));
    ClkMux I__2216 (
            .O(N__9818),
            .I(N__9761));
    Glb2LocalMux I__2215 (
            .O(N__9815),
            .I(N__9761));
    Glb2LocalMux I__2214 (
            .O(N__9812),
            .I(N__9761));
    GlobalMux I__2213 (
            .O(N__9761),
            .I(N__9758));
    gio2CtrlBuf I__2212 (
            .O(N__9758),
            .I(CLK40_IN_c_g));
    InMux I__2211 (
            .O(N__9755),
            .I(N__9752));
    LocalMux I__2210 (
            .O(N__9752),
            .I(N__9740));
    SRMux I__2209 (
            .O(N__9751),
            .I(N__9692));
    SRMux I__2208 (
            .O(N__9750),
            .I(N__9692));
    SRMux I__2207 (
            .O(N__9749),
            .I(N__9692));
    SRMux I__2206 (
            .O(N__9748),
            .I(N__9692));
    SRMux I__2205 (
            .O(N__9747),
            .I(N__9692));
    SRMux I__2204 (
            .O(N__9746),
            .I(N__9692));
    SRMux I__2203 (
            .O(N__9745),
            .I(N__9692));
    SRMux I__2202 (
            .O(N__9744),
            .I(N__9692));
    SRMux I__2201 (
            .O(N__9743),
            .I(N__9692));
    Glb2LocalMux I__2200 (
            .O(N__9740),
            .I(N__9692));
    SRMux I__2199 (
            .O(N__9739),
            .I(N__9692));
    SRMux I__2198 (
            .O(N__9738),
            .I(N__9692));
    SRMux I__2197 (
            .O(N__9737),
            .I(N__9692));
    SRMux I__2196 (
            .O(N__9736),
            .I(N__9692));
    SRMux I__2195 (
            .O(N__9735),
            .I(N__9692));
    SRMux I__2194 (
            .O(N__9734),
            .I(N__9692));
    SRMux I__2193 (
            .O(N__9733),
            .I(N__9692));
    SRMux I__2192 (
            .O(N__9732),
            .I(N__9692));
    SRMux I__2191 (
            .O(N__9731),
            .I(N__9692));
    GlobalMux I__2190 (
            .O(N__9692),
            .I(N__9689));
    gio2CtrlBuf I__2189 (
            .O(N__9689),
            .I(RESETn_c_i_g));
    InMux I__2188 (
            .O(N__9686),
            .I(N__9683));
    LocalMux I__2187 (
            .O(N__9683),
            .I(\U409_TICK.TICK603_11 ));
    InMux I__2186 (
            .O(N__9680),
            .I(bfn_15_7_0_));
    InMux I__2185 (
            .O(N__9677),
            .I(\U409_TICK.un2_COUNTER50_1_cry_9 ));
    InMux I__2184 (
            .O(N__9674),
            .I(\U409_TICK.un2_COUNTER50_1_cry_10 ));
    InMux I__2183 (
            .O(N__9671),
            .I(\U409_TICK.un2_COUNTER50_1_cry_11 ));
    InMux I__2182 (
            .O(N__9668),
            .I(\U409_TICK.un2_COUNTER50_1_cry_12 ));
    InMux I__2181 (
            .O(N__9665),
            .I(\U409_TICK.un2_COUNTER50_1_cry_13 ));
    InMux I__2180 (
            .O(N__9662),
            .I(\U409_TICK.un2_COUNTER50_1_cry_14 ));
    InMux I__2179 (
            .O(N__9659),
            .I(\U409_TICK.un2_COUNTER50_1_cry_15 ));
    InMux I__2178 (
            .O(N__9656),
            .I(N__9652));
    InMux I__2177 (
            .O(N__9655),
            .I(N__9649));
    LocalMux I__2176 (
            .O(N__9652),
            .I(N__9646));
    LocalMux I__2175 (
            .O(N__9649),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    Odrv4 I__2174 (
            .O(N__9646),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    IoInMux I__2173 (
            .O(N__9641),
            .I(N__9638));
    LocalMux I__2172 (
            .O(N__9638),
            .I(N__9635));
    IoSpan4Mux I__2171 (
            .O(N__9635),
            .I(N__9632));
    Span4Mux_s0_v I__2170 (
            .O(N__9632),
            .I(N__9629));
    Sp12to4 I__2169 (
            .O(N__9629),
            .I(N__9624));
    InMux I__2168 (
            .O(N__9628),
            .I(N__9621));
    CascadeMux I__2167 (
            .O(N__9627),
            .I(N__9617));
    Span12Mux_s11_v I__2166 (
            .O(N__9624),
            .I(N__9614));
    LocalMux I__2165 (
            .O(N__9621),
            .I(N__9611));
    InMux I__2164 (
            .O(N__9620),
            .I(N__9606));
    InMux I__2163 (
            .O(N__9617),
            .I(N__9606));
    Odrv12 I__2162 (
            .O(N__9614),
            .I(CLK_CIA_c));
    Odrv4 I__2161 (
            .O(N__9611),
            .I(CLK_CIA_c));
    LocalMux I__2160 (
            .O(N__9606),
            .I(CLK_CIA_c));
    InMux I__2159 (
            .O(N__9599),
            .I(N__9594));
    InMux I__2158 (
            .O(N__9598),
            .I(N__9589));
    InMux I__2157 (
            .O(N__9597),
            .I(N__9589));
    LocalMux I__2156 (
            .O(N__9594),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    LocalMux I__2155 (
            .O(N__9589),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    InMux I__2154 (
            .O(N__9584),
            .I(N__9579));
    InMux I__2153 (
            .O(N__9583),
            .I(N__9576));
    InMux I__2152 (
            .O(N__9582),
            .I(N__9573));
    LocalMux I__2151 (
            .O(N__9579),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    LocalMux I__2150 (
            .O(N__9576),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    LocalMux I__2149 (
            .O(N__9573),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    InMux I__2148 (
            .O(N__9566),
            .I(N__9562));
    InMux I__2147 (
            .O(N__9565),
            .I(N__9559));
    LocalMux I__2146 (
            .O(N__9562),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    LocalMux I__2145 (
            .O(N__9559),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    InMux I__2144 (
            .O(N__9554),
            .I(\U409_TICK.un2_COUNTER50_1_cry_1 ));
    InMux I__2143 (
            .O(N__9551),
            .I(\U409_TICK.un2_COUNTER50_1_cry_2 ));
    InMux I__2142 (
            .O(N__9548),
            .I(\U409_TICK.un2_COUNTER50_1_cry_3 ));
    InMux I__2141 (
            .O(N__9545),
            .I(\U409_TICK.un2_COUNTER50_1_cry_4 ));
    CascadeMux I__2140 (
            .O(N__9542),
            .I(N__9539));
    InMux I__2139 (
            .O(N__9539),
            .I(N__9536));
    LocalMux I__2138 (
            .O(N__9536),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ));
    InMux I__2137 (
            .O(N__9533),
            .I(\U409_TICK.un2_COUNTER50_1_cry_5 ));
    InMux I__2136 (
            .O(N__9530),
            .I(\U409_TICK.un2_COUNTER50_1_cry_6 ));
    CascadeMux I__2135 (
            .O(N__9527),
            .I(N__9524));
    InMux I__2134 (
            .O(N__9524),
            .I(N__9520));
    InMux I__2133 (
            .O(N__9523),
            .I(N__9517));
    LocalMux I__2132 (
            .O(N__9520),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    LocalMux I__2131 (
            .O(N__9517),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    InMux I__2130 (
            .O(N__9512),
            .I(\U409_TICK.un2_COUNTER50_1_cry_7 ));
    CascadeMux I__2129 (
            .O(N__9509),
            .I(N__9505));
    InMux I__2128 (
            .O(N__9508),
            .I(N__9500));
    InMux I__2127 (
            .O(N__9505),
            .I(N__9500));
    LocalMux I__2126 (
            .O(N__9500),
            .I(N__9497));
    Span4Mux_v I__2125 (
            .O(N__9497),
            .I(N__9494));
    Sp12to4 I__2124 (
            .O(N__9494),
            .I(N__9491));
    Span12Mux_v I__2123 (
            .O(N__9491),
            .I(N__9488));
    Span12Mux_h I__2122 (
            .O(N__9488),
            .I(N__9485));
    Odrv12 I__2121 (
            .O(N__9485),
            .I(ROM_DELAY_c_0));
    InMux I__2120 (
            .O(N__9482),
            .I(N__9475));
    InMux I__2119 (
            .O(N__9481),
            .I(N__9475));
    InMux I__2118 (
            .O(N__9480),
            .I(N__9472));
    LocalMux I__2117 (
            .O(N__9475),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__2116 (
            .O(N__9472),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    CascadeMux I__2115 (
            .O(N__9467),
            .I(N__9464));
    InMux I__2114 (
            .O(N__9464),
            .I(N__9458));
    InMux I__2113 (
            .O(N__9463),
            .I(N__9458));
    LocalMux I__2112 (
            .O(N__9458),
            .I(N__9455));
    Span4Mux_h I__2111 (
            .O(N__9455),
            .I(N__9452));
    Span4Mux_v I__2110 (
            .O(N__9452),
            .I(N__9449));
    Sp12to4 I__2109 (
            .O(N__9449),
            .I(N__9446));
    Span12Mux_h I__2108 (
            .O(N__9446),
            .I(N__9443));
    Span12Mux_v I__2107 (
            .O(N__9443),
            .I(N__9440));
    Odrv12 I__2106 (
            .O(N__9440),
            .I(ROM_DELAY_c_1));
    InMux I__2105 (
            .O(N__9437),
            .I(N__9432));
    InMux I__2104 (
            .O(N__9436),
            .I(N__9427));
    InMux I__2103 (
            .O(N__9435),
            .I(N__9427));
    LocalMux I__2102 (
            .O(N__9432),
            .I(N__9424));
    LocalMux I__2101 (
            .O(N__9427),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    Odrv4 I__2100 (
            .O(N__9424),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    InMux I__2099 (
            .O(N__9419),
            .I(N__9416));
    LocalMux I__2098 (
            .O(N__9416),
            .I(\U409_TRANSFER_ACK.N_19_mux ));
    IoInMux I__2097 (
            .O(N__9413),
            .I(N__9410));
    LocalMux I__2096 (
            .O(N__9410),
            .I(N__9407));
    IoSpan4Mux I__2095 (
            .O(N__9407),
            .I(N__9404));
    Span4Mux_s2_v I__2094 (
            .O(N__9404),
            .I(N__9401));
    Sp12to4 I__2093 (
            .O(N__9401),
            .I(N__9398));
    Span12Mux_s10_v I__2092 (
            .O(N__9398),
            .I(N__9394));
    InMux I__2091 (
            .O(N__9397),
            .I(N__9391));
    Odrv12 I__2090 (
            .O(N__9394),
            .I(TICK60_c));
    LocalMux I__2089 (
            .O(N__9391),
            .I(TICK60_c));
    CascadeMux I__2088 (
            .O(N__9386),
            .I(\U409_TICK.TICK603_9_cascade_ ));
    IoInMux I__2087 (
            .O(N__9383),
            .I(N__9380));
    LocalMux I__2086 (
            .O(N__9380),
            .I(N__9377));
    Span4Mux_s1_v I__2085 (
            .O(N__9377),
            .I(N__9374));
    Sp12to4 I__2084 (
            .O(N__9374),
            .I(N__9371));
    Span12Mux_h I__2083 (
            .O(N__9371),
            .I(N__9367));
    InMux I__2082 (
            .O(N__9370),
            .I(N__9364));
    Odrv12 I__2081 (
            .O(N__9367),
            .I(TICK50_c));
    LocalMux I__2080 (
            .O(N__9364),
            .I(TICK50_c));
    CascadeMux I__2079 (
            .O(N__9359),
            .I(\U409_TICK.TICK603_8_cascade_ ));
    CascadeMux I__2078 (
            .O(N__9356),
            .I(\U409_TICK.TICK603_14_cascade_ ));
    InMux I__2077 (
            .O(N__9353),
            .I(N__9350));
    LocalMux I__2076 (
            .O(N__9350),
            .I(\U409_TRANSFER_ACK.N_17_mux ));
    CascadeMux I__2075 (
            .O(N__9347),
            .I(\U409_TRANSFER_ACK.N_17_mux_cascade_ ));
    InMux I__2074 (
            .O(N__9344),
            .I(N__9341));
    LocalMux I__2073 (
            .O(N__9341),
            .I(\U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0 ));
    InMux I__2072 (
            .O(N__9338),
            .I(N__9335));
    LocalMux I__2071 (
            .O(N__9335),
            .I(\U409_TRANSFER_ACK.N_3_0 ));
    InMux I__2070 (
            .O(N__9332),
            .I(N__9326));
    InMux I__2069 (
            .O(N__9331),
            .I(N__9323));
    InMux I__2068 (
            .O(N__9330),
            .I(N__9318));
    InMux I__2067 (
            .O(N__9329),
            .I(N__9318));
    LocalMux I__2066 (
            .O(N__9326),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__2065 (
            .O(N__9323),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__2064 (
            .O(N__9318),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    InMux I__2063 (
            .O(N__9311),
            .I(N__9306));
    InMux I__2062 (
            .O(N__9310),
            .I(N__9301));
    InMux I__2061 (
            .O(N__9309),
            .I(N__9301));
    LocalMux I__2060 (
            .O(N__9306),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    LocalMux I__2059 (
            .O(N__9301),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    CascadeMux I__2058 (
            .O(N__9296),
            .I(\U409_TRANSFER_ACK.N_3_0_cascade_ ));
    InMux I__2057 (
            .O(N__9293),
            .I(N__9287));
    InMux I__2056 (
            .O(N__9292),
            .I(N__9284));
    InMux I__2055 (
            .O(N__9291),
            .I(N__9279));
    InMux I__2054 (
            .O(N__9290),
            .I(N__9279));
    LocalMux I__2053 (
            .O(N__9287),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__2052 (
            .O(N__9284),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__2051 (
            .O(N__9279),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    InMux I__2050 (
            .O(N__9272),
            .I(N__9269));
    LocalMux I__2049 (
            .O(N__9269),
            .I(\U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0 ));
    InMux I__2048 (
            .O(N__9266),
            .I(N__9260));
    InMux I__2047 (
            .O(N__9265),
            .I(N__9260));
    LocalMux I__2046 (
            .O(N__9260),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    InMux I__2045 (
            .O(N__9257),
            .I(N__9253));
    InMux I__2044 (
            .O(N__9256),
            .I(N__9250));
    LocalMux I__2043 (
            .O(N__9253),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__2042 (
            .O(N__9250),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    InMux I__2041 (
            .O(N__9245),
            .I(N__9241));
    InMux I__2040 (
            .O(N__9244),
            .I(N__9238));
    LocalMux I__2039 (
            .O(N__9241),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__2038 (
            .O(N__9238),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    CascadeMux I__2037 (
            .O(N__9233),
            .I(\U409_TRANSFER_ACK.N_7_cascade_ ));
    InMux I__2036 (
            .O(N__9230),
            .I(N__9227));
    LocalMux I__2035 (
            .O(N__9227),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_3 ));
    InMux I__2034 (
            .O(N__9224),
            .I(N__9221));
    LocalMux I__2033 (
            .O(N__9221),
            .I(N__9218));
    Span4Mux_v I__2032 (
            .O(N__9218),
            .I(N__9215));
    Odrv4 I__2031 (
            .O(N__9215),
            .I(AC_TACK));
    InMux I__2030 (
            .O(N__9212),
            .I(N__9208));
    InMux I__2029 (
            .O(N__9211),
            .I(N__9205));
    LocalMux I__2028 (
            .O(N__9208),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    LocalMux I__2027 (
            .O(N__9205),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    InMux I__2026 (
            .O(N__9200),
            .I(N__9197));
    LocalMux I__2025 (
            .O(N__9197),
            .I(\U409_TRANSFER_ACK.TACK_START_2_1 ));
    InMux I__2024 (
            .O(N__9194),
            .I(N__9189));
    CascadeMux I__2023 (
            .O(N__9193),
            .I(N__9186));
    CascadeMux I__2022 (
            .O(N__9192),
            .I(N__9182));
    LocalMux I__2021 (
            .O(N__9189),
            .I(N__9179));
    InMux I__2020 (
            .O(N__9186),
            .I(N__9174));
    InMux I__2019 (
            .O(N__9185),
            .I(N__9174));
    InMux I__2018 (
            .O(N__9182),
            .I(N__9171));
    Span4Mux_v I__2017 (
            .O(N__9179),
            .I(N__9166));
    LocalMux I__2016 (
            .O(N__9174),
            .I(N__9166));
    LocalMux I__2015 (
            .O(N__9171),
            .I(\U409_TRANSFER_ACK.TACK_STARTZ0 ));
    Odrv4 I__2014 (
            .O(N__9166),
            .I(\U409_TRANSFER_ACK.TACK_STARTZ0 ));
    ClkMux I__2013 (
            .O(N__9161),
            .I(N__9134));
    ClkMux I__2012 (
            .O(N__9160),
            .I(N__9134));
    ClkMux I__2011 (
            .O(N__9159),
            .I(N__9134));
    ClkMux I__2010 (
            .O(N__9158),
            .I(N__9134));
    ClkMux I__2009 (
            .O(N__9157),
            .I(N__9134));
    ClkMux I__2008 (
            .O(N__9156),
            .I(N__9134));
    ClkMux I__2007 (
            .O(N__9155),
            .I(N__9134));
    ClkMux I__2006 (
            .O(N__9154),
            .I(N__9134));
    ClkMux I__2005 (
            .O(N__9153),
            .I(N__9134));
    GlobalMux I__2004 (
            .O(N__9134),
            .I(CLK80_OUT));
    InMux I__2003 (
            .O(N__9131),
            .I(N__9128));
    LocalMux I__2002 (
            .O(N__9128),
            .I(N__9125));
    Odrv4 I__2001 (
            .O(N__9125),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_0 ));
    IoInMux I__2000 (
            .O(N__9122),
            .I(N__9118));
    IoInMux I__1999 (
            .O(N__9121),
            .I(N__9115));
    LocalMux I__1998 (
            .O(N__9118),
            .I(N__9112));
    LocalMux I__1997 (
            .O(N__9115),
            .I(N__9109));
    IoSpan4Mux I__1996 (
            .O(N__9112),
            .I(N__9103));
    IoSpan4Mux I__1995 (
            .O(N__9109),
            .I(N__9103));
    IoInMux I__1994 (
            .O(N__9108),
            .I(N__9100));
    Span4Mux_s3_v I__1993 (
            .O(N__9103),
            .I(N__9097));
    LocalMux I__1992 (
            .O(N__9100),
            .I(N__9093));
    Span4Mux_v I__1991 (
            .O(N__9097),
            .I(N__9090));
    InMux I__1990 (
            .O(N__9096),
            .I(N__9087));
    Span12Mux_s7_v I__1989 (
            .O(N__9093),
            .I(N__9082));
    Sp12to4 I__1988 (
            .O(N__9090),
            .I(N__9082));
    LocalMux I__1987 (
            .O(N__9087),
            .I(N__9079));
    Span12Mux_h I__1986 (
            .O(N__9082),
            .I(N__9075));
    Span4Mux_v I__1985 (
            .O(N__9079),
            .I(N__9072));
    InMux I__1984 (
            .O(N__9078),
            .I(N__9069));
    Odrv12 I__1983 (
            .O(N__9075),
            .I(TACK_EN));
    Odrv4 I__1982 (
            .O(N__9072),
            .I(TACK_EN));
    LocalMux I__1981 (
            .O(N__9069),
            .I(TACK_EN));
    InMux I__1980 (
            .O(N__9062),
            .I(N__9059));
    LocalMux I__1979 (
            .O(N__9059),
            .I(N__9055));
    InMux I__1978 (
            .O(N__9058),
            .I(N__9052));
    Span4Mux_v I__1977 (
            .O(N__9055),
            .I(N__9049));
    LocalMux I__1976 (
            .O(N__9052),
            .I(N__9042));
    Span4Mux_h I__1975 (
            .O(N__9049),
            .I(N__9037));
    CascadeMux I__1974 (
            .O(N__9048),
            .I(N__9031));
    CascadeMux I__1973 (
            .O(N__9047),
            .I(N__9028));
    InMux I__1972 (
            .O(N__9046),
            .I(N__9016));
    InMux I__1971 (
            .O(N__9045),
            .I(N__9016));
    Span4Mux_v I__1970 (
            .O(N__9042),
            .I(N__9013));
    InMux I__1969 (
            .O(N__9041),
            .I(N__9008));
    InMux I__1968 (
            .O(N__9040),
            .I(N__9008));
    Span4Mux_h I__1967 (
            .O(N__9037),
            .I(N__9004));
    InMux I__1966 (
            .O(N__9036),
            .I(N__9001));
    InMux I__1965 (
            .O(N__9035),
            .I(N__8998));
    InMux I__1964 (
            .O(N__9034),
            .I(N__8985));
    InMux I__1963 (
            .O(N__9031),
            .I(N__8985));
    InMux I__1962 (
            .O(N__9028),
            .I(N__8985));
    InMux I__1961 (
            .O(N__9027),
            .I(N__8985));
    InMux I__1960 (
            .O(N__9026),
            .I(N__8985));
    InMux I__1959 (
            .O(N__9025),
            .I(N__8985));
    CascadeMux I__1958 (
            .O(N__9024),
            .I(N__8980));
    CascadeMux I__1957 (
            .O(N__9023),
            .I(N__8977));
    CascadeMux I__1956 (
            .O(N__9022),
            .I(N__8973));
    CascadeMux I__1955 (
            .O(N__9021),
            .I(N__8970));
    LocalMux I__1954 (
            .O(N__9016),
            .I(N__8966));
    Span4Mux_v I__1953 (
            .O(N__9013),
            .I(N__8961));
    LocalMux I__1952 (
            .O(N__9008),
            .I(N__8961));
    InMux I__1951 (
            .O(N__9007),
            .I(N__8958));
    Span4Mux_v I__1950 (
            .O(N__9004),
            .I(N__8949));
    LocalMux I__1949 (
            .O(N__9001),
            .I(N__8949));
    LocalMux I__1948 (
            .O(N__8998),
            .I(N__8949));
    LocalMux I__1947 (
            .O(N__8985),
            .I(N__8949));
    InMux I__1946 (
            .O(N__8984),
            .I(N__8945));
    InMux I__1945 (
            .O(N__8983),
            .I(N__8940));
    InMux I__1944 (
            .O(N__8980),
            .I(N__8940));
    InMux I__1943 (
            .O(N__8977),
            .I(N__8937));
    InMux I__1942 (
            .O(N__8976),
            .I(N__8934));
    InMux I__1941 (
            .O(N__8973),
            .I(N__8929));
    InMux I__1940 (
            .O(N__8970),
            .I(N__8929));
    InMux I__1939 (
            .O(N__8969),
            .I(N__8925));
    Span4Mux_h I__1938 (
            .O(N__8966),
            .I(N__8918));
    Span4Mux_h I__1937 (
            .O(N__8961),
            .I(N__8918));
    LocalMux I__1936 (
            .O(N__8958),
            .I(N__8918));
    Span4Mux_v I__1935 (
            .O(N__8949),
            .I(N__8915));
    InMux I__1934 (
            .O(N__8948),
            .I(N__8912));
    LocalMux I__1933 (
            .O(N__8945),
            .I(N__8901));
    LocalMux I__1932 (
            .O(N__8940),
            .I(N__8901));
    LocalMux I__1931 (
            .O(N__8937),
            .I(N__8901));
    LocalMux I__1930 (
            .O(N__8934),
            .I(N__8901));
    LocalMux I__1929 (
            .O(N__8929),
            .I(N__8901));
    InMux I__1928 (
            .O(N__8928),
            .I(N__8898));
    LocalMux I__1927 (
            .O(N__8925),
            .I(N__8895));
    Span4Mux_v I__1926 (
            .O(N__8918),
            .I(N__8892));
    Span4Mux_h I__1925 (
            .O(N__8915),
            .I(N__8887));
    LocalMux I__1924 (
            .O(N__8912),
            .I(N__8887));
    Span4Mux_v I__1923 (
            .O(N__8901),
            .I(N__8882));
    LocalMux I__1922 (
            .O(N__8898),
            .I(N__8882));
    Span12Mux_v I__1921 (
            .O(N__8895),
            .I(N__8879));
    Sp12to4 I__1920 (
            .O(N__8892),
            .I(N__8876));
    Span4Mux_v I__1919 (
            .O(N__8887),
            .I(N__8871));
    Span4Mux_v I__1918 (
            .O(N__8882),
            .I(N__8871));
    Span12Mux_v I__1917 (
            .O(N__8879),
            .I(N__8868));
    Span12Mux_h I__1916 (
            .O(N__8876),
            .I(N__8865));
    Sp12to4 I__1915 (
            .O(N__8871),
            .I(N__8862));
    Span12Mux_h I__1914 (
            .O(N__8868),
            .I(N__8857));
    Span12Mux_v I__1913 (
            .O(N__8865),
            .I(N__8857));
    Span12Mux_h I__1912 (
            .O(N__8862),
            .I(N__8854));
    Odrv12 I__1911 (
            .O(N__8857),
            .I(RESETn_c));
    Odrv12 I__1910 (
            .O(N__8854),
            .I(RESETn_c));
    SRMux I__1909 (
            .O(N__8849),
            .I(N__8846));
    LocalMux I__1908 (
            .O(N__8846),
            .I(N__8843));
    Span4Mux_v I__1907 (
            .O(N__8843),
            .I(N__8840));
    Span4Mux_v I__1906 (
            .O(N__8840),
            .I(N__8837));
    Odrv4 I__1905 (
            .O(N__8837),
            .I(\U409_TRANSFER_ACK.TACK_RST_0_i ));
    InMux I__1904 (
            .O(N__8834),
            .I(N__8829));
    InMux I__1903 (
            .O(N__8833),
            .I(N__8825));
    InMux I__1902 (
            .O(N__8832),
            .I(N__8822));
    LocalMux I__1901 (
            .O(N__8829),
            .I(N__8819));
    InMux I__1900 (
            .O(N__8828),
            .I(N__8816));
    LocalMux I__1899 (
            .O(N__8825),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__1898 (
            .O(N__8822),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    Odrv12 I__1897 (
            .O(N__8819),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__1896 (
            .O(N__8816),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    InMux I__1895 (
            .O(N__8807),
            .I(N__8803));
    CascadeMux I__1894 (
            .O(N__8806),
            .I(N__8796));
    LocalMux I__1893 (
            .O(N__8803),
            .I(N__8793));
    InMux I__1892 (
            .O(N__8802),
            .I(N__8788));
    InMux I__1891 (
            .O(N__8801),
            .I(N__8788));
    InMux I__1890 (
            .O(N__8800),
            .I(N__8783));
    InMux I__1889 (
            .O(N__8799),
            .I(N__8783));
    InMux I__1888 (
            .O(N__8796),
            .I(N__8780));
    Odrv4 I__1887 (
            .O(N__8793),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1886 (
            .O(N__8788),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1885 (
            .O(N__8783),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1884 (
            .O(N__8780),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    CascadeMux I__1883 (
            .O(N__8771),
            .I(N__8768));
    InMux I__1882 (
            .O(N__8768),
            .I(N__8764));
    InMux I__1881 (
            .O(N__8767),
            .I(N__8759));
    LocalMux I__1880 (
            .O(N__8764),
            .I(N__8756));
    InMux I__1879 (
            .O(N__8763),
            .I(N__8753));
    InMux I__1878 (
            .O(N__8762),
            .I(N__8750));
    LocalMux I__1877 (
            .O(N__8759),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    Odrv4 I__1876 (
            .O(N__8756),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    LocalMux I__1875 (
            .O(N__8753),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    LocalMux I__1874 (
            .O(N__8750),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    InMux I__1873 (
            .O(N__8741),
            .I(N__8738));
    LocalMux I__1872 (
            .O(N__8738),
            .I(N__8731));
    InMux I__1871 (
            .O(N__8737),
            .I(N__8723));
    InMux I__1870 (
            .O(N__8736),
            .I(N__8723));
    InMux I__1869 (
            .O(N__8735),
            .I(N__8723));
    InMux I__1868 (
            .O(N__8734),
            .I(N__8720));
    Span4Mux_v I__1867 (
            .O(N__8731),
            .I(N__8717));
    InMux I__1866 (
            .O(N__8730),
            .I(N__8714));
    LocalMux I__1865 (
            .O(N__8723),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__1864 (
            .O(N__8720),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    Odrv4 I__1863 (
            .O(N__8717),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__1862 (
            .O(N__8714),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    CascadeMux I__1861 (
            .O(N__8705),
            .I(\U409_CIA.CLK_CIA6_3_cascade_ ));
    InMux I__1860 (
            .O(N__8702),
            .I(N__8697));
    CascadeMux I__1859 (
            .O(N__8701),
            .I(N__8692));
    CascadeMux I__1858 (
            .O(N__8700),
            .I(N__8689));
    LocalMux I__1857 (
            .O(N__8697),
            .I(N__8686));
    InMux I__1856 (
            .O(N__8696),
            .I(N__8683));
    InMux I__1855 (
            .O(N__8695),
            .I(N__8678));
    InMux I__1854 (
            .O(N__8692),
            .I(N__8678));
    InMux I__1853 (
            .O(N__8689),
            .I(N__8675));
    Odrv12 I__1852 (
            .O(N__8686),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__1851 (
            .O(N__8683),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__1850 (
            .O(N__8678),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__1849 (
            .O(N__8675),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    InMux I__1848 (
            .O(N__8666),
            .I(N__8662));
    CascadeMux I__1847 (
            .O(N__8665),
            .I(N__8658));
    LocalMux I__1846 (
            .O(N__8662),
            .I(N__8654));
    InMux I__1845 (
            .O(N__8661),
            .I(N__8651));
    InMux I__1844 (
            .O(N__8658),
            .I(N__8648));
    InMux I__1843 (
            .O(N__8657),
            .I(N__8645));
    Odrv4 I__1842 (
            .O(N__8654),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__1841 (
            .O(N__8651),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__1840 (
            .O(N__8648),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__1839 (
            .O(N__8645),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    InMux I__1838 (
            .O(N__8636),
            .I(N__8633));
    LocalMux I__1837 (
            .O(N__8633),
            .I(N__8626));
    InMux I__1836 (
            .O(N__8632),
            .I(N__8623));
    InMux I__1835 (
            .O(N__8631),
            .I(N__8620));
    InMux I__1834 (
            .O(N__8630),
            .I(N__8615));
    InMux I__1833 (
            .O(N__8629),
            .I(N__8615));
    Odrv4 I__1832 (
            .O(N__8626),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__1831 (
            .O(N__8623),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__1830 (
            .O(N__8620),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__1829 (
            .O(N__8615),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    InMux I__1828 (
            .O(N__8606),
            .I(N__8603));
    LocalMux I__1827 (
            .O(N__8603),
            .I(N__8597));
    InMux I__1826 (
            .O(N__8602),
            .I(N__8594));
    InMux I__1825 (
            .O(N__8601),
            .I(N__8591));
    InMux I__1824 (
            .O(N__8600),
            .I(N__8588));
    Odrv4 I__1823 (
            .O(N__8597),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__1822 (
            .O(N__8594),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__1821 (
            .O(N__8591),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__1820 (
            .O(N__8588),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    InMux I__1819 (
            .O(N__8579),
            .I(N__8576));
    LocalMux I__1818 (
            .O(N__8576),
            .I(\U409_CIA.CLK_CIA_r_1_0 ));
    CascadeMux I__1817 (
            .O(N__8573),
            .I(N__8569));
    CascadeMux I__1816 (
            .O(N__8572),
            .I(N__8565));
    InMux I__1815 (
            .O(N__8569),
            .I(N__8562));
    InMux I__1814 (
            .O(N__8568),
            .I(N__8559));
    InMux I__1813 (
            .O(N__8565),
            .I(N__8556));
    LocalMux I__1812 (
            .O(N__8562),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__1811 (
            .O(N__8559),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__1810 (
            .O(N__8556),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    InMux I__1809 (
            .O(N__8549),
            .I(N__8546));
    LocalMux I__1808 (
            .O(N__8546),
            .I(N__8541));
    InMux I__1807 (
            .O(N__8545),
            .I(N__8538));
    InMux I__1806 (
            .O(N__8544),
            .I(N__8535));
    Odrv4 I__1805 (
            .O(N__8541),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__1804 (
            .O(N__8538),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__1803 (
            .O(N__8535),
            .I(\U409_CIA.VMAZ0 ));
    InMux I__1802 (
            .O(N__8528),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_0 ));
    InMux I__1801 (
            .O(N__8525),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_1 ));
    InMux I__1800 (
            .O(N__8522),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_2 ));
    InMux I__1799 (
            .O(N__8519),
            .I(N__8516));
    LocalMux I__1798 (
            .O(N__8516),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_2 ));
    InMux I__1797 (
            .O(N__8513),
            .I(N__8510));
    LocalMux I__1796 (
            .O(N__8510),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_1 ));
    InMux I__1795 (
            .O(N__8507),
            .I(N__8503));
    InMux I__1794 (
            .O(N__8506),
            .I(N__8500));
    LocalMux I__1793 (
            .O(N__8503),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    LocalMux I__1792 (
            .O(N__8500),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    InMux I__1791 (
            .O(N__8495),
            .I(N__8491));
    InMux I__1790 (
            .O(N__8494),
            .I(N__8488));
    LocalMux I__1789 (
            .O(N__8491),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    LocalMux I__1788 (
            .O(N__8488),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    InMux I__1787 (
            .O(N__8483),
            .I(N__8480));
    LocalMux I__1786 (
            .O(N__8480),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_2 ));
    InMux I__1785 (
            .O(N__8477),
            .I(N__8471));
    InMux I__1784 (
            .O(N__8476),
            .I(N__8471));
    LocalMux I__1783 (
            .O(N__8471),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ));
    CascadeMux I__1782 (
            .O(N__8468),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_cascade_ ));
    IoInMux I__1781 (
            .O(N__8465),
            .I(N__8462));
    LocalMux I__1780 (
            .O(N__8462),
            .I(N__8459));
    Odrv12 I__1779 (
            .O(N__8459),
            .I(RESETn_c_i));
    InMux I__1778 (
            .O(N__8456),
            .I(N__8452));
    CascadeMux I__1777 (
            .O(N__8455),
            .I(N__8448));
    LocalMux I__1776 (
            .O(N__8452),
            .I(N__8445));
    InMux I__1775 (
            .O(N__8451),
            .I(N__8442));
    InMux I__1774 (
            .O(N__8448),
            .I(N__8439));
    Span4Mux_v I__1773 (
            .O(N__8445),
            .I(N__8436));
    LocalMux I__1772 (
            .O(N__8442),
            .I(N__8431));
    LocalMux I__1771 (
            .O(N__8439),
            .I(N__8431));
    Span4Mux_h I__1770 (
            .O(N__8436),
            .I(N__8428));
    Span4Mux_v I__1769 (
            .O(N__8431),
            .I(N__8425));
    Sp12to4 I__1768 (
            .O(N__8428),
            .I(N__8420));
    Sp12to4 I__1767 (
            .O(N__8425),
            .I(N__8420));
    Odrv12 I__1766 (
            .O(N__8420),
            .I(A_c_12));
    IoInMux I__1765 (
            .O(N__8417),
            .I(N__8414));
    LocalMux I__1764 (
            .O(N__8414),
            .I(N__8411));
    IoSpan4Mux I__1763 (
            .O(N__8411),
            .I(N__8408));
    IoSpan4Mux I__1762 (
            .O(N__8408),
            .I(N__8405));
    Sp12to4 I__1761 (
            .O(N__8405),
            .I(N__8402));
    Span12Mux_s7_h I__1760 (
            .O(N__8402),
            .I(N__8399));
    Odrv12 I__1759 (
            .O(N__8399),
            .I(U409_ADDRESS_DECODE_un1_CIACS0n_i));
    InMux I__1758 (
            .O(N__8396),
            .I(N__8392));
    InMux I__1757 (
            .O(N__8395),
            .I(N__8389));
    LocalMux I__1756 (
            .O(N__8392),
            .I(CIA_ENABLE));
    LocalMux I__1755 (
            .O(N__8389),
            .I(CIA_ENABLE));
    InMux I__1754 (
            .O(N__8384),
            .I(N__8380));
    CascadeMux I__1753 (
            .O(N__8383),
            .I(N__8376));
    LocalMux I__1752 (
            .O(N__8380),
            .I(N__8373));
    InMux I__1751 (
            .O(N__8379),
            .I(N__8370));
    InMux I__1750 (
            .O(N__8376),
            .I(N__8367));
    Sp12to4 I__1749 (
            .O(N__8373),
            .I(N__8364));
    LocalMux I__1748 (
            .O(N__8370),
            .I(N__8359));
    LocalMux I__1747 (
            .O(N__8367),
            .I(N__8359));
    Span12Mux_v I__1746 (
            .O(N__8364),
            .I(N__8356));
    Span4Mux_v I__1745 (
            .O(N__8359),
            .I(N__8353));
    Span12Mux_h I__1744 (
            .O(N__8356),
            .I(N__8350));
    Sp12to4 I__1743 (
            .O(N__8353),
            .I(N__8347));
    Odrv12 I__1742 (
            .O(N__8350),
            .I(A_c_13));
    Odrv12 I__1741 (
            .O(N__8347),
            .I(A_c_13));
    IoInMux I__1740 (
            .O(N__8342),
            .I(N__8339));
    LocalMux I__1739 (
            .O(N__8339),
            .I(N__8336));
    IoSpan4Mux I__1738 (
            .O(N__8336),
            .I(N__8333));
    Span4Mux_s1_h I__1737 (
            .O(N__8333),
            .I(N__8330));
    Sp12to4 I__1736 (
            .O(N__8330),
            .I(N__8327));
    Span12Mux_h I__1735 (
            .O(N__8327),
            .I(N__8324));
    Odrv12 I__1734 (
            .O(N__8324),
            .I(U409_ADDRESS_DECODE_un1_CIACS1n_i));
    InMux I__1733 (
            .O(N__8321),
            .I(N__8318));
    LocalMux I__1732 (
            .O(N__8318),
            .I(\U409_TRANSFER_ACK.N_5_0 ));
    InMux I__1731 (
            .O(N__8315),
            .I(N__8304));
    InMux I__1730 (
            .O(N__8314),
            .I(N__8304));
    InMux I__1729 (
            .O(N__8313),
            .I(N__8304));
    InMux I__1728 (
            .O(N__8312),
            .I(N__8301));
    InMux I__1727 (
            .O(N__8311),
            .I(N__8298));
    LocalMux I__1726 (
            .O(N__8304),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__1725 (
            .O(N__8301),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__1724 (
            .O(N__8298),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    InMux I__1723 (
            .O(N__8291),
            .I(N__8285));
    InMux I__1722 (
            .O(N__8290),
            .I(N__8282));
    InMux I__1721 (
            .O(N__8289),
            .I(N__8277));
    InMux I__1720 (
            .O(N__8288),
            .I(N__8277));
    LocalMux I__1719 (
            .O(N__8285),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1718 (
            .O(N__8282),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1717 (
            .O(N__8277),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    CascadeMux I__1716 (
            .O(N__8270),
            .I(N__8264));
    InMux I__1715 (
            .O(N__8269),
            .I(N__8261));
    InMux I__1714 (
            .O(N__8268),
            .I(N__8258));
    InMux I__1713 (
            .O(N__8267),
            .I(N__8253));
    InMux I__1712 (
            .O(N__8264),
            .I(N__8253));
    LocalMux I__1711 (
            .O(N__8261),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__1710 (
            .O(N__8258),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__1709 (
            .O(N__8253),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    InMux I__1708 (
            .O(N__8246),
            .I(N__8241));
    InMux I__1707 (
            .O(N__8245),
            .I(N__8236));
    InMux I__1706 (
            .O(N__8244),
            .I(N__8236));
    LocalMux I__1705 (
            .O(N__8241),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    LocalMux I__1704 (
            .O(N__8236),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    CascadeMux I__1703 (
            .O(N__8231),
            .I(N__8225));
    InMux I__1702 (
            .O(N__8230),
            .I(N__8220));
    InMux I__1701 (
            .O(N__8229),
            .I(N__8220));
    InMux I__1700 (
            .O(N__8228),
            .I(N__8215));
    InMux I__1699 (
            .O(N__8225),
            .I(N__8215));
    LocalMux I__1698 (
            .O(N__8220),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__1697 (
            .O(N__8215),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    CascadeMux I__1696 (
            .O(N__8210),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_ ));
    InMux I__1695 (
            .O(N__8207),
            .I(N__8200));
    InMux I__1694 (
            .O(N__8206),
            .I(N__8191));
    InMux I__1693 (
            .O(N__8205),
            .I(N__8191));
    InMux I__1692 (
            .O(N__8204),
            .I(N__8191));
    InMux I__1691 (
            .O(N__8203),
            .I(N__8191));
    LocalMux I__1690 (
            .O(N__8200),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1689 (
            .O(N__8191),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    CascadeMux I__1688 (
            .O(N__8186),
            .I(N__8181));
    InMux I__1687 (
            .O(N__8185),
            .I(N__8177));
    InMux I__1686 (
            .O(N__8184),
            .I(N__8170));
    InMux I__1685 (
            .O(N__8181),
            .I(N__8170));
    InMux I__1684 (
            .O(N__8180),
            .I(N__8170));
    LocalMux I__1683 (
            .O(N__8177),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1682 (
            .O(N__8170),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    InMux I__1681 (
            .O(N__8165),
            .I(N__8159));
    InMux I__1680 (
            .O(N__8164),
            .I(N__8159));
    LocalMux I__1679 (
            .O(N__8159),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ));
    CascadeMux I__1678 (
            .O(N__8156),
            .I(N__8152));
    InMux I__1677 (
            .O(N__8155),
            .I(N__8149));
    InMux I__1676 (
            .O(N__8152),
            .I(N__8146));
    LocalMux I__1675 (
            .O(N__8149),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ));
    LocalMux I__1674 (
            .O(N__8146),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ));
    InMux I__1673 (
            .O(N__8141),
            .I(N__8134));
    InMux I__1672 (
            .O(N__8140),
            .I(N__8134));
    InMux I__1671 (
            .O(N__8139),
            .I(N__8131));
    LocalMux I__1670 (
            .O(N__8134),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    LocalMux I__1669 (
            .O(N__8131),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    InMux I__1668 (
            .O(N__8126),
            .I(N__8121));
    InMux I__1667 (
            .O(N__8125),
            .I(N__8114));
    InMux I__1666 (
            .O(N__8124),
            .I(N__8111));
    LocalMux I__1665 (
            .O(N__8121),
            .I(N__8108));
    InMux I__1664 (
            .O(N__8120),
            .I(N__8099));
    InMux I__1663 (
            .O(N__8119),
            .I(N__8099));
    InMux I__1662 (
            .O(N__8118),
            .I(N__8099));
    InMux I__1661 (
            .O(N__8117),
            .I(N__8099));
    LocalMux I__1660 (
            .O(N__8114),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1659 (
            .O(N__8111),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    Odrv4 I__1658 (
            .O(N__8108),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1657 (
            .O(N__8099),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    SRMux I__1656 (
            .O(N__8090),
            .I(N__8087));
    LocalMux I__1655 (
            .O(N__8087),
            .I(N__8082));
    SRMux I__1654 (
            .O(N__8086),
            .I(N__8079));
    SRMux I__1653 (
            .O(N__8085),
            .I(N__8076));
    Span4Mux_h I__1652 (
            .O(N__8082),
            .I(N__8073));
    LocalMux I__1651 (
            .O(N__8079),
            .I(N__8070));
    LocalMux I__1650 (
            .O(N__8076),
            .I(N__8067));
    Span4Mux_h I__1649 (
            .O(N__8073),
            .I(N__8062));
    Span4Mux_h I__1648 (
            .O(N__8070),
            .I(N__8062));
    Span4Mux_v I__1647 (
            .O(N__8067),
            .I(N__8059));
    Odrv4 I__1646 (
            .O(N__8062),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    Odrv4 I__1645 (
            .O(N__8059),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    InMux I__1644 (
            .O(N__8054),
            .I(N__8051));
    LocalMux I__1643 (
            .O(N__8051),
            .I(N__8048));
    Span4Mux_v I__1642 (
            .O(N__8048),
            .I(N__8044));
    InMux I__1641 (
            .O(N__8047),
            .I(N__8041));
    Span4Mux_h I__1640 (
            .O(N__8044),
            .I(N__8036));
    LocalMux I__1639 (
            .O(N__8041),
            .I(N__8036));
    Odrv4 I__1638 (
            .O(N__8036),
            .I(U409_ADDRESS_DECODE_un1_RTC_ENn));
    CascadeMux I__1637 (
            .O(N__8033),
            .I(N__8030));
    InMux I__1636 (
            .O(N__8030),
            .I(N__8027));
    LocalMux I__1635 (
            .O(N__8027),
            .I(N__8024));
    Span4Mux_v I__1634 (
            .O(N__8024),
            .I(N__8021));
    Span4Mux_v I__1633 (
            .O(N__8021),
            .I(N__8018));
    Span4Mux_v I__1632 (
            .O(N__8018),
            .I(N__8015));
    Span4Mux_h I__1631 (
            .O(N__8015),
            .I(N__8012));
    Odrv4 I__1630 (
            .O(N__8012),
            .I(U409_ADDRESS_DECODE_AUTOVECTOR_10));
    InMux I__1629 (
            .O(N__8009),
            .I(N__8004));
    InMux I__1628 (
            .O(N__8008),
            .I(N__8001));
    InMux I__1627 (
            .O(N__8007),
            .I(N__7998));
    LocalMux I__1626 (
            .O(N__8004),
            .I(N__7994));
    LocalMux I__1625 (
            .O(N__8001),
            .I(N__7991));
    LocalMux I__1624 (
            .O(N__7998),
            .I(N__7988));
    InMux I__1623 (
            .O(N__7997),
            .I(N__7984));
    Span4Mux_v I__1622 (
            .O(N__7994),
            .I(N__7981));
    Span4Mux_v I__1621 (
            .O(N__7991),
            .I(N__7976));
    Span4Mux_v I__1620 (
            .O(N__7988),
            .I(N__7976));
    InMux I__1619 (
            .O(N__7987),
            .I(N__7973));
    LocalMux I__1618 (
            .O(N__7984),
            .I(N__7964));
    Sp12to4 I__1617 (
            .O(N__7981),
            .I(N__7964));
    Sp12to4 I__1616 (
            .O(N__7976),
            .I(N__7964));
    LocalMux I__1615 (
            .O(N__7973),
            .I(N__7964));
    Span12Mux_h I__1614 (
            .O(N__7964),
            .I(N__7961));
    Span12Mux_v I__1613 (
            .O(N__7961),
            .I(N__7958));
    Odrv12 I__1612 (
            .O(N__7958),
            .I(TSn_c));
    CascadeMux I__1611 (
            .O(N__7955),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_2_cascade_ ));
    InMux I__1610 (
            .O(N__7952),
            .I(N__7949));
    LocalMux I__1609 (
            .O(N__7949),
            .I(N__7943));
    InMux I__1608 (
            .O(N__7948),
            .I(N__7938));
    InMux I__1607 (
            .O(N__7947),
            .I(N__7938));
    InMux I__1606 (
            .O(N__7946),
            .I(N__7935));
    Odrv12 I__1605 (
            .O(N__7943),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_5 ));
    LocalMux I__1604 (
            .O(N__7938),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_5 ));
    LocalMux I__1603 (
            .O(N__7935),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_5 ));
    InMux I__1602 (
            .O(N__7928),
            .I(N__7925));
    LocalMux I__1601 (
            .O(N__7925),
            .I(N__7922));
    Odrv12 I__1600 (
            .O(N__7922),
            .I(\U409_ADDRESS_DECODE.AUTOVECTOR_4Z0Z_0 ));
    InMux I__1599 (
            .O(N__7919),
            .I(N__7916));
    LocalMux I__1598 (
            .O(N__7916),
            .I(N__7913));
    Span4Mux_v I__1597 (
            .O(N__7913),
            .I(N__7910));
    Span4Mux_v I__1596 (
            .O(N__7910),
            .I(N__7907));
    Sp12to4 I__1595 (
            .O(N__7907),
            .I(N__7904));
    Odrv12 I__1594 (
            .O(N__7904),
            .I(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8 ));
    InMux I__1593 (
            .O(N__7901),
            .I(N__7898));
    LocalMux I__1592 (
            .O(N__7898),
            .I(U409_ADDRESS_DECODE_AUTOVECTOR_11));
    InMux I__1591 (
            .O(N__7895),
            .I(N__7892));
    LocalMux I__1590 (
            .O(N__7892),
            .I(\U409_CIA.CLK_CIA6_4 ));
    CascadeMux I__1589 (
            .O(N__7889),
            .I(\U409_CIA.un1_CIA_CLK_COUNT_3_2_cascade_ ));
    InMux I__1588 (
            .O(N__7886),
            .I(N__7883));
    LocalMux I__1587 (
            .O(N__7883),
            .I(N__7880));
    Span4Mux_v I__1586 (
            .O(N__7880),
            .I(N__7877));
    Span4Mux_h I__1585 (
            .O(N__7877),
            .I(N__7873));
    InMux I__1584 (
            .O(N__7876),
            .I(N__7870));
    Odrv4 I__1583 (
            .O(N__7873),
            .I(CIA_SPACE));
    LocalMux I__1582 (
            .O(N__7870),
            .I(CIA_SPACE));
    CascadeMux I__1581 (
            .O(N__7865),
            .I(\U409_CIA.VMA_RNOZ0Z_0_cascade_ ));
    InMux I__1580 (
            .O(N__7862),
            .I(N__7853));
    InMux I__1579 (
            .O(N__7861),
            .I(N__7853));
    InMux I__1578 (
            .O(N__7860),
            .I(N__7853));
    LocalMux I__1577 (
            .O(N__7853),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ));
    CascadeMux I__1576 (
            .O(N__7850),
            .I(N__7844));
    InMux I__1575 (
            .O(N__7849),
            .I(N__7840));
    InMux I__1574 (
            .O(N__7848),
            .I(N__7833));
    InMux I__1573 (
            .O(N__7847),
            .I(N__7833));
    InMux I__1572 (
            .O(N__7844),
            .I(N__7833));
    InMux I__1571 (
            .O(N__7843),
            .I(N__7830));
    LocalMux I__1570 (
            .O(N__7840),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__1569 (
            .O(N__7833),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__1568 (
            .O(N__7830),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    CascadeMux I__1567 (
            .O(N__7823),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_ ));
    InMux I__1566 (
            .O(N__7820),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ));
    InMux I__1565 (
            .O(N__7817),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ));
    InMux I__1564 (
            .O(N__7814),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ));
    InMux I__1563 (
            .O(N__7811),
            .I(N__7808));
    LocalMux I__1562 (
            .O(N__7808),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO ));
    InMux I__1561 (
            .O(N__7805),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ));
    InMux I__1560 (
            .O(N__7802),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ));
    InMux I__1559 (
            .O(N__7799),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ));
    InMux I__1558 (
            .O(N__7796),
            .I(N__7793));
    LocalMux I__1557 (
            .O(N__7793),
            .I(\U409_CIA.CIA_CLK_COUNT11_2_0 ));
    CascadeMux I__1556 (
            .O(N__7790),
            .I(N__7787));
    InMux I__1555 (
            .O(N__7787),
            .I(N__7783));
    InMux I__1554 (
            .O(N__7786),
            .I(N__7780));
    LocalMux I__1553 (
            .O(N__7783),
            .I(\U409_CIA.CIA_CLK_COUNT11_3 ));
    LocalMux I__1552 (
            .O(N__7780),
            .I(\U409_CIA.CIA_CLK_COUNT11_3 ));
    InMux I__1551 (
            .O(N__7775),
            .I(N__7772));
    LocalMux I__1550 (
            .O(N__7772),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ));
    CascadeMux I__1549 (
            .O(N__7769),
            .I(N__7766));
    InMux I__1548 (
            .O(N__7766),
            .I(N__7763));
    LocalMux I__1547 (
            .O(N__7763),
            .I(\U409_TRANSFER_ACK.TACK_EN8 ));
    InMux I__1546 (
            .O(N__7760),
            .I(N__7757));
    LocalMux I__1545 (
            .O(N__7757),
            .I(\U409_TRANSFER_ACK.TACK_STATE_ns_1_0 ));
    InMux I__1544 (
            .O(N__7754),
            .I(N__7748));
    InMux I__1543 (
            .O(N__7753),
            .I(N__7743));
    InMux I__1542 (
            .O(N__7752),
            .I(N__7743));
    InMux I__1541 (
            .O(N__7751),
            .I(N__7740));
    LocalMux I__1540 (
            .O(N__7748),
            .I(\U409_TRANSFER_ACK.TACK_STATEZ0Z_0 ));
    LocalMux I__1539 (
            .O(N__7743),
            .I(\U409_TRANSFER_ACK.TACK_STATEZ0Z_0 ));
    LocalMux I__1538 (
            .O(N__7740),
            .I(\U409_TRANSFER_ACK.TACK_STATEZ0Z_0 ));
    CascadeMux I__1537 (
            .O(N__7733),
            .I(N__7728));
    InMux I__1536 (
            .O(N__7732),
            .I(N__7721));
    InMux I__1535 (
            .O(N__7731),
            .I(N__7721));
    InMux I__1534 (
            .O(N__7728),
            .I(N__7721));
    LocalMux I__1533 (
            .O(N__7721),
            .I(\U409_TRANSFER_ACK.TACK_STATEZ0Z_1 ));
    InMux I__1532 (
            .O(N__7718),
            .I(N__7714));
    InMux I__1531 (
            .O(N__7717),
            .I(N__7711));
    LocalMux I__1530 (
            .O(N__7714),
            .I(N__7705));
    LocalMux I__1529 (
            .O(N__7711),
            .I(N__7705));
    InMux I__1528 (
            .O(N__7710),
            .I(N__7700));
    Span4Mux_v I__1527 (
            .O(N__7705),
            .I(N__7697));
    InMux I__1526 (
            .O(N__7704),
            .I(N__7694));
    InMux I__1525 (
            .O(N__7703),
            .I(N__7691));
    LocalMux I__1524 (
            .O(N__7700),
            .I(N__7687));
    Span4Mux_h I__1523 (
            .O(N__7697),
            .I(N__7680));
    LocalMux I__1522 (
            .O(N__7694),
            .I(N__7680));
    LocalMux I__1521 (
            .O(N__7691),
            .I(N__7680));
    InMux I__1520 (
            .O(N__7690),
            .I(N__7677));
    Span4Mux_v I__1519 (
            .O(N__7687),
            .I(N__7674));
    Span4Mux_h I__1518 (
            .O(N__7680),
            .I(N__7671));
    LocalMux I__1517 (
            .O(N__7677),
            .I(N__7668));
    Span4Mux_v I__1516 (
            .O(N__7674),
            .I(N__7665));
    Span4Mux_v I__1515 (
            .O(N__7671),
            .I(N__7662));
    Span12Mux_h I__1514 (
            .O(N__7668),
            .I(N__7659));
    Span4Mux_v I__1513 (
            .O(N__7665),
            .I(N__7656));
    Span4Mux_v I__1512 (
            .O(N__7662),
            .I(N__7653));
    Odrv12 I__1511 (
            .O(N__7659),
            .I(U409_ADDRESS_DECODE_Z2_SPACE));
    Odrv4 I__1510 (
            .O(N__7656),
            .I(U409_ADDRESS_DECODE_Z2_SPACE));
    Odrv4 I__1509 (
            .O(N__7653),
            .I(U409_ADDRESS_DECODE_Z2_SPACE));
    CascadeMux I__1508 (
            .O(N__7646),
            .I(N__7642));
    InMux I__1507 (
            .O(N__7645),
            .I(N__7639));
    InMux I__1506 (
            .O(N__7642),
            .I(N__7636));
    LocalMux I__1505 (
            .O(N__7639),
            .I(N__7631));
    LocalMux I__1504 (
            .O(N__7636),
            .I(N__7631));
    Span4Mux_v I__1503 (
            .O(N__7631),
            .I(N__7628));
    Span4Mux_h I__1502 (
            .O(N__7628),
            .I(N__7625));
    Odrv4 I__1501 (
            .O(N__7625),
            .I(U409_ADDRESS_DECODE_HIROM));
    IoInMux I__1500 (
            .O(N__7622),
            .I(N__7619));
    LocalMux I__1499 (
            .O(N__7619),
            .I(N__7616));
    IoSpan4Mux I__1498 (
            .O(N__7616),
            .I(N__7612));
    IoInMux I__1497 (
            .O(N__7615),
            .I(N__7609));
    Span4Mux_s2_v I__1496 (
            .O(N__7612),
            .I(N__7606));
    LocalMux I__1495 (
            .O(N__7609),
            .I(N__7602));
    Span4Mux_v I__1494 (
            .O(N__7606),
            .I(N__7599));
    CascadeMux I__1493 (
            .O(N__7605),
            .I(N__7596));
    Span12Mux_s8_v I__1492 (
            .O(N__7602),
            .I(N__7593));
    Sp12to4 I__1491 (
            .O(N__7599),
            .I(N__7590));
    InMux I__1490 (
            .O(N__7596),
            .I(N__7587));
    Span12Mux_h I__1489 (
            .O(N__7593),
            .I(N__7583));
    Span12Mux_v I__1488 (
            .O(N__7590),
            .I(N__7580));
    LocalMux I__1487 (
            .O(N__7587),
            .I(N__7577));
    InMux I__1486 (
            .O(N__7586),
            .I(N__7574));
    Odrv12 I__1485 (
            .O(N__7583),
            .I(TACK_OUT));
    Odrv12 I__1484 (
            .O(N__7580),
            .I(TACK_OUT));
    Odrv4 I__1483 (
            .O(N__7577),
            .I(TACK_OUT));
    LocalMux I__1482 (
            .O(N__7574),
            .I(TACK_OUT));
    InMux I__1481 (
            .O(N__7565),
            .I(N__7562));
    LocalMux I__1480 (
            .O(N__7562),
            .I(N__7558));
    InMux I__1479 (
            .O(N__7561),
            .I(N__7555));
    Span4Mux_h I__1478 (
            .O(N__7558),
            .I(N__7552));
    LocalMux I__1477 (
            .O(N__7555),
            .I(N__7549));
    Odrv4 I__1476 (
            .O(N__7552),
            .I(U409_ADDRESS_DECODE_LOWROM));
    Odrv12 I__1475 (
            .O(N__7549),
            .I(U409_ADDRESS_DECODE_LOWROM));
    IoInMux I__1474 (
            .O(N__7544),
            .I(N__7541));
    LocalMux I__1473 (
            .O(N__7541),
            .I(N__7538));
    Span4Mux_s2_v I__1472 (
            .O(N__7538),
            .I(N__7535));
    Sp12to4 I__1471 (
            .O(N__7535),
            .I(N__7532));
    Span12Mux_h I__1470 (
            .O(N__7532),
            .I(N__7529));
    Span12Mux_v I__1469 (
            .O(N__7529),
            .I(N__7526));
    Odrv12 I__1468 (
            .O(N__7526),
            .I(U409_TRANSFER_ACK_un1_TACK_OUT_0_i));
    IoInMux I__1467 (
            .O(N__7523),
            .I(N__7520));
    LocalMux I__1466 (
            .O(N__7520),
            .I(N__7517));
    Span4Mux_s2_v I__1465 (
            .O(N__7517),
            .I(N__7514));
    Span4Mux_v I__1464 (
            .O(N__7514),
            .I(N__7511));
    Odrv4 I__1463 (
            .O(N__7511),
            .I(GB_BUFFER_CLK40_IN_c_g_THRU_CO));
    CascadeMux I__1462 (
            .O(N__7508),
            .I(\U409_CIA.CIA_CLK_COUNT11_2_0_cascade_ ));
    CascadeMux I__1461 (
            .O(N__7505),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_ ));
    CascadeMux I__1460 (
            .O(N__7502),
            .I(N__7499));
    InMux I__1459 (
            .O(N__7499),
            .I(N__7496));
    LocalMux I__1458 (
            .O(N__7496),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ));
    CascadeMux I__1457 (
            .O(N__7493),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ));
    CascadeMux I__1456 (
            .O(N__7490),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ));
    InMux I__1455 (
            .O(N__7487),
            .I(N__7481));
    InMux I__1454 (
            .O(N__7486),
            .I(N__7481));
    LocalMux I__1453 (
            .O(N__7481),
            .I(N__7478));
    Span4Mux_v I__1452 (
            .O(N__7478),
            .I(N__7474));
    InMux I__1451 (
            .O(N__7477),
            .I(N__7471));
    Odrv4 I__1450 (
            .O(N__7474),
            .I(\U409_AUTOCONFIG.N_78 ));
    LocalMux I__1449 (
            .O(N__7471),
            .I(\U409_AUTOCONFIG.N_78 ));
    InMux I__1448 (
            .O(N__7466),
            .I(N__7460));
    InMux I__1447 (
            .O(N__7465),
            .I(N__7460));
    LocalMux I__1446 (
            .O(N__7460),
            .I(N__7457));
    Odrv12 I__1445 (
            .O(N__7457),
            .I(\U409_AUTOCONFIG.N_92 ));
    InMux I__1444 (
            .O(N__7454),
            .I(N__7451));
    LocalMux I__1443 (
            .O(N__7451),
            .I(N__7448));
    Odrv4 I__1442 (
            .O(N__7448),
            .I(\U409_AUTOCONFIG.PR_OUTZ0Z_0 ));
    InMux I__1441 (
            .O(N__7445),
            .I(N__7442));
    LocalMux I__1440 (
            .O(N__7442),
            .I(N__7439));
    Odrv12 I__1439 (
            .O(N__7439),
            .I(\U409_AUTOCONFIG.LIDE_OUT_7_i_a3_1_0 ));
    CascadeMux I__1438 (
            .O(N__7436),
            .I(N__7433));
    InMux I__1437 (
            .O(N__7433),
            .I(N__7430));
    LocalMux I__1436 (
            .O(N__7430),
            .I(N__7427));
    Span12Mux_h I__1435 (
            .O(N__7427),
            .I(N__7424));
    Odrv12 I__1434 (
            .O(N__7424),
            .I(\U409_AUTOCONFIG.LIDE_OUT_7_i_a3_0_0 ));
    InMux I__1433 (
            .O(N__7421),
            .I(N__7418));
    LocalMux I__1432 (
            .O(N__7418),
            .I(N__7415));
    Odrv12 I__1431 (
            .O(N__7415),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_0 ));
    CEMux I__1430 (
            .O(N__7412),
            .I(N__7408));
    CEMux I__1429 (
            .O(N__7411),
            .I(N__7403));
    LocalMux I__1428 (
            .O(N__7408),
            .I(N__7400));
    CEMux I__1427 (
            .O(N__7407),
            .I(N__7397));
    CEMux I__1426 (
            .O(N__7406),
            .I(N__7394));
    LocalMux I__1425 (
            .O(N__7403),
            .I(N__7391));
    Span4Mux_v I__1424 (
            .O(N__7400),
            .I(N__7385));
    LocalMux I__1423 (
            .O(N__7397),
            .I(N__7385));
    LocalMux I__1422 (
            .O(N__7394),
            .I(N__7382));
    Span4Mux_v I__1421 (
            .O(N__7391),
            .I(N__7379));
    CEMux I__1420 (
            .O(N__7390),
            .I(N__7376));
    Span4Mux_v I__1419 (
            .O(N__7385),
            .I(N__7371));
    Span4Mux_v I__1418 (
            .O(N__7382),
            .I(N__7371));
    Span4Mux_h I__1417 (
            .O(N__7379),
            .I(N__7368));
    LocalMux I__1416 (
            .O(N__7376),
            .I(N__7365));
    Span4Mux_h I__1415 (
            .O(N__7371),
            .I(N__7362));
    Odrv4 I__1414 (
            .O(N__7368),
            .I(\U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i ));
    Odrv12 I__1413 (
            .O(N__7365),
            .I(\U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i ));
    Odrv4 I__1412 (
            .O(N__7362),
            .I(\U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i ));
    InMux I__1411 (
            .O(N__7355),
            .I(N__7352));
    LocalMux I__1410 (
            .O(N__7352),
            .I(N__7348));
    InMux I__1409 (
            .O(N__7351),
            .I(N__7345));
    Odrv4 I__1408 (
            .O(N__7348),
            .I(\U409_AUTOCONFIG.N_133 ));
    LocalMux I__1407 (
            .O(N__7345),
            .I(\U409_AUTOCONFIG.N_133 ));
    CascadeMux I__1406 (
            .O(N__7340),
            .I(N__7334));
    InMux I__1405 (
            .O(N__7339),
            .I(N__7329));
    InMux I__1404 (
            .O(N__7338),
            .I(N__7326));
    CascadeMux I__1403 (
            .O(N__7337),
            .I(N__7317));
    InMux I__1402 (
            .O(N__7334),
            .I(N__7308));
    InMux I__1401 (
            .O(N__7333),
            .I(N__7308));
    InMux I__1400 (
            .O(N__7332),
            .I(N__7305));
    LocalMux I__1399 (
            .O(N__7329),
            .I(N__7300));
    LocalMux I__1398 (
            .O(N__7326),
            .I(N__7300));
    InMux I__1397 (
            .O(N__7325),
            .I(N__7297));
    InMux I__1396 (
            .O(N__7324),
            .I(N__7294));
    InMux I__1395 (
            .O(N__7323),
            .I(N__7291));
    InMux I__1394 (
            .O(N__7322),
            .I(N__7288));
    InMux I__1393 (
            .O(N__7321),
            .I(N__7285));
    InMux I__1392 (
            .O(N__7320),
            .I(N__7282));
    InMux I__1391 (
            .O(N__7317),
            .I(N__7275));
    InMux I__1390 (
            .O(N__7316),
            .I(N__7275));
    InMux I__1389 (
            .O(N__7315),
            .I(N__7275));
    InMux I__1388 (
            .O(N__7314),
            .I(N__7272));
    InMux I__1387 (
            .O(N__7313),
            .I(N__7269));
    LocalMux I__1386 (
            .O(N__7308),
            .I(N__7266));
    LocalMux I__1385 (
            .O(N__7305),
            .I(N__7263));
    Span4Mux_v I__1384 (
            .O(N__7300),
            .I(N__7250));
    LocalMux I__1383 (
            .O(N__7297),
            .I(N__7250));
    LocalMux I__1382 (
            .O(N__7294),
            .I(N__7250));
    LocalMux I__1381 (
            .O(N__7291),
            .I(N__7250));
    LocalMux I__1380 (
            .O(N__7288),
            .I(N__7250));
    LocalMux I__1379 (
            .O(N__7285),
            .I(N__7250));
    LocalMux I__1378 (
            .O(N__7282),
            .I(N__7247));
    LocalMux I__1377 (
            .O(N__7275),
            .I(N__7240));
    LocalMux I__1376 (
            .O(N__7272),
            .I(N__7240));
    LocalMux I__1375 (
            .O(N__7269),
            .I(N__7240));
    Span4Mux_v I__1374 (
            .O(N__7266),
            .I(N__7235));
    Span4Mux_v I__1373 (
            .O(N__7263),
            .I(N__7235));
    Span4Mux_v I__1372 (
            .O(N__7250),
            .I(N__7232));
    Span4Mux_v I__1371 (
            .O(N__7247),
            .I(N__7227));
    Span4Mux_v I__1370 (
            .O(N__7240),
            .I(N__7227));
    Sp12to4 I__1369 (
            .O(N__7235),
            .I(N__7220));
    Sp12to4 I__1368 (
            .O(N__7232),
            .I(N__7220));
    Sp12to4 I__1367 (
            .O(N__7227),
            .I(N__7220));
    Span12Mux_h I__1366 (
            .O(N__7220),
            .I(N__7217));
    Span12Mux_v I__1365 (
            .O(N__7217),
            .I(N__7214));
    Odrv12 I__1364 (
            .O(N__7214),
            .I(A_c_1));
    CascadeMux I__1363 (
            .O(N__7211),
            .I(N__7208));
    InMux I__1362 (
            .O(N__7208),
            .I(N__7205));
    LocalMux I__1361 (
            .O(N__7205),
            .I(N__7202));
    Span4Mux_v I__1360 (
            .O(N__7202),
            .I(N__7199));
    Span4Mux_h I__1359 (
            .O(N__7199),
            .I(N__7196));
    Sp12to4 I__1358 (
            .O(N__7196),
            .I(N__7193));
    Span12Mux_h I__1357 (
            .O(N__7193),
            .I(N__7190));
    Span12Mux_v I__1356 (
            .O(N__7190),
            .I(N__7187));
    Odrv12 I__1355 (
            .O(N__7187),
            .I(AUTOBOOT_c));
    CascadeMux I__1354 (
            .O(N__7184),
            .I(N__7180));
    InMux I__1353 (
            .O(N__7183),
            .I(N__7175));
    InMux I__1352 (
            .O(N__7180),
            .I(N__7175));
    LocalMux I__1351 (
            .O(N__7175),
            .I(N__7171));
    InMux I__1350 (
            .O(N__7174),
            .I(N__7168));
    Odrv4 I__1349 (
            .O(N__7171),
            .I(\U409_AUTOCONFIG.N_126 ));
    LocalMux I__1348 (
            .O(N__7168),
            .I(\U409_AUTOCONFIG.N_126 ));
    InMux I__1347 (
            .O(N__7163),
            .I(N__7160));
    LocalMux I__1346 (
            .O(N__7160),
            .I(\U409_AUTOCONFIG.LIDE_OUT_7_i_1_0 ));
    InMux I__1345 (
            .O(N__7157),
            .I(N__7154));
    LocalMux I__1344 (
            .O(N__7154),
            .I(N__7151));
    Span12Mux_h I__1343 (
            .O(N__7151),
            .I(N__7148));
    Span12Mux_v I__1342 (
            .O(N__7148),
            .I(N__7145));
    Odrv12 I__1341 (
            .O(N__7145),
            .I(TACKn_in));
    InMux I__1340 (
            .O(N__7142),
            .I(N__7139));
    LocalMux I__1339 (
            .O(N__7139),
            .I(N__7134));
    InMux I__1338 (
            .O(N__7138),
            .I(N__7129));
    InMux I__1337 (
            .O(N__7137),
            .I(N__7129));
    Odrv12 I__1336 (
            .O(N__7134),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn));
    LocalMux I__1335 (
            .O(N__7129),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn));
    CascadeMux I__1334 (
            .O(N__7124),
            .I(N__7121));
    InMux I__1333 (
            .O(N__7121),
            .I(N__7118));
    LocalMux I__1332 (
            .O(N__7118),
            .I(N__7114));
    InMux I__1331 (
            .O(N__7117),
            .I(N__7111));
    Span4Mux_v I__1330 (
            .O(N__7114),
            .I(N__7108));
    LocalMux I__1329 (
            .O(N__7111),
            .I(N__7105));
    Odrv4 I__1328 (
            .O(N__7108),
            .I(U409_ADDRESS_DECODE_un1_RAMSPACEn));
    Odrv4 I__1327 (
            .O(N__7105),
            .I(U409_ADDRESS_DECODE_un1_RAMSPACEn));
    InMux I__1326 (
            .O(N__7100),
            .I(N__7096));
    InMux I__1325 (
            .O(N__7099),
            .I(N__7090));
    LocalMux I__1324 (
            .O(N__7096),
            .I(N__7085));
    InMux I__1323 (
            .O(N__7095),
            .I(N__7082));
    InMux I__1322 (
            .O(N__7094),
            .I(N__7077));
    InMux I__1321 (
            .O(N__7093),
            .I(N__7077));
    LocalMux I__1320 (
            .O(N__7090),
            .I(N__7074));
    InMux I__1319 (
            .O(N__7089),
            .I(N__7069));
    InMux I__1318 (
            .O(N__7088),
            .I(N__7069));
    Span4Mux_h I__1317 (
            .O(N__7085),
            .I(N__7064));
    LocalMux I__1316 (
            .O(N__7082),
            .I(N__7064));
    LocalMux I__1315 (
            .O(N__7077),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    Odrv4 I__1314 (
            .O(N__7074),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    LocalMux I__1313 (
            .O(N__7069),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    Odrv4 I__1312 (
            .O(N__7064),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    CEMux I__1311 (
            .O(N__7055),
            .I(N__7052));
    LocalMux I__1310 (
            .O(N__7052),
            .I(N__7049));
    Odrv4 I__1309 (
            .O(N__7049),
            .I(\U409_AUTOCONFIG.STATE_ns_0_0_1 ));
    CascadeMux I__1308 (
            .O(N__7046),
            .I(N__7041));
    InMux I__1307 (
            .O(N__7045),
            .I(N__7037));
    InMux I__1306 (
            .O(N__7044),
            .I(N__7032));
    InMux I__1305 (
            .O(N__7041),
            .I(N__7032));
    InMux I__1304 (
            .O(N__7040),
            .I(N__7029));
    LocalMux I__1303 (
            .O(N__7037),
            .I(\U409_AUTOCONFIG.N_4 ));
    LocalMux I__1302 (
            .O(N__7032),
            .I(\U409_AUTOCONFIG.N_4 ));
    LocalMux I__1301 (
            .O(N__7029),
            .I(\U409_AUTOCONFIG.N_4 ));
    IoInMux I__1300 (
            .O(N__7022),
            .I(N__7019));
    LocalMux I__1299 (
            .O(N__7019),
            .I(N__7016));
    IoSpan4Mux I__1298 (
            .O(N__7016),
            .I(N__7013));
    Sp12to4 I__1297 (
            .O(N__7013),
            .I(N__7010));
    Span12Mux_s9_v I__1296 (
            .O(N__7010),
            .I(N__7007));
    Odrv12 I__1295 (
            .O(N__7007),
            .I(D_OUT_0));
    InMux I__1294 (
            .O(N__7004),
            .I(N__7001));
    LocalMux I__1293 (
            .O(N__7001),
            .I(N__6998));
    Odrv4 I__1292 (
            .O(N__6998),
            .I(\U409_AUTOCONFIG.LIDE_OUT_RNI7DMPZ0Z_1 ));
    InMux I__1291 (
            .O(N__6995),
            .I(N__6991));
    InMux I__1290 (
            .O(N__6994),
            .I(N__6988));
    LocalMux I__1289 (
            .O(N__6991),
            .I(N__6976));
    LocalMux I__1288 (
            .O(N__6988),
            .I(N__6976));
    InMux I__1287 (
            .O(N__6987),
            .I(N__6971));
    InMux I__1286 (
            .O(N__6986),
            .I(N__6971));
    InMux I__1285 (
            .O(N__6985),
            .I(N__6966));
    InMux I__1284 (
            .O(N__6984),
            .I(N__6966));
    InMux I__1283 (
            .O(N__6983),
            .I(N__6963));
    InMux I__1282 (
            .O(N__6982),
            .I(N__6958));
    InMux I__1281 (
            .O(N__6981),
            .I(N__6958));
    Odrv4 I__1280 (
            .O(N__6976),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    LocalMux I__1279 (
            .O(N__6971),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    LocalMux I__1278 (
            .O(N__6966),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    LocalMux I__1277 (
            .O(N__6963),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    LocalMux I__1276 (
            .O(N__6958),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    InMux I__1275 (
            .O(N__6947),
            .I(N__6944));
    LocalMux I__1274 (
            .O(N__6944),
            .I(\U409_AUTOCONFIG.LIDE_OUT_RNI5BMPZ0Z_0 ));
    CascadeMux I__1273 (
            .O(N__6941),
            .I(N__6932));
    CascadeMux I__1272 (
            .O(N__6940),
            .I(N__6929));
    CascadeMux I__1271 (
            .O(N__6939),
            .I(N__6925));
    InMux I__1270 (
            .O(N__6938),
            .I(N__6921));
    InMux I__1269 (
            .O(N__6937),
            .I(N__6916));
    InMux I__1268 (
            .O(N__6936),
            .I(N__6916));
    CascadeMux I__1267 (
            .O(N__6935),
            .I(N__6913));
    InMux I__1266 (
            .O(N__6932),
            .I(N__6906));
    InMux I__1265 (
            .O(N__6929),
            .I(N__6906));
    InMux I__1264 (
            .O(N__6928),
            .I(N__6906));
    InMux I__1263 (
            .O(N__6925),
            .I(N__6903));
    CascadeMux I__1262 (
            .O(N__6924),
            .I(N__6899));
    LocalMux I__1261 (
            .O(N__6921),
            .I(N__6896));
    LocalMux I__1260 (
            .O(N__6916),
            .I(N__6893));
    InMux I__1259 (
            .O(N__6913),
            .I(N__6890));
    LocalMux I__1258 (
            .O(N__6906),
            .I(N__6885));
    LocalMux I__1257 (
            .O(N__6903),
            .I(N__6885));
    InMux I__1256 (
            .O(N__6902),
            .I(N__6880));
    InMux I__1255 (
            .O(N__6899),
            .I(N__6880));
    Span4Mux_v I__1254 (
            .O(N__6896),
            .I(N__6876));
    Span4Mux_v I__1253 (
            .O(N__6893),
            .I(N__6871));
    LocalMux I__1252 (
            .O(N__6890),
            .I(N__6871));
    Span4Mux_h I__1251 (
            .O(N__6885),
            .I(N__6866));
    LocalMux I__1250 (
            .O(N__6880),
            .I(N__6866));
    InMux I__1249 (
            .O(N__6879),
            .I(N__6863));
    Odrv4 I__1248 (
            .O(N__6876),
            .I(AUTOCONFIG_SPACE));
    Odrv4 I__1247 (
            .O(N__6871),
            .I(AUTOCONFIG_SPACE));
    Odrv4 I__1246 (
            .O(N__6866),
            .I(AUTOCONFIG_SPACE));
    LocalMux I__1245 (
            .O(N__6863),
            .I(AUTOCONFIG_SPACE));
    CascadeMux I__1244 (
            .O(N__6854),
            .I(N__6849));
    InMux I__1243 (
            .O(N__6853),
            .I(N__6843));
    InMux I__1242 (
            .O(N__6852),
            .I(N__6839));
    InMux I__1241 (
            .O(N__6849),
            .I(N__6836));
    InMux I__1240 (
            .O(N__6848),
            .I(N__6831));
    InMux I__1239 (
            .O(N__6847),
            .I(N__6831));
    InMux I__1238 (
            .O(N__6846),
            .I(N__6828));
    LocalMux I__1237 (
            .O(N__6843),
            .I(N__6825));
    InMux I__1236 (
            .O(N__6842),
            .I(N__6822));
    LocalMux I__1235 (
            .O(N__6839),
            .I(CONFIGURED));
    LocalMux I__1234 (
            .O(N__6836),
            .I(CONFIGURED));
    LocalMux I__1233 (
            .O(N__6831),
            .I(CONFIGURED));
    LocalMux I__1232 (
            .O(N__6828),
            .I(CONFIGURED));
    Odrv4 I__1231 (
            .O(N__6825),
            .I(CONFIGURED));
    LocalMux I__1230 (
            .O(N__6822),
            .I(CONFIGURED));
    InMux I__1229 (
            .O(N__6809),
            .I(N__6805));
    InMux I__1228 (
            .O(N__6808),
            .I(N__6802));
    LocalMux I__1227 (
            .O(N__6805),
            .I(\U409_AUTOCONFIG.AC_STARTZ0 ));
    LocalMux I__1226 (
            .O(N__6802),
            .I(\U409_AUTOCONFIG.AC_STARTZ0 ));
    InMux I__1225 (
            .O(N__6797),
            .I(N__6794));
    LocalMux I__1224 (
            .O(N__6794),
            .I(N__6791));
    Odrv4 I__1223 (
            .O(N__6791),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0 ));
    InMux I__1222 (
            .O(N__6788),
            .I(N__6785));
    LocalMux I__1221 (
            .O(N__6785),
            .I(\U409_AUTOCONFIG.N_82 ));
    InMux I__1220 (
            .O(N__6782),
            .I(N__6779));
    LocalMux I__1219 (
            .O(N__6779),
            .I(N__6776));
    Odrv4 I__1218 (
            .O(N__6776),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ));
    CascadeMux I__1217 (
            .O(N__6773),
            .I(N__6770));
    InMux I__1216 (
            .O(N__6770),
            .I(N__6767));
    LocalMux I__1215 (
            .O(N__6767),
            .I(N__6764));
    Odrv4 I__1214 (
            .O(N__6764),
            .I(\U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_0Z0Z_3 ));
    InMux I__1213 (
            .O(N__6761),
            .I(N__6758));
    LocalMux I__1212 (
            .O(N__6758),
            .I(N__6755));
    Odrv12 I__1211 (
            .O(N__6755),
            .I(\U409_AUTOCONFIG.PR_OUTZ0Z_3 ));
    CascadeMux I__1210 (
            .O(N__6752),
            .I(N__6748));
    InMux I__1209 (
            .O(N__6751),
            .I(N__6743));
    InMux I__1208 (
            .O(N__6748),
            .I(N__6743));
    LocalMux I__1207 (
            .O(N__6743),
            .I(N__6740));
    Odrv4 I__1206 (
            .O(N__6740),
            .I(\U409_AUTOCONFIG.N_131 ));
    InMux I__1205 (
            .O(N__6737),
            .I(N__6734));
    LocalMux I__1204 (
            .O(N__6734),
            .I(\U409_AUTOCONFIG.N_93 ));
    CascadeMux I__1203 (
            .O(N__6731),
            .I(N__6728));
    InMux I__1202 (
            .O(N__6728),
            .I(N__6725));
    LocalMux I__1201 (
            .O(N__6725),
            .I(N__6722));
    Odrv12 I__1200 (
            .O(N__6722),
            .I(\U409_AUTOCONFIG.PR_OUTZ0Z_1 ));
    InMux I__1199 (
            .O(N__6719),
            .I(N__6713));
    InMux I__1198 (
            .O(N__6718),
            .I(N__6713));
    LocalMux I__1197 (
            .O(N__6713),
            .I(N__6709));
    InMux I__1196 (
            .O(N__6712),
            .I(N__6706));
    Span4Mux_v I__1195 (
            .O(N__6709),
            .I(N__6701));
    LocalMux I__1194 (
            .O(N__6706),
            .I(N__6698));
    InMux I__1193 (
            .O(N__6705),
            .I(N__6693));
    InMux I__1192 (
            .O(N__6704),
            .I(N__6693));
    Odrv4 I__1191 (
            .O(N__6701),
            .I(\U409_AUTOCONFIG.N_116 ));
    Odrv4 I__1190 (
            .O(N__6698),
            .I(\U409_AUTOCONFIG.N_116 ));
    LocalMux I__1189 (
            .O(N__6693),
            .I(\U409_AUTOCONFIG.N_116 ));
    InMux I__1188 (
            .O(N__6686),
            .I(N__6679));
    InMux I__1187 (
            .O(N__6685),
            .I(N__6679));
    InMux I__1186 (
            .O(N__6684),
            .I(N__6676));
    LocalMux I__1185 (
            .O(N__6679),
            .I(N__6665));
    LocalMux I__1184 (
            .O(N__6676),
            .I(N__6665));
    InMux I__1183 (
            .O(N__6675),
            .I(N__6660));
    InMux I__1182 (
            .O(N__6674),
            .I(N__6660));
    CascadeMux I__1181 (
            .O(N__6673),
            .I(N__6657));
    InMux I__1180 (
            .O(N__6672),
            .I(N__6652));
    InMux I__1179 (
            .O(N__6671),
            .I(N__6649));
    InMux I__1178 (
            .O(N__6670),
            .I(N__6646));
    Span4Mux_v I__1177 (
            .O(N__6665),
            .I(N__6641));
    LocalMux I__1176 (
            .O(N__6660),
            .I(N__6641));
    InMux I__1175 (
            .O(N__6657),
            .I(N__6636));
    InMux I__1174 (
            .O(N__6656),
            .I(N__6636));
    InMux I__1173 (
            .O(N__6655),
            .I(N__6633));
    LocalMux I__1172 (
            .O(N__6652),
            .I(N__6627));
    LocalMux I__1171 (
            .O(N__6649),
            .I(N__6627));
    LocalMux I__1170 (
            .O(N__6646),
            .I(N__6620));
    Span4Mux_v I__1169 (
            .O(N__6641),
            .I(N__6620));
    LocalMux I__1168 (
            .O(N__6636),
            .I(N__6620));
    LocalMux I__1167 (
            .O(N__6633),
            .I(N__6617));
    InMux I__1166 (
            .O(N__6632),
            .I(N__6614));
    Span4Mux_v I__1165 (
            .O(N__6627),
            .I(N__6611));
    Span4Mux_h I__1164 (
            .O(N__6620),
            .I(N__6604));
    Span4Mux_v I__1163 (
            .O(N__6617),
            .I(N__6604));
    LocalMux I__1162 (
            .O(N__6614),
            .I(N__6604));
    Span4Mux_v I__1161 (
            .O(N__6611),
            .I(N__6601));
    Span4Mux_v I__1160 (
            .O(N__6604),
            .I(N__6598));
    Sp12to4 I__1159 (
            .O(N__6601),
            .I(N__6593));
    Sp12to4 I__1158 (
            .O(N__6598),
            .I(N__6593));
    Span12Mux_h I__1157 (
            .O(N__6593),
            .I(N__6590));
    Odrv12 I__1156 (
            .O(N__6590),
            .I(A_c_2));
    InMux I__1155 (
            .O(N__6587),
            .I(N__6584));
    LocalMux I__1154 (
            .O(N__6584),
            .I(N__6581));
    Odrv4 I__1153 (
            .O(N__6581),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1 ));
    InMux I__1152 (
            .O(N__6578),
            .I(N__6575));
    LocalMux I__1151 (
            .O(N__6575),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2 ));
    InMux I__1150 (
            .O(N__6572),
            .I(N__6569));
    LocalMux I__1149 (
            .O(N__6569),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ));
    InMux I__1148 (
            .O(N__6566),
            .I(N__6563));
    LocalMux I__1147 (
            .O(N__6563),
            .I(N__6560));
    Odrv12 I__1146 (
            .O(N__6560),
            .I(\U409_AUTOCONFIG.LIDE_OUT_RNI9FMPZ0Z_2 ));
    InMux I__1145 (
            .O(N__6557),
            .I(N__6554));
    LocalMux I__1144 (
            .O(N__6554),
            .I(N__6550));
    CascadeMux I__1143 (
            .O(N__6553),
            .I(N__6547));
    Span4Mux_v I__1142 (
            .O(N__6550),
            .I(N__6544));
    InMux I__1141 (
            .O(N__6547),
            .I(N__6541));
    Odrv4 I__1140 (
            .O(N__6544),
            .I(\U409_AUTOCONFIG.N_129 ));
    LocalMux I__1139 (
            .O(N__6541),
            .I(\U409_AUTOCONFIG.N_129 ));
    CascadeMux I__1138 (
            .O(N__6536),
            .I(\U409_AUTOCONFIG.N_133_cascade_ ));
    InMux I__1137 (
            .O(N__6533),
            .I(N__6527));
    InMux I__1136 (
            .O(N__6532),
            .I(N__6527));
    LocalMux I__1135 (
            .O(N__6527),
            .I(\U409_AUTOCONFIG.N_127 ));
    CascadeMux I__1134 (
            .O(N__6524),
            .I(N__6521));
    InMux I__1133 (
            .O(N__6521),
            .I(N__6515));
    InMux I__1132 (
            .O(N__6520),
            .I(N__6515));
    LocalMux I__1131 (
            .O(N__6515),
            .I(N__6508));
    InMux I__1130 (
            .O(N__6514),
            .I(N__6505));
    InMux I__1129 (
            .O(N__6513),
            .I(N__6502));
    InMux I__1128 (
            .O(N__6512),
            .I(N__6497));
    InMux I__1127 (
            .O(N__6511),
            .I(N__6497));
    Span4Mux_v I__1126 (
            .O(N__6508),
            .I(N__6492));
    LocalMux I__1125 (
            .O(N__6505),
            .I(N__6489));
    LocalMux I__1124 (
            .O(N__6502),
            .I(N__6486));
    LocalMux I__1123 (
            .O(N__6497),
            .I(N__6483));
    InMux I__1122 (
            .O(N__6496),
            .I(N__6480));
    InMux I__1121 (
            .O(N__6495),
            .I(N__6477));
    Odrv4 I__1120 (
            .O(N__6492),
            .I(\U409_AUTOCONFIG.N_110 ));
    Odrv4 I__1119 (
            .O(N__6489),
            .I(\U409_AUTOCONFIG.N_110 ));
    Odrv12 I__1118 (
            .O(N__6486),
            .I(\U409_AUTOCONFIG.N_110 ));
    Odrv12 I__1117 (
            .O(N__6483),
            .I(\U409_AUTOCONFIG.N_110 ));
    LocalMux I__1116 (
            .O(N__6480),
            .I(\U409_AUTOCONFIG.N_110 ));
    LocalMux I__1115 (
            .O(N__6477),
            .I(\U409_AUTOCONFIG.N_110 ));
    CascadeMux I__1114 (
            .O(N__6464),
            .I(N__6458));
    CascadeMux I__1113 (
            .O(N__6463),
            .I(N__6452));
    CascadeMux I__1112 (
            .O(N__6462),
            .I(N__6446));
    CascadeMux I__1111 (
            .O(N__6461),
            .I(N__6442));
    InMux I__1110 (
            .O(N__6458),
            .I(N__6439));
    InMux I__1109 (
            .O(N__6457),
            .I(N__6436));
    InMux I__1108 (
            .O(N__6456),
            .I(N__6433));
    InMux I__1107 (
            .O(N__6455),
            .I(N__6428));
    InMux I__1106 (
            .O(N__6452),
            .I(N__6428));
    CascadeMux I__1105 (
            .O(N__6451),
            .I(N__6425));
    CascadeMux I__1104 (
            .O(N__6450),
            .I(N__6422));
    InMux I__1103 (
            .O(N__6449),
            .I(N__6417));
    InMux I__1102 (
            .O(N__6446),
            .I(N__6417));
    InMux I__1101 (
            .O(N__6445),
            .I(N__6412));
    InMux I__1100 (
            .O(N__6442),
            .I(N__6412));
    LocalMux I__1099 (
            .O(N__6439),
            .I(N__6401));
    LocalMux I__1098 (
            .O(N__6436),
            .I(N__6401));
    LocalMux I__1097 (
            .O(N__6433),
            .I(N__6401));
    LocalMux I__1096 (
            .O(N__6428),
            .I(N__6401));
    InMux I__1095 (
            .O(N__6425),
            .I(N__6396));
    InMux I__1094 (
            .O(N__6422),
            .I(N__6396));
    LocalMux I__1093 (
            .O(N__6417),
            .I(N__6391));
    LocalMux I__1092 (
            .O(N__6412),
            .I(N__6391));
    InMux I__1091 (
            .O(N__6411),
            .I(N__6386));
    InMux I__1090 (
            .O(N__6410),
            .I(N__6386));
    Span4Mux_v I__1089 (
            .O(N__6401),
            .I(N__6383));
    LocalMux I__1088 (
            .O(N__6396),
            .I(N__6380));
    Span4Mux_v I__1087 (
            .O(N__6391),
            .I(N__6375));
    LocalMux I__1086 (
            .O(N__6386),
            .I(N__6375));
    Span4Mux_h I__1085 (
            .O(N__6383),
            .I(N__6372));
    Span4Mux_v I__1084 (
            .O(N__6380),
            .I(N__6369));
    Sp12to4 I__1083 (
            .O(N__6375),
            .I(N__6362));
    Sp12to4 I__1082 (
            .O(N__6372),
            .I(N__6362));
    Sp12to4 I__1081 (
            .O(N__6369),
            .I(N__6362));
    Odrv12 I__1080 (
            .O(N__6362),
            .I(A_c_4));
    IoInMux I__1079 (
            .O(N__6359),
            .I(N__6356));
    LocalMux I__1078 (
            .O(N__6356),
            .I(N__6353));
    Span4Mux_s3_v I__1077 (
            .O(N__6353),
            .I(N__6350));
    Span4Mux_v I__1076 (
            .O(N__6350),
            .I(N__6347));
    Span4Mux_v I__1075 (
            .O(N__6347),
            .I(N__6344));
    Odrv4 I__1074 (
            .O(N__6344),
            .I(D_OUT_1));
    InMux I__1073 (
            .O(N__6341),
            .I(N__6338));
    LocalMux I__1072 (
            .O(N__6338),
            .I(N__6335));
    Span4Mux_v I__1071 (
            .O(N__6335),
            .I(N__6332));
    Span4Mux_v I__1070 (
            .O(N__6332),
            .I(N__6329));
    Odrv4 I__1069 (
            .O(N__6329),
            .I(\U409_AUTOCONFIG.LIDE_OUT_RNIBHMPZ0Z_3 ));
    IoInMux I__1068 (
            .O(N__6326),
            .I(N__6323));
    LocalMux I__1067 (
            .O(N__6323),
            .I(N__6320));
    IoSpan4Mux I__1066 (
            .O(N__6320),
            .I(N__6317));
    Span4Mux_s3_v I__1065 (
            .O(N__6317),
            .I(N__6314));
    Span4Mux_v I__1064 (
            .O(N__6314),
            .I(N__6311));
    Odrv4 I__1063 (
            .O(N__6311),
            .I(D_OUT_3));
    InMux I__1062 (
            .O(N__6308),
            .I(N__6302));
    InMux I__1061 (
            .O(N__6307),
            .I(N__6302));
    LocalMux I__1060 (
            .O(N__6302),
            .I(\U409_AUTOCONFIG.CONFIGENn_1_sqmuxa ));
    IoInMux I__1059 (
            .O(N__6299),
            .I(N__6296));
    LocalMux I__1058 (
            .O(N__6296),
            .I(N__6293));
    Span4Mux_s0_v I__1057 (
            .O(N__6293),
            .I(N__6290));
    Sp12to4 I__1056 (
            .O(N__6290),
            .I(N__6287));
    Span12Mux_h I__1055 (
            .O(N__6287),
            .I(N__6284));
    Span12Mux_v I__1054 (
            .O(N__6284),
            .I(N__6280));
    InMux I__1053 (
            .O(N__6283),
            .I(N__6277));
    Odrv12 I__1052 (
            .O(N__6280),
            .I(CONFIGENn_c));
    LocalMux I__1051 (
            .O(N__6277),
            .I(CONFIGENn_c));
    CascadeMux I__1050 (
            .O(N__6272),
            .I(\U409_AUTOCONFIG.STATE_ns_1_cascade_ ));
    InMux I__1049 (
            .O(N__6269),
            .I(N__6263));
    InMux I__1048 (
            .O(N__6268),
            .I(N__6260));
    InMux I__1047 (
            .O(N__6267),
            .I(N__6257));
    InMux I__1046 (
            .O(N__6266),
            .I(N__6254));
    LocalMux I__1045 (
            .O(N__6263),
            .I(N__6248));
    LocalMux I__1044 (
            .O(N__6260),
            .I(N__6248));
    LocalMux I__1043 (
            .O(N__6257),
            .I(N__6239));
    LocalMux I__1042 (
            .O(N__6254),
            .I(N__6239));
    InMux I__1041 (
            .O(N__6253),
            .I(N__6235));
    Span4Mux_v I__1040 (
            .O(N__6248),
            .I(N__6232));
    InMux I__1039 (
            .O(N__6247),
            .I(N__6225));
    InMux I__1038 (
            .O(N__6246),
            .I(N__6225));
    InMux I__1037 (
            .O(N__6245),
            .I(N__6225));
    InMux I__1036 (
            .O(N__6244),
            .I(N__6222));
    Span4Mux_v I__1035 (
            .O(N__6239),
            .I(N__6219));
    InMux I__1034 (
            .O(N__6238),
            .I(N__6216));
    LocalMux I__1033 (
            .O(N__6235),
            .I(N__6203));
    Sp12to4 I__1032 (
            .O(N__6232),
            .I(N__6203));
    LocalMux I__1031 (
            .O(N__6225),
            .I(N__6203));
    LocalMux I__1030 (
            .O(N__6222),
            .I(N__6203));
    Sp12to4 I__1029 (
            .O(N__6219),
            .I(N__6203));
    LocalMux I__1028 (
            .O(N__6216),
            .I(N__6203));
    Span12Mux_h I__1027 (
            .O(N__6203),
            .I(N__6200));
    Span12Mux_v I__1026 (
            .O(N__6200),
            .I(N__6197));
    Odrv12 I__1025 (
            .O(N__6197),
            .I(A_c_22));
    InMux I__1024 (
            .O(N__6194),
            .I(N__6191));
    LocalMux I__1023 (
            .O(N__6191),
            .I(N__6188));
    Odrv4 I__1022 (
            .O(N__6188),
            .I(\U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_1 ));
    CascadeMux I__1021 (
            .O(N__6185),
            .I(N__6180));
    InMux I__1020 (
            .O(N__6184),
            .I(N__6177));
    InMux I__1019 (
            .O(N__6183),
            .I(N__6174));
    InMux I__1018 (
            .O(N__6180),
            .I(N__6171));
    LocalMux I__1017 (
            .O(N__6177),
            .I(N__6166));
    LocalMux I__1016 (
            .O(N__6174),
            .I(N__6166));
    LocalMux I__1015 (
            .O(N__6171),
            .I(N__6163));
    Span4Mux_v I__1014 (
            .O(N__6166),
            .I(N__6160));
    Span4Mux_v I__1013 (
            .O(N__6163),
            .I(N__6157));
    Sp12to4 I__1012 (
            .O(N__6160),
            .I(N__6152));
    Sp12to4 I__1011 (
            .O(N__6157),
            .I(N__6152));
    Span12Mux_h I__1010 (
            .O(N__6152),
            .I(N__6149));
    Span12Mux_v I__1009 (
            .O(N__6149),
            .I(N__6146));
    Odrv12 I__1008 (
            .O(N__6146),
            .I(OVL_c));
    CascadeMux I__1007 (
            .O(N__6143),
            .I(N__6140));
    InMux I__1006 (
            .O(N__6140),
            .I(N__6132));
    InMux I__1005 (
            .O(N__6139),
            .I(N__6128));
    InMux I__1004 (
            .O(N__6138),
            .I(N__6121));
    InMux I__1003 (
            .O(N__6137),
            .I(N__6121));
    InMux I__1002 (
            .O(N__6136),
            .I(N__6121));
    CascadeMux I__1001 (
            .O(N__6135),
            .I(N__6118));
    LocalMux I__1000 (
            .O(N__6132),
            .I(N__6114));
    InMux I__999 (
            .O(N__6131),
            .I(N__6111));
    LocalMux I__998 (
            .O(N__6128),
            .I(N__6106));
    LocalMux I__997 (
            .O(N__6121),
            .I(N__6106));
    InMux I__996 (
            .O(N__6118),
            .I(N__6101));
    InMux I__995 (
            .O(N__6117),
            .I(N__6101));
    Span4Mux_v I__994 (
            .O(N__6114),
            .I(N__6098));
    LocalMux I__993 (
            .O(N__6111),
            .I(N__6095));
    Span4Mux_h I__992 (
            .O(N__6106),
            .I(N__6090));
    LocalMux I__991 (
            .O(N__6101),
            .I(N__6090));
    Span4Mux_h I__990 (
            .O(N__6098),
            .I(N__6085));
    Span4Mux_v I__989 (
            .O(N__6095),
            .I(N__6085));
    Span4Mux_h I__988 (
            .O(N__6090),
            .I(N__6082));
    Span4Mux_v I__987 (
            .O(N__6085),
            .I(N__6079));
    Span4Mux_v I__986 (
            .O(N__6082),
            .I(N__6076));
    Sp12to4 I__985 (
            .O(N__6079),
            .I(N__6071));
    Sp12to4 I__984 (
            .O(N__6076),
            .I(N__6071));
    Odrv12 I__983 (
            .O(N__6071),
            .I(A_c_23));
    IoInMux I__982 (
            .O(N__6068),
            .I(N__6065));
    LocalMux I__981 (
            .O(N__6065),
            .I(N__6062));
    Span4Mux_s3_v I__980 (
            .O(N__6062),
            .I(N__6059));
    Span4Mux_h I__979 (
            .O(N__6059),
            .I(N__6056));
    Sp12to4 I__978 (
            .O(N__6056),
            .I(N__6053));
    Odrv12 I__977 (
            .O(N__6053),
            .I(U409_ADDRESS_DECODE_un1_RAMSPACEn_i));
    InMux I__976 (
            .O(N__6050),
            .I(N__6044));
    InMux I__975 (
            .O(N__6049),
            .I(N__6039));
    InMux I__974 (
            .O(N__6048),
            .I(N__6036));
    InMux I__973 (
            .O(N__6047),
            .I(N__6033));
    LocalMux I__972 (
            .O(N__6044),
            .I(N__6030));
    InMux I__971 (
            .O(N__6043),
            .I(N__6025));
    InMux I__970 (
            .O(N__6042),
            .I(N__6025));
    LocalMux I__969 (
            .O(N__6039),
            .I(N__6022));
    LocalMux I__968 (
            .O(N__6036),
            .I(\U409_AUTOCONFIG.STATEZ0Z_1 ));
    LocalMux I__967 (
            .O(N__6033),
            .I(\U409_AUTOCONFIG.STATEZ0Z_1 ));
    Odrv4 I__966 (
            .O(N__6030),
            .I(\U409_AUTOCONFIG.STATEZ0Z_1 ));
    LocalMux I__965 (
            .O(N__6025),
            .I(\U409_AUTOCONFIG.STATEZ0Z_1 ));
    Odrv4 I__964 (
            .O(N__6022),
            .I(\U409_AUTOCONFIG.STATEZ0Z_1 ));
    InMux I__963 (
            .O(N__6011),
            .I(N__6002));
    InMux I__962 (
            .O(N__6010),
            .I(N__6002));
    InMux I__961 (
            .O(N__6009),
            .I(N__6002));
    LocalMux I__960 (
            .O(N__6002),
            .I(N__5996));
    InMux I__959 (
            .O(N__6001),
            .I(N__5993));
    CascadeMux I__958 (
            .O(N__6000),
            .I(N__5990));
    CascadeMux I__957 (
            .O(N__5999),
            .I(N__5986));
    Span4Mux_v I__956 (
            .O(N__5996),
            .I(N__5976));
    LocalMux I__955 (
            .O(N__5993),
            .I(N__5976));
    InMux I__954 (
            .O(N__5990),
            .I(N__5971));
    InMux I__953 (
            .O(N__5989),
            .I(N__5971));
    InMux I__952 (
            .O(N__5986),
            .I(N__5968));
    InMux I__951 (
            .O(N__5985),
            .I(N__5965));
    InMux I__950 (
            .O(N__5984),
            .I(N__5962));
    InMux I__949 (
            .O(N__5983),
            .I(N__5959));
    InMux I__948 (
            .O(N__5982),
            .I(N__5954));
    InMux I__947 (
            .O(N__5981),
            .I(N__5954));
    Span4Mux_h I__946 (
            .O(N__5976),
            .I(N__5949));
    LocalMux I__945 (
            .O(N__5971),
            .I(N__5949));
    LocalMux I__944 (
            .O(N__5968),
            .I(N__5938));
    LocalMux I__943 (
            .O(N__5965),
            .I(N__5938));
    LocalMux I__942 (
            .O(N__5962),
            .I(N__5938));
    LocalMux I__941 (
            .O(N__5959),
            .I(N__5938));
    LocalMux I__940 (
            .O(N__5954),
            .I(N__5938));
    Span4Mux_v I__939 (
            .O(N__5949),
            .I(N__5935));
    Span4Mux_v I__938 (
            .O(N__5938),
            .I(N__5932));
    Span4Mux_v I__937 (
            .O(N__5935),
            .I(N__5929));
    Sp12to4 I__936 (
            .O(N__5932),
            .I(N__5926));
    Sp12to4 I__935 (
            .O(N__5929),
            .I(N__5923));
    Span12Mux_h I__934 (
            .O(N__5926),
            .I(N__5920));
    Span12Mux_h I__933 (
            .O(N__5923),
            .I(N__5915));
    Span12Mux_v I__932 (
            .O(N__5920),
            .I(N__5915));
    Odrv12 I__931 (
            .O(N__5915),
            .I(RnW_c));
    CascadeMux I__930 (
            .O(N__5912),
            .I(N__5909));
    InMux I__929 (
            .O(N__5909),
            .I(N__5906));
    LocalMux I__928 (
            .O(N__5906),
            .I(N__5902));
    InMux I__927 (
            .O(N__5905),
            .I(N__5899));
    Span4Mux_h I__926 (
            .O(N__5902),
            .I(N__5894));
    LocalMux I__925 (
            .O(N__5899),
            .I(N__5894));
    Span4Mux_v I__924 (
            .O(N__5894),
            .I(N__5891));
    Sp12to4 I__923 (
            .O(N__5891),
            .I(N__5888));
    Span12Mux_h I__922 (
            .O(N__5888),
            .I(N__5885));
    Span12Mux_v I__921 (
            .O(N__5885),
            .I(N__5882));
    Odrv12 I__920 (
            .O(N__5882),
            .I(CPUCONFn_c));
    CascadeMux I__919 (
            .O(N__5879),
            .I(\U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_a3_1_cascade_ ));
    CascadeMux I__918 (
            .O(N__5876),
            .I(\U409_AUTOCONFIG.N_227_3_cascade_ ));
    CascadeMux I__917 (
            .O(N__5873),
            .I(N__5870));
    InMux I__916 (
            .O(N__5870),
            .I(N__5867));
    LocalMux I__915 (
            .O(N__5867),
            .I(N__5864));
    Span4Mux_v I__914 (
            .O(N__5864),
            .I(N__5861));
    Sp12to4 I__913 (
            .O(N__5861),
            .I(N__5857));
    InMux I__912 (
            .O(N__5860),
            .I(N__5854));
    Span12Mux_h I__911 (
            .O(N__5857),
            .I(N__5849));
    LocalMux I__910 (
            .O(N__5854),
            .I(N__5849));
    Span12Mux_v I__909 (
            .O(N__5849),
            .I(N__5846));
    Odrv12 I__908 (
            .O(N__5846),
            .I(D_in_5));
    CascadeMux I__907 (
            .O(N__5843),
            .I(\U409_AUTOCONFIG.N_49_cascade_ ));
    InMux I__906 (
            .O(N__5840),
            .I(N__5837));
    LocalMux I__905 (
            .O(N__5837),
            .I(\U409_AUTOCONFIG.N_107 ));
    InMux I__904 (
            .O(N__5834),
            .I(N__5831));
    LocalMux I__903 (
            .O(N__5831),
            .I(\U409_AUTOCONFIG.N_95 ));
    CascadeMux I__902 (
            .O(N__5828),
            .I(\U409_AUTOCONFIG.N_48_cascade_ ));
    InMux I__901 (
            .O(N__5825),
            .I(N__5822));
    LocalMux I__900 (
            .O(N__5822),
            .I(N__5818));
    InMux I__899 (
            .O(N__5821),
            .I(N__5815));
    Span4Mux_h I__898 (
            .O(N__5818),
            .I(N__5810));
    LocalMux I__897 (
            .O(N__5815),
            .I(N__5810));
    Span4Mux_v I__896 (
            .O(N__5810),
            .I(N__5807));
    Odrv4 I__895 (
            .O(N__5807),
            .I(\U409_AUTOCONFIG.un1_A_13 ));
    InMux I__894 (
            .O(N__5804),
            .I(N__5801));
    LocalMux I__893 (
            .O(N__5801),
            .I(\U409_AUTOCONFIG.STATE_d_2 ));
    InMux I__892 (
            .O(N__5798),
            .I(N__5792));
    InMux I__891 (
            .O(N__5797),
            .I(N__5792));
    LocalMux I__890 (
            .O(N__5792),
            .I(LIDE_BASE_7));
    InMux I__889 (
            .O(N__5789),
            .I(N__5786));
    LocalMux I__888 (
            .O(N__5786),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_4 ));
    CascadeMux I__887 (
            .O(N__5783),
            .I(N__5776));
    CascadeMux I__886 (
            .O(N__5782),
            .I(N__5773));
    CascadeMux I__885 (
            .O(N__5781),
            .I(N__5770));
    CascadeMux I__884 (
            .O(N__5780),
            .I(N__5766));
    InMux I__883 (
            .O(N__5779),
            .I(N__5763));
    InMux I__882 (
            .O(N__5776),
            .I(N__5757));
    InMux I__881 (
            .O(N__5773),
            .I(N__5757));
    InMux I__880 (
            .O(N__5770),
            .I(N__5750));
    InMux I__879 (
            .O(N__5769),
            .I(N__5750));
    InMux I__878 (
            .O(N__5766),
            .I(N__5750));
    LocalMux I__877 (
            .O(N__5763),
            .I(N__5746));
    InMux I__876 (
            .O(N__5762),
            .I(N__5743));
    LocalMux I__875 (
            .O(N__5757),
            .I(N__5740));
    LocalMux I__874 (
            .O(N__5750),
            .I(N__5737));
    InMux I__873 (
            .O(N__5749),
            .I(N__5734));
    Span4Mux_v I__872 (
            .O(N__5746),
            .I(N__5729));
    LocalMux I__871 (
            .O(N__5743),
            .I(N__5729));
    Odrv4 I__870 (
            .O(N__5740),
            .I(\U409_AUTOCONFIG.un1_STATE_6_0 ));
    Odrv4 I__869 (
            .O(N__5737),
            .I(\U409_AUTOCONFIG.un1_STATE_6_0 ));
    LocalMux I__868 (
            .O(N__5734),
            .I(\U409_AUTOCONFIG.un1_STATE_6_0 ));
    Odrv4 I__867 (
            .O(N__5729),
            .I(\U409_AUTOCONFIG.un1_STATE_6_0 ));
    InMux I__866 (
            .O(N__5720),
            .I(N__5713));
    InMux I__865 (
            .O(N__5719),
            .I(N__5713));
    InMux I__864 (
            .O(N__5718),
            .I(N__5706));
    LocalMux I__863 (
            .O(N__5713),
            .I(N__5703));
    InMux I__862 (
            .O(N__5712),
            .I(N__5698));
    InMux I__861 (
            .O(N__5711),
            .I(N__5698));
    InMux I__860 (
            .O(N__5710),
            .I(N__5694));
    InMux I__859 (
            .O(N__5709),
            .I(N__5691));
    LocalMux I__858 (
            .O(N__5706),
            .I(N__5684));
    Span4Mux_v I__857 (
            .O(N__5703),
            .I(N__5684));
    LocalMux I__856 (
            .O(N__5698),
            .I(N__5684));
    InMux I__855 (
            .O(N__5697),
            .I(N__5681));
    LocalMux I__854 (
            .O(N__5694),
            .I(\U409_AUTOCONFIG.N_48 ));
    LocalMux I__853 (
            .O(N__5691),
            .I(\U409_AUTOCONFIG.N_48 ));
    Odrv4 I__852 (
            .O(N__5684),
            .I(\U409_AUTOCONFIG.N_48 ));
    LocalMux I__851 (
            .O(N__5681),
            .I(\U409_AUTOCONFIG.N_48 ));
    CascadeMux I__850 (
            .O(N__5672),
            .I(N__5669));
    InMux I__849 (
            .O(N__5669),
            .I(N__5658));
    InMux I__848 (
            .O(N__5668),
            .I(N__5658));
    InMux I__847 (
            .O(N__5667),
            .I(N__5658));
    InMux I__846 (
            .O(N__5666),
            .I(N__5655));
    InMux I__845 (
            .O(N__5665),
            .I(N__5652));
    LocalMux I__844 (
            .O(N__5658),
            .I(N__5649));
    LocalMux I__843 (
            .O(N__5655),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    LocalMux I__842 (
            .O(N__5652),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    Odrv4 I__841 (
            .O(N__5649),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    InMux I__840 (
            .O(N__5642),
            .I(N__5639));
    LocalMux I__839 (
            .O(N__5639),
            .I(N__5636));
    Odrv4 I__838 (
            .O(N__5636),
            .I(\U409_ADDRESS_DECODE.LOWROMZ0Z_3 ));
    CascadeMux I__837 (
            .O(N__5633),
            .I(N__5628));
    CascadeMux I__836 (
            .O(N__5632),
            .I(N__5625));
    CascadeMux I__835 (
            .O(N__5631),
            .I(N__5620));
    InMux I__834 (
            .O(N__5628),
            .I(N__5614));
    InMux I__833 (
            .O(N__5625),
            .I(N__5609));
    InMux I__832 (
            .O(N__5624),
            .I(N__5609));
    InMux I__831 (
            .O(N__5623),
            .I(N__5604));
    InMux I__830 (
            .O(N__5620),
            .I(N__5604));
    InMux I__829 (
            .O(N__5619),
            .I(N__5600));
    InMux I__828 (
            .O(N__5618),
            .I(N__5597));
    InMux I__827 (
            .O(N__5617),
            .I(N__5594));
    LocalMux I__826 (
            .O(N__5614),
            .I(N__5587));
    LocalMux I__825 (
            .O(N__5609),
            .I(N__5587));
    LocalMux I__824 (
            .O(N__5604),
            .I(N__5587));
    InMux I__823 (
            .O(N__5603),
            .I(N__5584));
    LocalMux I__822 (
            .O(N__5600),
            .I(N__5576));
    LocalMux I__821 (
            .O(N__5597),
            .I(N__5576));
    LocalMux I__820 (
            .O(N__5594),
            .I(N__5576));
    Span4Mux_v I__819 (
            .O(N__5587),
            .I(N__5571));
    LocalMux I__818 (
            .O(N__5584),
            .I(N__5571));
    InMux I__817 (
            .O(N__5583),
            .I(N__5568));
    Span4Mux_v I__816 (
            .O(N__5576),
            .I(N__5565));
    Span4Mux_h I__815 (
            .O(N__5571),
            .I(N__5560));
    LocalMux I__814 (
            .O(N__5568),
            .I(N__5560));
    Span4Mux_v I__813 (
            .O(N__5565),
            .I(N__5557));
    Span4Mux_v I__812 (
            .O(N__5560),
            .I(N__5554));
    Sp12to4 I__811 (
            .O(N__5557),
            .I(N__5549));
    Sp12to4 I__810 (
            .O(N__5554),
            .I(N__5549));
    Odrv12 I__809 (
            .O(N__5549),
            .I(A_c_21));
    InMux I__808 (
            .O(N__5546),
            .I(N__5542));
    InMux I__807 (
            .O(N__5545),
            .I(N__5537));
    LocalMux I__806 (
            .O(N__5542),
            .I(N__5533));
    InMux I__805 (
            .O(N__5541),
            .I(N__5530));
    InMux I__804 (
            .O(N__5540),
            .I(N__5527));
    LocalMux I__803 (
            .O(N__5537),
            .I(N__5524));
    InMux I__802 (
            .O(N__5536),
            .I(N__5521));
    Span4Mux_v I__801 (
            .O(N__5533),
            .I(N__5512));
    LocalMux I__800 (
            .O(N__5530),
            .I(N__5512));
    LocalMux I__799 (
            .O(N__5527),
            .I(N__5512));
    Span4Mux_h I__798 (
            .O(N__5524),
            .I(N__5507));
    LocalMux I__797 (
            .O(N__5521),
            .I(N__5507));
    InMux I__796 (
            .O(N__5520),
            .I(N__5504));
    InMux I__795 (
            .O(N__5519),
            .I(N__5501));
    Span4Mux_v I__794 (
            .O(N__5512),
            .I(N__5498));
    Span4Mux_v I__793 (
            .O(N__5507),
            .I(N__5495));
    LocalMux I__792 (
            .O(N__5504),
            .I(N__5492));
    LocalMux I__791 (
            .O(N__5501),
            .I(N__5489));
    Sp12to4 I__790 (
            .O(N__5498),
            .I(N__5482));
    Sp12to4 I__789 (
            .O(N__5495),
            .I(N__5482));
    Span12Mux_v I__788 (
            .O(N__5492),
            .I(N__5482));
    Span12Mux_h I__787 (
            .O(N__5489),
            .I(N__5479));
    Odrv12 I__786 (
            .O(N__5482),
            .I(A_c_20));
    Odrv12 I__785 (
            .O(N__5479),
            .I(A_c_20));
    CascadeMux I__784 (
            .O(N__5474),
            .I(N__5471));
    InMux I__783 (
            .O(N__5471),
            .I(N__5468));
    LocalMux I__782 (
            .O(N__5468),
            .I(N__5465));
    Odrv4 I__781 (
            .O(N__5465),
            .I(\U409_AUTOCONFIG.PR_OUTZ0Z_2 ));
    IoInMux I__780 (
            .O(N__5462),
            .I(N__5459));
    LocalMux I__779 (
            .O(N__5459),
            .I(N__5456));
    Span12Mux_s6_v I__778 (
            .O(N__5456),
            .I(N__5453));
    Odrv12 I__777 (
            .O(N__5453),
            .I(D_OUT_2));
    InMux I__776 (
            .O(N__5450),
            .I(N__5447));
    LocalMux I__775 (
            .O(N__5447),
            .I(N__5444));
    Span4Mux_h I__774 (
            .O(N__5444),
            .I(N__5441));
    Odrv4 I__773 (
            .O(N__5441),
            .I(\U409_AUTOCONFIG.N_97 ));
    CascadeMux I__772 (
            .O(N__5438),
            .I(\U409_AUTOCONFIG.STATE_d_2_cascade_ ));
    InMux I__771 (
            .O(N__5435),
            .I(N__5429));
    InMux I__770 (
            .O(N__5434),
            .I(N__5429));
    LocalMux I__769 (
            .O(N__5429),
            .I(N__5426));
    Span12Mux_v I__768 (
            .O(N__5426),
            .I(N__5423));
    Odrv12 I__767 (
            .O(N__5423),
            .I(D_in_6));
    InMux I__766 (
            .O(N__5420),
            .I(N__5417));
    LocalMux I__765 (
            .O(N__5417),
            .I(\U409_AUTOCONFIG.N_105 ));
    InMux I__764 (
            .O(N__5414),
            .I(N__5411));
    LocalMux I__763 (
            .O(N__5411),
            .I(N__5404));
    InMux I__762 (
            .O(N__5410),
            .I(N__5399));
    InMux I__761 (
            .O(N__5409),
            .I(N__5399));
    InMux I__760 (
            .O(N__5408),
            .I(N__5396));
    InMux I__759 (
            .O(N__5407),
            .I(N__5393));
    Odrv12 I__758 (
            .O(N__5404),
            .I(\U409_AUTOCONFIG.N_49 ));
    LocalMux I__757 (
            .O(N__5399),
            .I(\U409_AUTOCONFIG.N_49 ));
    LocalMux I__756 (
            .O(N__5396),
            .I(\U409_AUTOCONFIG.N_49 ));
    LocalMux I__755 (
            .O(N__5393),
            .I(\U409_AUTOCONFIG.N_49 ));
    InMux I__754 (
            .O(N__5384),
            .I(N__5381));
    LocalMux I__753 (
            .O(N__5381),
            .I(\U409_AUTOCONFIG.PR_OUT_cnst_i_i_0_0_2 ));
    CascadeMux I__752 (
            .O(N__5378),
            .I(\U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_1_cascade_ ));
    CascadeMux I__751 (
            .O(N__5375),
            .I(N__5372));
    InMux I__750 (
            .O(N__5372),
            .I(N__5365));
    InMux I__749 (
            .O(N__5371),
            .I(N__5360));
    InMux I__748 (
            .O(N__5370),
            .I(N__5360));
    InMux I__747 (
            .O(N__5369),
            .I(N__5356));
    InMux I__746 (
            .O(N__5368),
            .I(N__5353));
    LocalMux I__745 (
            .O(N__5365),
            .I(N__5348));
    LocalMux I__744 (
            .O(N__5360),
            .I(N__5348));
    CascadeMux I__743 (
            .O(N__5359),
            .I(N__5345));
    LocalMux I__742 (
            .O(N__5356),
            .I(N__5340));
    LocalMux I__741 (
            .O(N__5353),
            .I(N__5340));
    Span4Mux_v I__740 (
            .O(N__5348),
            .I(N__5337));
    InMux I__739 (
            .O(N__5345),
            .I(N__5334));
    Span4Mux_v I__738 (
            .O(N__5340),
            .I(N__5331));
    Sp12to4 I__737 (
            .O(N__5337),
            .I(N__5324));
    LocalMux I__736 (
            .O(N__5334),
            .I(N__5324));
    Sp12to4 I__735 (
            .O(N__5331),
            .I(N__5324));
    Span12Mux_h I__734 (
            .O(N__5324),
            .I(N__5321));
    Span12Mux_v I__733 (
            .O(N__5321),
            .I(N__5318));
    Odrv12 I__732 (
            .O(N__5318),
            .I(A_c_19));
    InMux I__731 (
            .O(N__5315),
            .I(N__5309));
    InMux I__730 (
            .O(N__5314),
            .I(N__5309));
    LocalMux I__729 (
            .O(N__5309),
            .I(\U409_AUTOCONFIG.N_84 ));
    InMux I__728 (
            .O(N__5306),
            .I(N__5303));
    LocalMux I__727 (
            .O(N__5303),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ));
    InMux I__726 (
            .O(N__5300),
            .I(N__5297));
    LocalMux I__725 (
            .O(N__5297),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ));
    InMux I__724 (
            .O(N__5294),
            .I(N__5291));
    LocalMux I__723 (
            .O(N__5291),
            .I(N__5287));
    InMux I__722 (
            .O(N__5290),
            .I(N__5284));
    Span4Mux_v I__721 (
            .O(N__5287),
            .I(N__5281));
    LocalMux I__720 (
            .O(N__5284),
            .I(N__5278));
    Span4Mux_h I__719 (
            .O(N__5281),
            .I(N__5273));
    Span4Mux_h I__718 (
            .O(N__5278),
            .I(N__5273));
    Span4Mux_v I__717 (
            .O(N__5273),
            .I(N__5270));
    Span4Mux_v I__716 (
            .O(N__5270),
            .I(N__5267));
    Odrv4 I__715 (
            .O(N__5267),
            .I(D_in_7));
    InMux I__714 (
            .O(N__5264),
            .I(N__5261));
    LocalMux I__713 (
            .O(N__5261),
            .I(\U409_ADDRESS_DECODE.PORTSIZEZ0Z_1 ));
    CascadeMux I__712 (
            .O(N__5258),
            .I(\U409_ADDRESS_DECODE.PORTSIZEZ0Z_0_cascade_ ));
    IoInMux I__711 (
            .O(N__5255),
            .I(N__5252));
    LocalMux I__710 (
            .O(N__5252),
            .I(N__5249));
    IoSpan4Mux I__709 (
            .O(N__5249),
            .I(N__5246));
    Span4Mux_s2_v I__708 (
            .O(N__5246),
            .I(N__5243));
    Sp12to4 I__707 (
            .O(N__5243),
            .I(N__5240));
    Span12Mux_s8_v I__706 (
            .O(N__5240),
            .I(N__5237));
    Odrv12 I__705 (
            .O(N__5237),
            .I(PORTSIZE_0_i));
    IoInMux I__704 (
            .O(N__5234),
            .I(N__5231));
    LocalMux I__703 (
            .O(N__5231),
            .I(N__5228));
    Span4Mux_s3_v I__702 (
            .O(N__5228),
            .I(N__5225));
    Span4Mux_v I__701 (
            .O(N__5225),
            .I(N__5222));
    Sp12to4 I__700 (
            .O(N__5222),
            .I(N__5219));
    Span12Mux_h I__699 (
            .O(N__5219),
            .I(N__5216));
    Odrv12 I__698 (
            .O(N__5216),
            .I(BUFENn_c));
    IoInMux I__697 (
            .O(N__5213),
            .I(N__5210));
    LocalMux I__696 (
            .O(N__5210),
            .I(N__5207));
    IoSpan4Mux I__695 (
            .O(N__5207),
            .I(N__5204));
    Span4Mux_s2_h I__694 (
            .O(N__5204),
            .I(N__5201));
    Sp12to4 I__693 (
            .O(N__5201),
            .I(N__5198));
    Span12Mux_s9_h I__692 (
            .O(N__5198),
            .I(N__5195));
    Odrv12 I__691 (
            .O(N__5195),
            .I(U409_ADDRESS_DECODE_un1_ATA_ENn_i));
    CascadeMux I__690 (
            .O(N__5192),
            .I(N__5188));
    InMux I__689 (
            .O(N__5191),
            .I(N__5183));
    InMux I__688 (
            .O(N__5188),
            .I(N__5180));
    InMux I__687 (
            .O(N__5187),
            .I(N__5177));
    InMux I__686 (
            .O(N__5186),
            .I(N__5174));
    LocalMux I__685 (
            .O(N__5183),
            .I(N__5169));
    LocalMux I__684 (
            .O(N__5180),
            .I(N__5169));
    LocalMux I__683 (
            .O(N__5177),
            .I(N__5164));
    LocalMux I__682 (
            .O(N__5174),
            .I(N__5164));
    Span4Mux_h I__681 (
            .O(N__5169),
            .I(N__5161));
    Span12Mux_h I__680 (
            .O(N__5164),
            .I(N__5156));
    Sp12to4 I__679 (
            .O(N__5161),
            .I(N__5156));
    Span12Mux_v I__678 (
            .O(N__5156),
            .I(N__5153));
    Odrv12 I__677 (
            .O(N__5153),
            .I(A_c_18));
    InMux I__676 (
            .O(N__5150),
            .I(N__5146));
    InMux I__675 (
            .O(N__5149),
            .I(N__5143));
    LocalMux I__674 (
            .O(N__5146),
            .I(LIDE_BASE_2));
    LocalMux I__673 (
            .O(N__5143),
            .I(LIDE_BASE_2));
    CascadeMux I__672 (
            .O(N__5138),
            .I(N__5134));
    CascadeMux I__671 (
            .O(N__5137),
            .I(N__5131));
    InMux I__670 (
            .O(N__5134),
            .I(N__5128));
    InMux I__669 (
            .O(N__5131),
            .I(N__5122));
    LocalMux I__668 (
            .O(N__5128),
            .I(N__5119));
    InMux I__667 (
            .O(N__5127),
            .I(N__5116));
    InMux I__666 (
            .O(N__5126),
            .I(N__5113));
    InMux I__665 (
            .O(N__5125),
            .I(N__5110));
    LocalMux I__664 (
            .O(N__5122),
            .I(N__5107));
    Span4Mux_h I__663 (
            .O(N__5119),
            .I(N__5100));
    LocalMux I__662 (
            .O(N__5116),
            .I(N__5100));
    LocalMux I__661 (
            .O(N__5113),
            .I(N__5100));
    LocalMux I__660 (
            .O(N__5110),
            .I(N__5093));
    Sp12to4 I__659 (
            .O(N__5107),
            .I(N__5093));
    Sp12to4 I__658 (
            .O(N__5100),
            .I(N__5093));
    Span12Mux_v I__657 (
            .O(N__5093),
            .I(N__5090));
    Odrv12 I__656 (
            .O(N__5090),
            .I(A_c_17));
    InMux I__655 (
            .O(N__5087),
            .I(N__5083));
    InMux I__654 (
            .O(N__5086),
            .I(N__5080));
    LocalMux I__653 (
            .O(N__5083),
            .I(LIDE_BASE_1));
    LocalMux I__652 (
            .O(N__5080),
            .I(LIDE_BASE_1));
    InMux I__651 (
            .O(N__5075),
            .I(N__5072));
    LocalMux I__650 (
            .O(N__5072),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3 ));
    CascadeMux I__649 (
            .O(N__5069),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1_cascade_ ));
    InMux I__648 (
            .O(N__5066),
            .I(N__5063));
    LocalMux I__647 (
            .O(N__5063),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2 ));
    InMux I__646 (
            .O(N__5060),
            .I(N__5051));
    InMux I__645 (
            .O(N__5059),
            .I(N__5051));
    InMux I__644 (
            .O(N__5058),
            .I(N__5051));
    LocalMux I__643 (
            .O(N__5051),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0 ));
    CascadeMux I__642 (
            .O(N__5048),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_ ));
    InMux I__641 (
            .O(N__5045),
            .I(N__5036));
    InMux I__640 (
            .O(N__5044),
            .I(N__5036));
    InMux I__639 (
            .O(N__5043),
            .I(N__5036));
    LocalMux I__638 (
            .O(N__5036),
            .I(\U409_ADDRESS_DECODE.ATA_ENZ0 ));
    CascadeMux I__637 (
            .O(N__5033),
            .I(\U409_AUTOCONFIG.N_121_cascade_ ));
    InMux I__636 (
            .O(N__5030),
            .I(N__5025));
    InMux I__635 (
            .O(N__5029),
            .I(N__5021));
    InMux I__634 (
            .O(N__5028),
            .I(N__5018));
    LocalMux I__633 (
            .O(N__5025),
            .I(N__5015));
    CascadeMux I__632 (
            .O(N__5024),
            .I(N__5012));
    LocalMux I__631 (
            .O(N__5021),
            .I(N__5007));
    LocalMux I__630 (
            .O(N__5018),
            .I(N__5007));
    Span4Mux_v I__629 (
            .O(N__5015),
            .I(N__5004));
    InMux I__628 (
            .O(N__5012),
            .I(N__5001));
    Span12Mux_v I__627 (
            .O(N__5007),
            .I(N__4994));
    Sp12to4 I__626 (
            .O(N__5004),
            .I(N__4994));
    LocalMux I__625 (
            .O(N__5001),
            .I(N__4994));
    Odrv12 I__624 (
            .O(N__4994),
            .I(A_c_7));
    InMux I__623 (
            .O(N__4991),
            .I(N__4987));
    InMux I__622 (
            .O(N__4990),
            .I(N__4984));
    LocalMux I__621 (
            .O(N__4987),
            .I(N__4981));
    LocalMux I__620 (
            .O(N__4984),
            .I(N__4978));
    Span4Mux_v I__619 (
            .O(N__4981),
            .I(N__4968));
    Span4Mux_v I__618 (
            .O(N__4978),
            .I(N__4968));
    InMux I__617 (
            .O(N__4977),
            .I(N__4961));
    InMux I__616 (
            .O(N__4976),
            .I(N__4961));
    InMux I__615 (
            .O(N__4975),
            .I(N__4961));
    InMux I__614 (
            .O(N__4974),
            .I(N__4956));
    InMux I__613 (
            .O(N__4973),
            .I(N__4956));
    Sp12to4 I__612 (
            .O(N__4968),
            .I(N__4949));
    LocalMux I__611 (
            .O(N__4961),
            .I(N__4949));
    LocalMux I__610 (
            .O(N__4956),
            .I(N__4949));
    Odrv12 I__609 (
            .O(N__4949),
            .I(A_c_6));
    CascadeMux I__608 (
            .O(N__4946),
            .I(N__4942));
    InMux I__607 (
            .O(N__4945),
            .I(N__4939));
    InMux I__606 (
            .O(N__4942),
            .I(N__4935));
    LocalMux I__605 (
            .O(N__4939),
            .I(N__4932));
    InMux I__604 (
            .O(N__4938),
            .I(N__4929));
    LocalMux I__603 (
            .O(N__4935),
            .I(N__4925));
    Span4Mux_v I__602 (
            .O(N__4932),
            .I(N__4922));
    LocalMux I__601 (
            .O(N__4929),
            .I(N__4919));
    InMux I__600 (
            .O(N__4928),
            .I(N__4916));
    Span12Mux_v I__599 (
            .O(N__4925),
            .I(N__4907));
    Sp12to4 I__598 (
            .O(N__4922),
            .I(N__4907));
    Sp12to4 I__597 (
            .O(N__4919),
            .I(N__4907));
    LocalMux I__596 (
            .O(N__4916),
            .I(N__4907));
    Odrv12 I__595 (
            .O(N__4907),
            .I(A_c_5));
    InMux I__594 (
            .O(N__4904),
            .I(N__4894));
    InMux I__593 (
            .O(N__4903),
            .I(N__4894));
    InMux I__592 (
            .O(N__4902),
            .I(N__4889));
    InMux I__591 (
            .O(N__4901),
            .I(N__4889));
    InMux I__590 (
            .O(N__4900),
            .I(N__4884));
    InMux I__589 (
            .O(N__4899),
            .I(N__4884));
    LocalMux I__588 (
            .O(N__4894),
            .I(N__4879));
    LocalMux I__587 (
            .O(N__4889),
            .I(N__4879));
    LocalMux I__586 (
            .O(N__4884),
            .I(N__4876));
    Sp12to4 I__585 (
            .O(N__4879),
            .I(N__4873));
    Span12Mux_h I__584 (
            .O(N__4876),
            .I(N__4870));
    Span12Mux_v I__583 (
            .O(N__4873),
            .I(N__4867));
    Span12Mux_v I__582 (
            .O(N__4870),
            .I(N__4864));
    Odrv12 I__581 (
            .O(N__4867),
            .I(A_c_3));
    Odrv12 I__580 (
            .O(N__4864),
            .I(A_c_3));
    InMux I__579 (
            .O(N__4859),
            .I(N__4854));
    InMux I__578 (
            .O(N__4858),
            .I(N__4849));
    InMux I__577 (
            .O(N__4857),
            .I(N__4849));
    LocalMux I__576 (
            .O(N__4854),
            .I(\U409_AUTOCONFIG.N_121 ));
    LocalMux I__575 (
            .O(N__4849),
            .I(\U409_AUTOCONFIG.N_121 ));
    CascadeMux I__574 (
            .O(N__4844),
            .I(N__4841));
    InMux I__573 (
            .O(N__4841),
            .I(N__4838));
    LocalMux I__572 (
            .O(N__4838),
            .I(N__4835));
    Odrv12 I__571 (
            .O(N__4835),
            .I(\U409_AUTOCONFIG.N_123 ));
    CascadeMux I__570 (
            .O(N__4832),
            .I(N__4828));
    InMux I__569 (
            .O(N__4831),
            .I(N__4825));
    InMux I__568 (
            .O(N__4828),
            .I(N__4822));
    LocalMux I__567 (
            .O(N__4825),
            .I(N__4819));
    LocalMux I__566 (
            .O(N__4822),
            .I(N__4816));
    Span4Mux_v I__565 (
            .O(N__4819),
            .I(N__4811));
    Span4Mux_v I__564 (
            .O(N__4816),
            .I(N__4808));
    InMux I__563 (
            .O(N__4815),
            .I(N__4805));
    InMux I__562 (
            .O(N__4814),
            .I(N__4802));
    Span4Mux_v I__561 (
            .O(N__4811),
            .I(N__4799));
    Span4Mux_v I__560 (
            .O(N__4808),
            .I(N__4792));
    LocalMux I__559 (
            .O(N__4805),
            .I(N__4792));
    LocalMux I__558 (
            .O(N__4802),
            .I(N__4792));
    Span4Mux_v I__557 (
            .O(N__4799),
            .I(N__4789));
    Span4Mux_v I__556 (
            .O(N__4792),
            .I(N__4786));
    Sp12to4 I__555 (
            .O(N__4789),
            .I(N__4781));
    Sp12to4 I__554 (
            .O(N__4786),
            .I(N__4781));
    Odrv12 I__553 (
            .O(N__4781),
            .I(A_c_16));
    InMux I__552 (
            .O(N__4778),
            .I(N__4774));
    InMux I__551 (
            .O(N__4777),
            .I(N__4771));
    LocalMux I__550 (
            .O(N__4774),
            .I(N__4766));
    LocalMux I__549 (
            .O(N__4771),
            .I(N__4766));
    Span4Mux_v I__548 (
            .O(N__4766),
            .I(N__4763));
    Sp12to4 I__547 (
            .O(N__4763),
            .I(N__4760));
    Odrv12 I__546 (
            .O(N__4760),
            .I(A_c_15));
    IoInMux I__545 (
            .O(N__4757),
            .I(N__4754));
    LocalMux I__544 (
            .O(N__4754),
            .I(N__4749));
    IoInMux I__543 (
            .O(N__4753),
            .I(N__4746));
    IoInMux I__542 (
            .O(N__4752),
            .I(N__4743));
    IoSpan4Mux I__541 (
            .O(N__4749),
            .I(N__4739));
    LocalMux I__540 (
            .O(N__4746),
            .I(N__4734));
    LocalMux I__539 (
            .O(N__4743),
            .I(N__4734));
    IoInMux I__538 (
            .O(N__4742),
            .I(N__4731));
    Span4Mux_s3_v I__537 (
            .O(N__4739),
            .I(N__4728));
    Span4Mux_s3_v I__536 (
            .O(N__4734),
            .I(N__4725));
    LocalMux I__535 (
            .O(N__4731),
            .I(N__4722));
    Span4Mux_v I__534 (
            .O(N__4728),
            .I(N__4717));
    Span4Mux_v I__533 (
            .O(N__4725),
            .I(N__4717));
    Span12Mux_s8_v I__532 (
            .O(N__4722),
            .I(N__4714));
    Odrv4 I__531 (
            .O(N__4717),
            .I(D_1_i));
    Odrv12 I__530 (
            .O(N__4714),
            .I(D_1_i));
    InMux I__529 (
            .O(N__4709),
            .I(N__4706));
    LocalMux I__528 (
            .O(N__4706),
            .I(N__4703));
    Odrv4 I__527 (
            .O(N__4703),
            .I(\U409_AUTOCONFIG.N_103 ));
    CascadeMux I__526 (
            .O(N__4700),
            .I(N__4697));
    InMux I__525 (
            .O(N__4697),
            .I(N__4694));
    LocalMux I__524 (
            .O(N__4694),
            .I(N__4690));
    InMux I__523 (
            .O(N__4693),
            .I(N__4687));
    Odrv4 I__522 (
            .O(N__4690),
            .I(LIDE_BASE_4));
    LocalMux I__521 (
            .O(N__4687),
            .I(LIDE_BASE_4));
    InMux I__520 (
            .O(N__4682),
            .I(N__4678));
    InMux I__519 (
            .O(N__4681),
            .I(N__4675));
    LocalMux I__518 (
            .O(N__4678),
            .I(LIDE_BASE_3));
    LocalMux I__517 (
            .O(N__4675),
            .I(LIDE_BASE_3));
    InMux I__516 (
            .O(N__4670),
            .I(N__4667));
    LocalMux I__515 (
            .O(N__4667),
            .I(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_5 ));
    CascadeMux I__514 (
            .O(N__4664),
            .I(\U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_0Z0Z_3_cascade_ ));
    InMux I__513 (
            .O(N__4661),
            .I(N__4658));
    LocalMux I__512 (
            .O(N__4658),
            .I(\U409_ADDRESS_DECODE.HIROMZ0Z_0 ));
    CascadeMux I__511 (
            .O(N__4655),
            .I(N__4652));
    InMux I__510 (
            .O(N__4652),
            .I(N__4649));
    LocalMux I__509 (
            .O(N__4649),
            .I(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_0 ));
    CascadeMux I__508 (
            .O(N__4646),
            .I(\U409_AUTOCONFIG.N_99_cascade_ ));
    InMux I__507 (
            .O(N__4643),
            .I(N__4637));
    InMux I__506 (
            .O(N__4642),
            .I(N__4637));
    LocalMux I__505 (
            .O(N__4637),
            .I(LIDE_BASE_5));
    InMux I__504 (
            .O(N__4634),
            .I(N__4631));
    LocalMux I__503 (
            .O(N__4631),
            .I(N__4628));
    Sp12to4 I__502 (
            .O(N__4628),
            .I(N__4625));
    Span12Mux_v I__501 (
            .O(N__4625),
            .I(N__4622));
    Odrv12 I__500 (
            .O(N__4622),
            .I(D_in_4));
    InMux I__499 (
            .O(N__4619),
            .I(N__4616));
    LocalMux I__498 (
            .O(N__4616),
            .I(\U409_AUTOCONFIG.N_101 ));
    CascadeMux I__497 (
            .O(N__4613),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2_cascade_ ));
    CascadeMux I__496 (
            .O(N__4610),
            .I(N__4607));
    InMux I__495 (
            .O(N__4607),
            .I(N__4604));
    LocalMux I__494 (
            .O(N__4604),
            .I(N__4597));
    InMux I__493 (
            .O(N__4603),
            .I(N__4594));
    InMux I__492 (
            .O(N__4602),
            .I(N__4589));
    InMux I__491 (
            .O(N__4601),
            .I(N__4589));
    InMux I__490 (
            .O(N__4600),
            .I(N__4586));
    Odrv4 I__489 (
            .O(N__4597),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4 ));
    LocalMux I__488 (
            .O(N__4594),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4 ));
    LocalMux I__487 (
            .O(N__4589),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4 ));
    LocalMux I__486 (
            .O(N__4586),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4 ));
    InMux I__485 (
            .O(N__4577),
            .I(N__4574));
    LocalMux I__484 (
            .O(N__4574),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2 ));
    IoInMux I__483 (
            .O(N__4571),
            .I(N__4568));
    LocalMux I__482 (
            .O(N__4568),
            .I(N__4565));
    Span4Mux_s3_v I__481 (
            .O(N__4565),
            .I(N__4562));
    Span4Mux_h I__480 (
            .O(N__4562),
            .I(N__4559));
    Sp12to4 I__479 (
            .O(N__4559),
            .I(N__4556));
    Span12Mux_v I__478 (
            .O(N__4556),
            .I(N__4553));
    Span12Mux_h I__477 (
            .O(N__4553),
            .I(N__4550));
    Odrv12 I__476 (
            .O(N__4550),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn_i));
    InMux I__475 (
            .O(N__4547),
            .I(N__4544));
    LocalMux I__474 (
            .O(N__4544),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0Z0Z_0 ));
    InMux I__473 (
            .O(N__4541),
            .I(N__4538));
    LocalMux I__472 (
            .O(N__4538),
            .I(N__4535));
    Span4Mux_h I__471 (
            .O(N__4535),
            .I(N__4532));
    Odrv4 I__470 (
            .O(N__4532),
            .I(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7 ));
    InMux I__469 (
            .O(N__4529),
            .I(N__4526));
    LocalMux I__468 (
            .O(N__4526),
            .I(N__4523));
    Span4Mux_v I__467 (
            .O(N__4523),
            .I(N__4520));
    IoSpan4Mux I__466 (
            .O(N__4520),
            .I(N__4517));
    Odrv4 I__465 (
            .O(N__4517),
            .I(TT_c_1));
    InMux I__464 (
            .O(N__4514),
            .I(N__4511));
    LocalMux I__463 (
            .O(N__4511),
            .I(N__4508));
    Span4Mux_h I__462 (
            .O(N__4508),
            .I(N__4505));
    Span4Mux_v I__461 (
            .O(N__4505),
            .I(N__4502));
    Odrv4 I__460 (
            .O(N__4502),
            .I(TT_c_0));
    InMux I__459 (
            .O(N__4499),
            .I(N__4495));
    InMux I__458 (
            .O(N__4498),
            .I(N__4492));
    LocalMux I__457 (
            .O(N__4495),
            .I(LIDE_BASE_6));
    LocalMux I__456 (
            .O(N__4492),
            .I(LIDE_BASE_6));
    CascadeMux I__455 (
            .O(N__4487),
            .I(\U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_5_cascade_ ));
    InMux I__454 (
            .O(N__4484),
            .I(N__4480));
    InMux I__453 (
            .O(N__4483),
            .I(N__4477));
    LocalMux I__452 (
            .O(N__4480),
            .I(N__4472));
    LocalMux I__451 (
            .O(N__4477),
            .I(N__4472));
    Span4Mux_v I__450 (
            .O(N__4472),
            .I(N__4469));
    Span4Mux_h I__449 (
            .O(N__4469),
            .I(N__4466));
    Odrv4 I__448 (
            .O(N__4466),
            .I(A_c_25));
    CascadeMux I__447 (
            .O(N__4463),
            .I(N__4460));
    InMux I__446 (
            .O(N__4460),
            .I(N__4457));
    LocalMux I__445 (
            .O(N__4457),
            .I(N__4453));
    InMux I__444 (
            .O(N__4456),
            .I(N__4450));
    Span4Mux_h I__443 (
            .O(N__4453),
            .I(N__4445));
    LocalMux I__442 (
            .O(N__4450),
            .I(N__4445));
    Span4Mux_v I__441 (
            .O(N__4445),
            .I(N__4442));
    Span4Mux_h I__440 (
            .O(N__4442),
            .I(N__4439));
    Odrv4 I__439 (
            .O(N__4439),
            .I(A_c_24));
    InMux I__438 (
            .O(N__4436),
            .I(N__4433));
    LocalMux I__437 (
            .O(N__4433),
            .I(\U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4 ));
    InMux I__436 (
            .O(N__4430),
            .I(N__4424));
    InMux I__435 (
            .O(N__4429),
            .I(N__4424));
    LocalMux I__434 (
            .O(N__4424),
            .I(N__4421));
    Span4Mux_v I__433 (
            .O(N__4421),
            .I(N__4418));
    Span4Mux_h I__432 (
            .O(N__4418),
            .I(N__4415));
    Odrv4 I__431 (
            .O(N__4415),
            .I(A_c_29));
    InMux I__430 (
            .O(N__4412),
            .I(N__4406));
    InMux I__429 (
            .O(N__4411),
            .I(N__4406));
    LocalMux I__428 (
            .O(N__4406),
            .I(N__4403));
    Span4Mux_v I__427 (
            .O(N__4403),
            .I(N__4400));
    Span4Mux_h I__426 (
            .O(N__4400),
            .I(N__4397));
    Odrv4 I__425 (
            .O(N__4397),
            .I(A_c_31));
    CascadeMux I__424 (
            .O(N__4394),
            .I(N__4390));
    InMux I__423 (
            .O(N__4393),
            .I(N__4385));
    InMux I__422 (
            .O(N__4390),
            .I(N__4385));
    LocalMux I__421 (
            .O(N__4385),
            .I(N__4382));
    Span4Mux_v I__420 (
            .O(N__4382),
            .I(N__4379));
    Span4Mux_h I__419 (
            .O(N__4379),
            .I(N__4376));
    Odrv4 I__418 (
            .O(N__4376),
            .I(A_c_30));
    InMux I__417 (
            .O(N__4373),
            .I(N__4367));
    InMux I__416 (
            .O(N__4372),
            .I(N__4367));
    LocalMux I__415 (
            .O(N__4367),
            .I(N__4364));
    Span4Mux_v I__414 (
            .O(N__4364),
            .I(N__4361));
    Span4Mux_v I__413 (
            .O(N__4361),
            .I(N__4358));
    Sp12to4 I__412 (
            .O(N__4358),
            .I(N__4355));
    Odrv12 I__411 (
            .O(N__4355),
            .I(A_c_28));
    IoInMux I__410 (
            .O(N__4352),
            .I(N__4349));
    LocalMux I__409 (
            .O(N__4349),
            .I(N__4346));
    IoSpan4Mux I__408 (
            .O(N__4346),
            .I(N__4343));
    Span4Mux_s3_h I__407 (
            .O(N__4343),
            .I(N__4340));
    Sp12to4 I__406 (
            .O(N__4340),
            .I(N__4337));
    Span12Mux_s11_h I__405 (
            .O(N__4337),
            .I(N__4334));
    Span12Mux_h I__404 (
            .O(N__4334),
            .I(N__4331));
    Odrv12 I__403 (
            .O(N__4331),
            .I(U409_ADDRESS_DECODE_un1_RTC_ENn_i));
    InMux I__402 (
            .O(N__4328),
            .I(N__4325));
    LocalMux I__401 (
            .O(N__4325),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0 ));
    CascadeMux I__400 (
            .O(N__4322),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0_cascade_ ));
    CascadeMux I__399 (
            .O(N__4319),
            .I(\U409_ADDRESS_DECODE.HIROMZ0Z_0_cascade_ ));
    IoInMux I__398 (
            .O(N__4316),
            .I(N__4313));
    LocalMux I__397 (
            .O(N__4313),
            .I(N__4310));
    Span12Mux_s2_h I__396 (
            .O(N__4310),
            .I(N__4307));
    Span12Mux_v I__395 (
            .O(N__4307),
            .I(N__4304));
    Odrv12 I__394 (
            .O(N__4304),
            .I(SPIO_c));
    InMux I__393 (
            .O(N__4301),
            .I(N__4298));
    LocalMux I__392 (
            .O(N__4298),
            .I(N__4294));
    InMux I__391 (
            .O(N__4297),
            .I(N__4291));
    Span4Mux_v I__390 (
            .O(N__4294),
            .I(N__4286));
    LocalMux I__389 (
            .O(N__4291),
            .I(N__4286));
    Span4Mux_h I__388 (
            .O(N__4286),
            .I(N__4283));
    Span4Mux_v I__387 (
            .O(N__4283),
            .I(N__4280));
    Odrv4 I__386 (
            .O(N__4280),
            .I(A_c_26));
    CascadeMux I__385 (
            .O(N__4277),
            .I(N__4274));
    InMux I__384 (
            .O(N__4274),
            .I(N__4270));
    InMux I__383 (
            .O(N__4273),
            .I(N__4267));
    LocalMux I__382 (
            .O(N__4270),
            .I(N__4262));
    LocalMux I__381 (
            .O(N__4267),
            .I(N__4262));
    Span4Mux_v I__380 (
            .O(N__4262),
            .I(N__4259));
    Span4Mux_h I__379 (
            .O(N__4259),
            .I(N__4256));
    Odrv4 I__378 (
            .O(N__4256),
            .I(A_c_27));
    IoInMux I__377 (
            .O(N__4253),
            .I(N__4250));
    LocalMux I__376 (
            .O(N__4250),
            .I(N__4247));
    IoSpan4Mux I__375 (
            .O(N__4247),
            .I(N__4244));
    Sp12to4 I__374 (
            .O(N__4244),
            .I(N__4241));
    Span12Mux_s1_h I__373 (
            .O(N__4241),
            .I(N__4238));
    Span12Mux_v I__372 (
            .O(N__4238),
            .I(N__4235));
    Odrv12 I__371 (
            .O(N__4235),
            .I(PPIO_c));
    INV \INVU409_TRANSFER_ACK.LASTCLK_0C  (
            .O(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .I(N__9161));
    INV \INVU409_TRANSFER_ACK.LASTCLK_1C  (
            .O(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .I(N__9160));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .I(N__9155));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_1C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .I(N__9153));
    INV \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC  (
            .O(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .I(N__9158));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ),
            .I(N__9156));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ),
            .I(N__9154));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .I(N__9157));
    INV \INVU409_AUTOCONFIG.AC_TACK_nesrC  (
            .O(\INVU409_AUTOCONFIG.AC_TACK_nesrC_net ),
            .I(N__9821));
    INV \INVU409_AUTOCONFIG.LIDE_OUT_0C  (
            .O(\INVU409_AUTOCONFIG.LIDE_OUT_0C_net ),
            .I(N__9820));
    INV \INVU409_AUTOCONFIG.BRIDGE_OUT_0C  (
            .O(\INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ),
            .I(N__9824));
    INV \INVU409_AUTOCONFIG.CONFIGUREDC  (
            .O(\INVU409_AUTOCONFIG.CONFIGUREDC_net ),
            .I(N__9839));
    INV \INVU409_AUTOCONFIG.LIDE_OUT_2C  (
            .O(\INVU409_AUTOCONFIG.LIDE_OUT_2C_net ),
            .I(N__9823));
    INV \INVU409_AUTOCONFIG.STATE_0C  (
            .O(\INVU409_AUTOCONFIG.STATE_0C_net ),
            .I(N__9833));
    INV \INVU409_AUTOCONFIG.LIDE_BASE_7C  (
            .O(\INVU409_AUTOCONFIG.LIDE_BASE_7C_net ),
            .I(N__9838));
    INV \INVU409_AUTOCONFIG.BRIDGE_OUT_3C  (
            .O(\INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net ),
            .I(N__9830));
    INV \INVU409_AUTOCONFIG.PR_OUT_2C  (
            .O(\INVU409_AUTOCONFIG.PR_OUT_2C_net ),
            .I(N__9837));
    INV \INVU409_AUTOCONFIG.LIDE_BASE_1C  (
            .O(\INVU409_AUTOCONFIG.LIDE_BASE_1C_net ),
            .I(N__9842));
    INV \INVU409_AUTOCONFIG.LIDE_BASE_5C  (
            .O(\INVU409_AUTOCONFIG.LIDE_BASE_5C_net ),
            .I(N__9841));
    INV \INVU409_AUTOCONFIG.LIDE_BASE_3C  (
            .O(\INVU409_AUTOCONFIG.LIDE_BASE_3C_net ),
            .I(N__9846));
    defparam IN_MUX_bfv_17_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_5_0_));
    defparam IN_MUX_bfv_17_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_6_0_ (
            .carryinitin(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .carryinitout(bfn_17_6_0_));
    defparam IN_MUX_bfv_15_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_6_0_));
    defparam IN_MUX_bfv_15_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_7_0_ (
            .carryinitin(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .carryinitout(bfn_15_7_0_));
    defparam IN_MUX_bfv_12_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_6_0_));
    defparam IN_MUX_bfv_13_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_8_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__8465),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_1_17_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_1_17_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_1_17_4  (
            .in0(N__4483),
            .in1(N__4273),
            .in2(N__4463),
            .in3(N__4301),
            .lcout(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_5_LC_1_18_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_5_LC_1_18_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_5_LC_1_18_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_5_LC_1_18_1  (
            .in0(N__4297),
            .in1(N__4412),
            .in2(N__4277),
            .in3(N__4373),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_1_18_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_1_18_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_1_18_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_1_18_2  (
            .in0(N__4436),
            .in1(N__4393),
            .in2(N__4487),
            .in3(N__4430),
            .lcout(U409_ADDRESS_DECODE_Z2_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_4_LC_1_18_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_4_LC_1_18_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_4_LC_1_18_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_4_LC_1_18_5  (
            .in0(N__4484),
            .in1(N__9062),
            .in2(_gnd_net_),
            .in3(N__4456),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_1_18_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_1_18_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_1_18_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_1_18_7  (
            .in0(N__4429),
            .in1(N__4411),
            .in2(N__4394),
            .in3(N__4372),
            .lcout(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_5_7_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_5_7_3 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_5_7_3  (
            .in0(N__5126),
            .in1(N__4328),
            .in2(N__4610),
            .in3(N__5619),
            .lcout(U409_ADDRESS_DECODE_un1_RTC_ENn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_0_LC_5_8_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_0_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_0_LC_5_8_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_0_LC_5_8_4  (
            .in0(N__6267),
            .in1(N__5545),
            .in2(N__5192),
            .in3(N__5368),
            .lcout(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0 ),
            .ltout(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_5_8_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_5_8_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_5_8_5  (
            .in0(N__5127),
            .in1(N__4603),
            .in2(N__4322),
            .in3(N__5618),
            .lcout(U409_ADDRESS_DECODE_un1_RTC_ENn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.HIROM_0_LC_5_9_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.HIROM_0_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.HIROM_0_LC_5_9_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_ADDRESS_DECODE.HIROM_0_LC_5_9_5  (
            .in0(N__5536),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5617),
            .lcout(\U409_ADDRESS_DECODE.HIROMZ0Z_0 ),
            .ltout(\U409_ADDRESS_DECODE.HIROMZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_5_9_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_5_9_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_LC_5_9_6  (
            .in0(N__6266),
            .in1(N__7946),
            .in2(N__4319),
            .in3(N__4600),
            .lcout(CIA_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_5_9_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_5_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_5_9_7  (
            .in0(_gnd_net_),
            .in1(N__7710),
            .in2(_gnd_net_),
            .in3(N__6131),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0_LC_5_10_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0_LC_5_10_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0_LC_5_10_2  (
            .in0(N__6655),
            .in1(N__4547),
            .in2(N__5024),
            .in3(N__7314),
            .lcout(\U409_AUTOCONFIG.N_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_5_LC_5_10_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_5_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_5_LC_5_10_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_5_LC_5_10_7  (
            .in0(N__5186),
            .in1(N__5369),
            .in2(N__5137),
            .in3(N__4831),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0_0_LC_5_11_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0_0_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0_0_LC_5_11_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0_0_LC_5_11_1  (
            .in0(N__4928),
            .in1(N__4973),
            .in2(N__6450),
            .in3(N__4901),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_0_LC_5_11_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_0_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_0_LC_5_11_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_2_0_LC_5_11_5  (
            .in0(N__5030),
            .in1(N__4974),
            .in2(N__6451),
            .in3(N__4902),
            .lcout(\U409_AUTOCONFIG.LIDE_OUT_7_i_a3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_5_12_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_5_12_3 .LUT_INIT=16'b1010101000100010;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_5_12_3  (
            .in0(N__7313),
            .in1(N__4945),
            .in2(_gnd_net_),
            .in3(N__6632),
            .lcout(\U409_AUTOCONFIG.LIDE_OUT_7_i_a3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_5_20_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_5_20_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_5_20_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_5_20_7  (
            .in0(N__4541),
            .in1(N__4529),
            .in2(_gnd_net_),
            .in3(N__4514),
            .lcout(U409_ADDRESS_DECODE_AUTOVECTOR_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_BASE_3_LC_6_7_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_3_LC_6_7_0 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_3_LC_6_7_0 .LUT_INIT=16'b1110111111000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_3_LC_6_7_0  (
            .in0(N__5414),
            .in1(N__4709),
            .in2(N__5780),
            .in3(N__4682),
            .lcout(LIDE_BASE_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_3C_net ),
            .ce(),
            .sr(N__9751));
    defparam \U409_AUTOCONFIG.LIDE_BASE_6_LC_6_7_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_6_LC_6_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_6_LC_6_7_4 .LUT_INIT=16'b1110111111000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_6_LC_6_7_4  (
            .in0(N__5719),
            .in1(N__5450),
            .in2(N__5781),
            .in3(N__4499),
            .lcout(LIDE_BASE_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_3C_net ),
            .ce(),
            .sr(N__9751));
    defparam \U409_AUTOCONFIG.LIDE_BASE_4_LC_6_7_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_4_LC_6_7_5 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_4_LC_6_7_5 .LUT_INIT=16'b1110101011110000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_4_LC_6_7_5  (
            .in0(N__4619),
            .in1(N__5720),
            .in2(N__4700),
            .in3(N__5769),
            .lcout(LIDE_BASE_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_3C_net ),
            .ce(),
            .sr(N__9751));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_6_8_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_6_8_0 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_6_8_0  (
            .in0(N__4498),
            .in1(N__6269),
            .in2(N__5633),
            .in3(N__4642),
            .lcout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_5_LC_6_8_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_5_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_5_LC_6_8_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_RNO_0_5_LC_6_8_3  (
            .in0(N__5982),
            .in1(N__5718),
            .in2(N__5873),
            .in3(N__6902),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.N_99_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_BASE_5_LC_6_8_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_5_LC_6_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_5_LC_6_8_4 .LUT_INIT=16'b1111110110100000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_5_LC_6_8_4  (
            .in0(N__5749),
            .in1(N__5712),
            .in2(N__4646),
            .in3(N__4643),
            .lcout(LIDE_BASE_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_5C_net ),
            .ce(),
            .sr(N__9749));
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_4_LC_6_8_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_4_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_4_LC_6_8_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_RNO_0_4_LC_6_8_6  (
            .in0(N__4634),
            .in1(N__5981),
            .in2(N__6924),
            .in3(N__5711),
            .lcout(\U409_AUTOCONFIG.N_101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_2_LC_6_9_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_2_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_2_LC_6_9_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_2_LC_6_9_1  (
            .in0(N__5541),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6268),
            .lcout(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2 ),
            .ltout(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_9_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_9_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_9_2  (
            .in0(N__7947),
            .in1(N__4601),
            .in2(N__4613),
            .in3(N__5624),
            .lcout(U409_ADDRESS_DECODE_un1_REGSPACEn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_9_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_9_5 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_9_5  (
            .in0(N__4602),
            .in1(N__4577),
            .in2(N__5632),
            .in3(N__7948),
            .lcout(U409_ADDRESS_DECODE_un1_REGSPACEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PORTSIZE_1_LC_6_9_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_1_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_1_LC_6_9_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_ADDRESS_DECODE.PORTSIZE_1_LC_6_9_6  (
            .in0(N__7876),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6879),
            .lcout(\U409_ADDRESS_DECODE.PORTSIZEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNIU6QK1_1_LC_6_9_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNIU6QK1_1_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNIU6QK1_1_LC_6_9_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNIU6QK1_1_LC_6_9_7  (
            .in0(N__4991),
            .in1(N__6050),
            .in2(N__4844),
            .in3(N__7099),
            .lcout(\U409_AUTOCONFIG.un1_STATE_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_LC_6_10_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_LC_6_10_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_LC_6_10_0  (
            .in0(N__5370),
            .in1(N__4670),
            .in2(N__4655),
            .in3(N__5603),
            .lcout(AUTOCONFIG_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_5_LC_6_10_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_5_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_5_LC_6_10_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_5_LC_6_10_3  (
            .in0(N__7703),
            .in1(N__5187),
            .in2(N__4832),
            .in3(N__5125),
            .lcout(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_0_3_LC_6_10_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_0_3_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_0_3_LC_6_10_4 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_0_3_LC_6_10_4  (
            .in0(N__6513),
            .in1(N__6456),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_0Z0Z_3 ),
            .ltout(\U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_RNO_0_2_LC_6_10_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_RNO_0_2_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_RNO_0_2_LC_6_10_5 .LUT_INIT=16'b1111111101110101;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_RNO_0_2_LC_6_10_5  (
            .in0(N__9058),
            .in1(N__7320),
            .in2(N__4664),
            .in3(N__7477),
            .lcout(\U409_AUTOCONFIG.PR_OUT_cnst_i_i_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.HIROM_LC_6_10_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.HIROM_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.HIROM_LC_6_10_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.HIROM_LC_6_10_6  (
            .in0(N__5371),
            .in1(N__4661),
            .in2(N__6135),
            .in3(N__6244),
            .lcout(U409_ADDRESS_DECODE_HIROM),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_0_LC_6_10_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_0_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_0_LC_6_10_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_0_LC_6_10_7  (
            .in0(N__5520),
            .in1(N__6238),
            .in2(_gnd_net_),
            .in3(N__6117),
            .lcout(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_0_a3_3_LC_6_11_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_0_a3_3_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_0_a3_3_LC_6_11_0 .LUT_INIT=16'b1000000000001000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_7_0_a3_3_LC_6_11_0  (
            .in0(N__7315),
            .in1(N__6495),
            .in2(N__6463),
            .in3(N__6656),
            .lcout(\U409_AUTOCONFIG.N_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_2_LC_6_11_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_2_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_2_LC_6_11_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_2_LC_6_11_3  (
            .in0(N__4857),
            .in1(N__4976),
            .in2(_gnd_net_),
            .in3(N__7316),
            .lcout(\U409_AUTOCONFIG.N_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_A_13_0_a2_LC_6_11_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_A_13_0_a2_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_A_13_0_a2_LC_6_11_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_AUTOCONFIG.un1_A_13_0_a2_LC_6_11_4  (
            .in0(N__4977),
            .in1(N__4858),
            .in2(N__7337),
            .in3(N__4904),
            .lcout(\U409_AUTOCONFIG.un1_A_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_2_LC_6_11_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_2_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_2_LC_6_11_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_2_LC_6_11_5  (
            .in0(N__4938),
            .in1(N__5028),
            .in2(N__6673),
            .in3(N__6455),
            .lcout(\U409_AUTOCONFIG.N_121 ),
            .ltout(\U409_AUTOCONFIG.N_121_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_3_LC_6_11_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_3_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_3_LC_6_11_6 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_3_LC_6_11_6  (
            .in0(N__4975),
            .in1(_gnd_net_),
            .in2(N__5033),
            .in3(N__4903),
            .lcout(\U409_AUTOCONFIG.N_129 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_0_3_LC_6_12_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_0_3_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_0_3_LC_6_12_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_0_3_LC_6_12_4  (
            .in0(N__5029),
            .in1(N__4990),
            .in2(N__4946),
            .in3(N__4900),
            .lcout(\U409_AUTOCONFIG.N_110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_0_3_LC_6_12_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_0_3_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_0_3_LC_6_12_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_0_3_LC_6_12_7  (
            .in0(N__4899),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4859),
            .lcout(\U409_AUTOCONFIG.N_123 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CS0_LC_7_2_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CS0_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CS0_LC_7_2_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_ADDRESS_DECODE.CS0_LC_7_2_5  (
            .in0(N__4814),
            .in1(N__4777),
            .in2(N__8383),
            .in3(N__8451),
            .lcout(\U409_ADDRESS_DECODE.CSZ0Z0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CS1_LC_7_3_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CS1_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CS1_LC_7_3_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U409_ADDRESS_DECODE.CS1_LC_7_3_2  (
            .in0(N__4815),
            .in1(N__8379),
            .in2(N__8455),
            .in3(N__4778),
            .lcout(\U409_ADDRESS_DECODE.CSZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.D_1_i_LC_7_6_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.D_1_i_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.D_1_i_LC_7_6_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_ADDRESS_DECODE.D_1_i_LC_7_6_1  (
            .in0(N__5985),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6936),
            .lcout(D_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_3_LC_7_6_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_3_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_3_LC_7_6_4 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_RNO_0_3_LC_7_6_4  (
            .in0(N__6937),
            .in1(N__5290),
            .in2(N__5999),
            .in3(N__5408),
            .lcout(\U409_AUTOCONFIG.N_103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_7_7_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_7_7_0 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_7_7_0  (
            .in0(N__5546),
            .in1(N__4693),
            .in2(N__5359),
            .in3(N__4681),
            .lcout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_BASE_1_LC_7_7_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_1_LC_7_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_1_LC_7_7_4 .LUT_INIT=16'b1110111111000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_1_LC_7_7_4  (
            .in0(N__5409),
            .in1(N__5840),
            .in2(N__5782),
            .in3(N__5087),
            .lcout(LIDE_BASE_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_1C_net ),
            .ce(),
            .sr(N__9750));
    defparam \U409_AUTOCONFIG.LIDE_BASE_2_LC_7_7_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_2_LC_7_7_6 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_2_LC_7_7_6 .LUT_INIT=16'b1110111111000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_2_LC_7_7_6  (
            .in0(N__5410),
            .in1(N__5420),
            .in2(N__5783),
            .in3(N__5150),
            .lcout(LIDE_BASE_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_1C_net ),
            .ce(),
            .sr(N__9750));
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_7_LC_7_7_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_7_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_7_LC_7_7_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_RNO_0_7_LC_7_7_7  (
            .in0(N__5294),
            .in1(N__5984),
            .in2(N__6939),
            .in3(N__5709),
            .lcout(\U409_AUTOCONFIG.N_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_LC_7_8_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_LC_7_8_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_ADDRESS_DECODE.PORTSIZE_0_LC_7_8_1  (
            .in0(N__8047),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7138),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.PORTSIZEZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNIOGLSO_LC_7_8_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNIOGLSO_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNIOGLSO_LC_7_8_2 .LUT_INIT=16'b1011111100111111;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_EN_RNIOGLSO_LC_7_8_2  (
            .in0(N__5044),
            .in1(N__5264),
            .in2(N__5258),
            .in3(N__5058),
            .lcout(PORTSIZE_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.LV_SPACE_LC_7_8_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.LV_SPACE_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.LV_SPACE_LC_7_8_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.LV_SPACE_LC_7_8_3  (
            .in0(N__5060),
            .in1(N__7137),
            .in2(N__6935),
            .in3(N__7117),
            .lcout(BUFENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNITH4D5_LC_7_8_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNITH4D5_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNITH4D5_LC_7_8_4 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_EN_RNITH4D5_LC_7_8_4  (
            .in0(N__5045),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5059),
            .lcout(U409_ADDRESS_DECODE_un1_ATA_ENn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_1_LC_7_8_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_1_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_1_LC_7_8_5 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_1_LC_7_8_5  (
            .in0(N__5191),
            .in1(N__5149),
            .in2(N__5138),
            .in3(N__5086),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_LC_7_8_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_LC_7_8_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_LC_7_8_6  (
            .in0(N__5075),
            .in1(N__5789),
            .in2(N__5069),
            .in3(N__5066),
            .lcout(\U409_ADDRESS_DECODE.ATA_SPACEZ0 ),
            .ltout(\U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_EN_LC_7_8_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_EN_LC_7_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_ADDRESS_DECODE.ATA_EN_LC_7_8_7 .LUT_INIT=16'b1111111101010000;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_EN_LC_7_8_7  (
            .in0(N__5983),
            .in1(_gnd_net_),
            .in2(N__5048),
            .in3(N__5043),
            .lcout(\U409_ADDRESS_DECODE.ATA_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9840),
            .ce(),
            .sr(N__9748));
    defparam \U409_AUTOCONFIG.PR_OUT_2_LC_7_9_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_2_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.PR_OUT_2_LC_7_9_3 .LUT_INIT=16'b0000000011011111;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_2_LC_7_9_3  (
            .in0(N__6712),
            .in1(N__6672),
            .in2(N__6464),
            .in3(N__5384),
            .lcout(\U409_AUTOCONFIG.PR_OUTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.PR_OUT_2C_net ),
            .ce(N__7407),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_1_LC_7_10_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_1_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_1_LC_7_10_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_1_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(N__5623),
            .in2(_gnd_net_),
            .in3(N__7704),
            .lcout(\U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_1 ),
            .ltout(\U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_7_10_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_7_10_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_7_10_3  (
            .in0(N__6247),
            .in1(N__6184),
            .in2(N__5378),
            .in3(N__6138),
            .lcout(U409_ADDRESS_DECODE_un1_RAMSPACEn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.LOWROM_3_LC_7_10_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.LOWROM_3_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.LOWROM_3_LC_7_10_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U409_ADDRESS_DECODE.LOWROM_3_LC_7_10_4  (
            .in0(N__6137),
            .in1(N__6183),
            .in2(N__5375),
            .in3(N__6246),
            .lcout(\U409_ADDRESS_DECODE.LOWROMZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_4_0_LC_7_10_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_4_0_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_4_0_LC_7_10_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_4_0_LC_7_10_5  (
            .in0(N__6245),
            .in1(N__6136),
            .in2(N__5631),
            .in3(N__5540),
            .lcout(\U409_ADDRESS_DECODE.AUTOVECTOR_4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_1_LC_7_10_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_1_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_1_LC_7_10_7 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_1_LC_7_10_7  (
            .in0(N__6514),
            .in1(N__6457),
            .in2(_gnd_net_),
            .in3(N__6671),
            .lcout(\U409_AUTOCONFIG.N_131 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_7_11_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_7_11_0 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_7_11_0 .LUT_INIT=16'b0000000010001010;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_7_11_0  (
            .in0(N__9045),
            .in1(N__7322),
            .in2(N__6553),
            .in3(N__5314),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net ),
            .ce(N__7412),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_3_LC_7_11_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_3_LC_7_11_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_3_LC_7_11_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_3_LC_7_11_1  (
            .in0(N__5315),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9046),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net ),
            .ce(N__7412),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIBHMP_3_LC_7_11_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIBHMP_3_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIBHMP_3_LC_7_11_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNIBHMP_3_LC_7_11_2  (
            .in0(N__5306),
            .in1(N__5300),
            .in2(_gnd_net_),
            .in3(N__6995),
            .lcout(\U409_AUTOCONFIG.LIDE_OUT_RNIBHMPZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_3_LC_7_12_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_3_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_3_LC_7_12_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_3_LC_7_12_4  (
            .in0(N__6496),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7321),
            .lcout(\U409_AUTOCONFIG.N_116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.LOWROM_LC_7_12_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.LOWROM_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.LOWROM_LC_7_12_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_ADDRESS_DECODE.LOWROM_LC_7_12_7  (
            .in0(N__5642),
            .in1(N__5583),
            .in2(_gnd_net_),
            .in3(N__5519),
            .lcout(U409_ADDRESS_DECODE_LOWROM),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_RNIVV912_2_LC_8_6_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_RNIVV912_2_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_RNIVV912_2_LC_8_6_7 .LUT_INIT=16'b1011101110111000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_RNIVV912_2_LC_8_6_7  (
            .in0(N__6566),
            .in1(N__7040),
            .in2(N__5474),
            .in3(N__6852),
            .lcout(D_OUT_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_6_LC_8_7_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_6_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_6_LC_8_7_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_RNO_0_6_LC_8_7_0  (
            .in0(N__5435),
            .in1(N__6011),
            .in2(N__6941),
            .in3(N__5697),
            .lcout(\U409_AUTOCONFIG.N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNIF4QU_1_LC_8_7_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNIF4QU_1_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNIF4QU_1_LC_8_7_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNIF4QU_1_LC_8_7_2  (
            .in0(_gnd_net_),
            .in1(N__6049),
            .in2(_gnd_net_),
            .in3(N__7095),
            .lcout(\U409_AUTOCONFIG.STATE_d_2 ),
            .ltout(\U409_AUTOCONFIG.STATE_d_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2_LC_8_7_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2_LC_8_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2_LC_8_7_3  (
            .in0(N__5668),
            .in1(N__6984),
            .in2(N__5438),
            .in3(N__5825),
            .lcout(\U409_AUTOCONFIG.CONFIGENn_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_2_LC_8_7_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_2_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_2_LC_8_7_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_RNO_0_2_LC_8_7_4  (
            .in0(N__5434),
            .in1(N__6010),
            .in2(N__6940),
            .in3(N__5407),
            .lcout(\U409_AUTOCONFIG.N_105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIH4AI_LC_8_7_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIH4AI_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIH4AI_LC_8_7_5 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNIH4AI_LC_8_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5672),
            .in3(N__6985),
            .lcout(\U409_AUTOCONFIG.N_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI0CVL_0_LC_8_7_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI0CVL_0_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI0CVL_0_LC_8_7_6 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNI0CVL_0_LC_8_7_6  (
            .in0(N__7339),
            .in1(N__5667),
            .in2(_gnd_net_),
            .in3(N__6983),
            .lcout(\U409_AUTOCONFIG.N_49 ),
            .ltout(\U409_AUTOCONFIG.N_49_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_1_LC_8_7_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_1_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_1_LC_8_7_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_RNO_0_1_LC_8_7_7  (
            .in0(N__6009),
            .in1(N__5860),
            .in2(N__5843),
            .in3(N__6928),
            .lcout(\U409_AUTOCONFIG.N_107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI0CVL_LC_8_8_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI0CVL_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI0CVL_LC_8_8_0 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNI0CVL_LC_8_8_0  (
            .in0(N__7338),
            .in1(N__5665),
            .in2(_gnd_net_),
            .in3(N__6981),
            .lcout(\U409_AUTOCONFIG.N_48 ),
            .ltout(\U409_AUTOCONFIG.N_48_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_BASE_7_LC_8_8_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_7_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_7_LC_8_8_1 .LUT_INIT=16'b1111110110001000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_7_LC_8_8_1  (
            .in0(N__5779),
            .in1(N__5834),
            .in2(N__5828),
            .in3(N__5798),
            .lcout(LIDE_BASE_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_7C_net ),
            .ce(),
            .sr(N__9746));
    defparam \U409_AUTOCONFIG.BRIDGE_CONF_LC_8_8_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_CONF_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_CONF_LC_8_8_6 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_CONF_LC_8_8_6  (
            .in0(N__5821),
            .in1(N__5804),
            .in2(_gnd_net_),
            .in3(N__6982),
            .lcout(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_7C_net ),
            .ce(),
            .sr(N__9746));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_4_LC_8_8_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_4_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_4_LC_8_8_7 .LUT_INIT=16'b1000001000000000;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_4_LC_8_8_7  (
            .in0(N__7690),
            .in1(N__5797),
            .in2(N__6143),
            .in3(N__6842),
            .lcout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_0_LC_8_9_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_0_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.STATE_0_LC_8_9_2 .LUT_INIT=16'b0010001100100010;
    LogicCell40 \U409_AUTOCONFIG.STATE_0_LC_8_9_2  (
            .in0(N__6048),
            .in1(N__7094),
            .in2(N__5912),
            .in3(N__6809),
            .lcout(\U409_AUTOCONFIG.STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.STATE_0C_net ),
            .ce(),
            .sr(N__9743));
    defparam \U409_AUTOCONFIG.STATE_1_LC_8_9_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_1_LC_8_9_4 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.STATE_1_LC_8_9_4 .LUT_INIT=16'b0001000111001100;
    LogicCell40 \U409_AUTOCONFIG.STATE_1_LC_8_9_4  (
            .in0(N__6001),
            .in1(N__6047),
            .in2(_gnd_net_),
            .in3(N__7093),
            .lcout(\U409_AUTOCONFIG.STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.STATE_0C_net ),
            .ce(),
            .sr(N__9743));
    defparam \U409_AUTOCONFIG.LIDE_CONF_LC_8_9_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_LC_8_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_LC_8_9_6 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_LC_8_9_6  (
            .in0(N__5762),
            .in1(N__5666),
            .in2(_gnd_net_),
            .in3(N__5710),
            .lcout(\U409_AUTOCONFIG.LIDE_CONFZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.STATE_0C_net ),
            .ce(),
            .sr(N__9743));
    defparam \U409_AUTOCONFIG.STATE_ns_1_0__m4_LC_8_10_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_ns_1_0__m4_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_ns_1_0__m4_LC_8_10_0 .LUT_INIT=16'b0101010100001010;
    LogicCell40 \U409_AUTOCONFIG.STATE_ns_1_0__m4_LC_8_10_0  (
            .in0(N__7088),
            .in1(_gnd_net_),
            .in2(N__6000),
            .in3(N__6042),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.STATE_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_TACK_nesr_RNO_LC_8_10_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_TACK_nesr_RNO_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.AC_TACK_nesr_RNO_LC_8_10_1 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \U409_AUTOCONFIG.AC_TACK_nesr_RNO_LC_8_10_1  (
            .in0(N__9755),
            .in1(_gnd_net_),
            .in2(N__6272),
            .in3(_gnd_net_),
            .lcout(\U409_AUTOCONFIG.STATE_ns_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_8_10_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_8_10_2 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_8_10_2  (
            .in0(N__6253),
            .in1(N__6194),
            .in2(N__6185),
            .in3(N__6139),
            .lcout(U409_ADDRESS_DECODE_un1_RAMSPACEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNIBIND1_1_LC_8_10_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNIBIND1_1_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNIBIND1_1_LC_8_10_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNIBIND1_1_LC_8_10_3  (
            .in0(N__6043),
            .in1(N__5989),
            .in2(_gnd_net_),
            .in3(N__7089),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_a3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_START_RNI10V92_LC_8_10_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_START_RNI10V92_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.AC_START_RNI10V92_LC_8_10_4 .LUT_INIT=16'b0111001100110011;
    LogicCell40 \U409_AUTOCONFIG.AC_START_RNI10V92_LC_8_10_4  (
            .in0(N__5905),
            .in1(N__9035),
            .in2(N__5879),
            .in3(N__6808),
            .lcout(\U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_RNO_0_1_LC_8_10_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_RNO_0_1_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_RNO_0_1_LC_8_10_5 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_RNO_0_1_LC_8_10_5  (
            .in0(_gnd_net_),
            .in1(N__6449),
            .in2(N__6524),
            .in3(N__7325),
            .lcout(\U409_AUTOCONFIG.N_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_8_10_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_8_10_6 .LUT_INIT=16'b0100100000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_8_10_6  (
            .in0(N__6684),
            .in1(N__6520),
            .in2(N__6462),
            .in3(N__7324),
            .lcout(\U409_AUTOCONFIG.N_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_8_11_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_8_11_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(N__6445),
            .in2(_gnd_net_),
            .in3(N__6670),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.N_227_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_2_LC_8_11_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_2_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_2_LC_8_11_1 .LUT_INIT=16'b0000000001001100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_2_LC_8_11_1  (
            .in0(N__6705),
            .in1(N__9041),
            .in2(N__5876),
            .in3(N__6533),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_2C_net ),
            .ce(N__7406),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_8_11_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_8_11_3 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_8_11_3 .LUT_INIT=16'b0000000011000100;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_8_11_3  (
            .in0(N__6704),
            .in1(N__9040),
            .in2(N__6461),
            .in3(N__6532),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_2C_net ),
            .ce(N__7406),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNI9FMP_2_LC_8_11_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNI9FMP_2_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNI9FMP_2_LC_8_11_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNI9FMP_2_LC_8_11_4  (
            .in0(N__6578),
            .in1(N__6994),
            .in2(_gnd_net_),
            .in3(N__6572),
            .lcout(\U409_AUTOCONFIG.LIDE_OUT_RNI9FMPZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_0_LC_8_12_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_0_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_0_LC_8_12_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_0_LC_8_12_1  (
            .in0(N__6675),
            .in1(N__6512),
            .in2(_gnd_net_),
            .in3(N__6411),
            .lcout(\U409_AUTOCONFIG.N_133 ),
            .ltout(\U409_AUTOCONFIG.N_133_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_0_a2_2_LC_8_12_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_0_a2_2_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_7_0_a2_2_LC_8_12_2 .LUT_INIT=16'b0000000011111010;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_7_0_a2_2_LC_8_12_2  (
            .in0(N__6557),
            .in1(_gnd_net_),
            .in2(N__6536),
            .in3(N__7323),
            .lcout(\U409_AUTOCONFIG.N_127 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_1_LC_8_12_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_1_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_1_LC_8_12_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_1_LC_8_12_7  (
            .in0(N__6674),
            .in1(N__6511),
            .in2(_gnd_net_),
            .in3(N__6410),
            .lcout(\U409_AUTOCONFIG.N_126 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_RNISS912_1_LC_9_6_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_RNISS912_1_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_RNISS912_1_LC_9_6_1 .LUT_INIT=16'b1011101110111000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_RNISS912_1_LC_9_6_1  (
            .in0(N__7004),
            .in1(N__7044),
            .in2(N__6731),
            .in3(N__6848),
            .lcout(D_OUT_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_RNI23A12_3_LC_9_6_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_RNI23A12_3_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_RNI23A12_3_LC_9_6_2 .LUT_INIT=16'b1100111111001010;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_RNI23A12_3_LC_9_6_2  (
            .in0(N__6847),
            .in1(N__6341),
            .in2(N__7046),
            .in3(N__6761),
            .lcout(D_OUT_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.CONFIGURED_LC_9_7_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.CONFIGURED_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.CONFIGURED_LC_9_7_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U409_AUTOCONFIG.CONFIGURED_LC_9_7_3  (
            .in0(N__6308),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6846),
            .lcout(CONFIGURED),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.CONFIGUREDC_net ),
            .ce(),
            .sr(N__9747));
    defparam \U409_AUTOCONFIG.CONFIGENn_LC_9_7_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.CONFIGENn_LC_9_7_6 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.CONFIGENn_LC_9_7_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U409_AUTOCONFIG.CONFIGENn_LC_9_7_6  (
            .in0(_gnd_net_),
            .in1(N__6283),
            .in2(_gnd_net_),
            .in3(N__6307),
            .lcout(CONFIGENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.CONFIGUREDC_net ),
            .ce(),
            .sr(N__9747));
    defparam \U409_AUTOCONFIG.PR_OUT_RNIPP912_0_LC_9_8_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_RNIPP912_0_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_RNIPP912_0_LC_9_8_0 .LUT_INIT=16'b1011101110111000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_RNIPP912_0_LC_9_8_0  (
            .in0(N__6947),
            .in1(N__7045),
            .in2(N__6854),
            .in3(N__7454),
            .lcout(D_OUT_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNI7DMP_1_LC_9_8_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNI7DMP_1_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNI7DMP_1_LC_9_8_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNI7DMP_1_LC_9_8_6  (
            .in0(N__6987),
            .in1(N__6782),
            .in2(_gnd_net_),
            .in3(N__6587),
            .lcout(\U409_AUTOCONFIG.LIDE_OUT_RNI7DMPZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNI5BMP_0_LC_9_8_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNI5BMP_0_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNI5BMP_0_LC_9_8_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNI5BMP_0_LC_9_8_7  (
            .in0(N__7421),
            .in1(N__6797),
            .in2(_gnd_net_),
            .in3(N__6986),
            .lcout(\U409_AUTOCONFIG.LIDE_OUT_RNI5BMPZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_START_LC_9_9_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_START_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.AC_START_LC_9_9_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_AUTOCONFIG.AC_START_LC_9_9_2  (
            .in0(N__6938),
            .in1(N__7987),
            .in2(_gnd_net_),
            .in3(N__6853),
            .lcout(\U409_AUTOCONFIG.AC_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9831),
            .ce(),
            .sr(N__9736));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_9_10_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_9_10_0 .LUT_INIT=16'b0100010000000100;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_9_10_0  (
            .in0(N__7465),
            .in1(N__9025),
            .in2(N__6752),
            .in3(N__7333),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ),
            .ce(N__7390),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_1_LC_9_10_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_1_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_1_LC_9_10_1 .LUT_INIT=16'b0000000010100010;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_1_LC_9_10_1  (
            .in0(N__9027),
            .in1(N__7183),
            .in2(N__7340),
            .in3(N__6788),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ),
            .ce(N__7390),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_3_LC_9_10_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_3_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.PR_OUT_3_LC_9_10_2 .LUT_INIT=16'b0000010001000100;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_3_LC_9_10_2  (
            .in0(N__6719),
            .in1(N__9034),
            .in2(N__6773),
            .in3(N__6686),
            .lcout(\U409_AUTOCONFIG.PR_OUTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ),
            .ce(N__7390),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_1_LC_9_10_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_1_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.PR_OUT_1_LC_9_10_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_1_LC_9_10_5  (
            .in0(N__7487),
            .in1(N__6751),
            .in2(N__9048),
            .in3(N__6737),
            .lcout(\U409_AUTOCONFIG.PR_OUTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ),
            .ce(N__7390),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_9_10_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_9_10_6 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_9_10_6 .LUT_INIT=16'b0000110100000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_9_10_6  (
            .in0(N__6718),
            .in1(N__6685),
            .in2(N__7184),
            .in3(N__9026),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ),
            .ce(N__7390),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_0_LC_9_10_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_0_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.PR_OUT_0_LC_9_10_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_0_LC_9_10_7  (
            .in0(N__7486),
            .in1(N__7466),
            .in2(N__9047),
            .in3(N__7355),
            .lcout(\U409_AUTOCONFIG.PR_OUTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ),
            .ce(N__7390),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_0_LC_9_11_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_0_LC_9_11_5 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_0_LC_9_11_5 .LUT_INIT=16'b0001001100000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_0_LC_9_11_5  (
            .in0(N__7445),
            .in1(N__7163),
            .in2(N__7436),
            .in3(N__9036),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_0C_net ),
            .ce(N__7411),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_9_12_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_9_12_5 .LUT_INIT=16'b0010111100100010;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_9_12_5  (
            .in0(N__7351),
            .in1(N__7332),
            .in2(N__7211),
            .in3(N__7174),
            .lcout(\U409_AUTOCONFIG.LIDE_OUT_7_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_10_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_10_9_3 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_10_9_3  (
            .in0(N__7157),
            .in1(N__7142),
            .in2(N__7124),
            .in3(N__9007),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_TACK_nesr_LC_10_10_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_TACK_nesr_LC_10_10_0 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.AC_TACK_nesr_LC_10_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_AUTOCONFIG.AC_TACK_nesr_LC_10_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7100),
            .lcout(AC_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.AC_TACK_nesrC_net ),
            .ce(N__7055),
            .sr(N__9733));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIQ2ND1_7_LC_11_6_0 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIQ2ND1_7_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIQ2ND1_7_LC_11_6_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIQ2ND1_7_LC_11_6_0  (
            .in0(N__8763),
            .in1(N__8832),
            .in2(N__8665),
            .in3(N__8734),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_11_6_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_11_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_11_6_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_0_LC_11_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8802),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11149),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_11_6_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_11_6_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_11_6_6  (
            .in0(N__8602),
            .in1(N__8632),
            .in2(N__8701),
            .in3(N__8801),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_2_0 ),
            .ltout(\U409_CIA.CIA_CLK_COUNT11_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_11_6_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_11_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_11_6_7 .LUT_INIT=16'b0001001101001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_5_LC_11_6_7  (
            .in0(N__7786),
            .in1(N__8695),
            .in2(N__7508),
            .in3(N__7811),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11149),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_8_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_8_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_8_0 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_8_0  (
            .in0(N__8314),
            .in1(N__7862),
            .in2(N__7850),
            .in3(N__8269),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__8086));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_8_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_8_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_8_1  (
            .in0(N__7860),
            .in1(N__8268),
            .in2(_gnd_net_),
            .in3(N__8313),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_8_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_8_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_8_2 .LUT_INIT=16'b0000001100110000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(N__7843),
            .in2(N__7505),
            .in3(N__8230),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__8086));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_8_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_8_3 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_8_3 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_8_3  (
            .in0(N__8229),
            .in1(N__8246),
            .in2(N__7502),
            .in3(N__7848),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__8086));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_11_8_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_11_8_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_11_8_4  (
            .in0(N__8124),
            .in1(N__8185),
            .in2(_gnd_net_),
            .in3(N__8207),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_8_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_8_5 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_8_5 .LUT_INIT=16'b0000000000111100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(N__8291),
            .in2(N__7493),
            .in3(N__7847),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__8086));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_5_LC_11_8_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_5_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_5_LC_11_8_6 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_5_LC_11_8_6  (
            .in0(N__8008),
            .in1(N__9869),
            .in2(N__8156),
            .in3(N__8139),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_8_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_8_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_8_7 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_8_7  (
            .in0(N__7861),
            .in1(_gnd_net_),
            .in2(N__7490),
            .in3(N__8315),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__8086));
    defparam \U409_TRANSFER_ACK.TACK_OUT_RNO_0_LC_11_9_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUT_RNO_0_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_OUT_RNO_0_LC_11_9_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUT_RNO_0_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__10062),
            .in2(_gnd_net_),
            .in3(N__9185),
            .lcout(\U409_TRANSFER_ACK.TACK_EN8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_RNO_0_LC_11_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_RNO_0_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_EN_RNO_0_LC_11_9_6 .LUT_INIT=16'b0000000011111010;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_RNO_0_LC_11_9_6  (
            .in0(N__10063),
            .in1(_gnd_net_),
            .in2(N__9193),
            .in3(N__7751),
            .lcout(\U409_TRANSFER_ACK.TACK_STATE_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUT_LC_11_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUT_LC_11_10_0 .SEQ_MODE=4'b1001;
    defparam \U409_TRANSFER_ACK.TACK_OUT_LC_11_10_0 .LUT_INIT=16'b1101110111001000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUT_LC_11_10_0  (
            .in0(N__7732),
            .in1(N__7586),
            .in2(N__7769),
            .in3(N__7752),
            .lcout(TACK_OUT),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9818),
            .ce(),
            .sr(N__9732));
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_11_10_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_11_10_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_11_10_1 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_LC_11_10_1  (
            .in0(N__9078),
            .in1(N__7731),
            .in2(_gnd_net_),
            .in3(N__7760),
            .lcout(TACK_EN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9818),
            .ce(),
            .sr(N__9732));
    defparam \U409_TRANSFER_ACK.TACK_STATE_0_LC_11_10_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_STATE_0_LC_11_10_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_STATE_0_LC_11_10_2 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \U409_TRANSFER_ACK.TACK_STATE_0_LC_11_10_2  (
            .in0(N__7754),
            .in1(N__10067),
            .in2(N__7733),
            .in3(N__9194),
            .lcout(\U409_TRANSFER_ACK.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9818),
            .ce(),
            .sr(N__9732));
    defparam \U409_TRANSFER_ACK.TACK_STATE_1_LC_11_10_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_STATE_1_LC_11_10_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_STATE_1_LC_11_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_STATE_1_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7753),
            .lcout(\U409_TRANSFER_ACK.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9818),
            .ce(),
            .sr(N__9732));
    defparam \U409_TRANSFER_ACK.ROM_TACK_STATE5_LC_11_11_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_STATE5_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_STATE5_LC_11_11_5 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_STATE5_LC_11_11_5  (
            .in0(N__7718),
            .in1(N__7565),
            .in2(N__7646),
            .in3(N__8007),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUT_RNIU3I06_LC_11_12_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUT_RNIU3I06_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_OUT_RNIU3I06_LC_11_12_5 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUT_RNIU3I06_LC_11_12_5  (
            .in0(N__7717),
            .in1(N__7645),
            .in2(N__7605),
            .in3(N__7561),
            .lcout(U409_TRANSFER_ACK_un1_TACK_OUT_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_2.C_ON=1'b0;
    defparam GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_2.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9871),
            .lcout(GB_BUFFER_CLK40_IN_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_6_0 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(N__8730),
            .in2(N__8806),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_6_0_),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_12_6_1 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_12_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_2_LC_12_6_1  (
            .in0(_gnd_net_),
            .in1(N__8600),
            .in2(_gnd_net_),
            .in3(N__7820),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .clk(N__11148),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_12_6_2 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_12_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_12_6_2  (
            .in0(_gnd_net_),
            .in1(N__8629),
            .in2(_gnd_net_),
            .in3(N__7817),
            .lcout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_12_6_3 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_12_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_12_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_4_LC_12_6_3  (
            .in0(_gnd_net_),
            .in1(N__8657),
            .in2(_gnd_net_),
            .in3(N__7814),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .clk(N__11148),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_LUT4_0_LC_12_6_4 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_LUT4_0_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_LUT4_0_LC_12_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_LUT4_0_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(N__8696),
            .in2(_gnd_net_),
            .in3(N__7805),
            .lcout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_12_6_5 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_12_6_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_12_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_6_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(N__8833),
            .in2(_gnd_net_),
            .in3(N__7802),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ),
            .clk(N__11148),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_12_6_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_12_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_12_6_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_7_LC_12_6_6  (
            .in0(_gnd_net_),
            .in1(N__8767),
            .in2(_gnd_net_),
            .in3(N__7799),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11148),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_12_6_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_12_6_7 .LUT_INIT=16'b0001010100101010;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_3_LC_12_6_7  (
            .in0(N__8630),
            .in1(N__7796),
            .in2(N__7790),
            .in3(N__7775),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11148),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_1_LC_12_7_0 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_1_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_1_LC_12_7_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_CIA.VMA_RNO_1_LC_12_7_0  (
            .in0(_gnd_net_),
            .in1(N__8762),
            .in2(_gnd_net_),
            .in3(N__8828),
            .lcout(\U409_CIA.CLK_CIA6_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_12_7_1 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_12_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_12_7_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_1_LC_12_7_1  (
            .in0(N__8736),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8800),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11147),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_2_LC_12_7_3 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_2_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_2_LC_12_7_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_CIA.VMA_RNO_2_LC_12_7_3  (
            .in0(N__8631),
            .in1(N__8601),
            .in2(N__8700),
            .in3(N__8799),
            .lcout(),
            .ltout(\U409_CIA.un1_CIA_CLK_COUNT_3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_0_LC_12_7_4 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_0_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_0_LC_12_7_4 .LUT_INIT=16'b0100000010000000;
    LogicCell40 \U409_CIA.VMA_RNO_0_LC_12_7_4  (
            .in0(N__8661),
            .in1(N__7895),
            .in2(N__7889),
            .in3(N__8735),
            .lcout(),
            .ltout(\U409_CIA.VMA_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_LC_12_7_5 .C_ON=1'b0;
    defparam \U409_CIA.VMA_LC_12_7_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.VMA_LC_12_7_5 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \U409_CIA.VMA_LC_12_7_5  (
            .in0(N__8737),
            .in1(N__7886),
            .in2(N__7865),
            .in3(N__8544),
            .lcout(\U409_CIA.VMAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11147),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_7_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_7_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_7_7  (
            .in0(_gnd_net_),
            .in1(N__9311),
            .in2(_gnd_net_),
            .in3(N__9292),
            .lcout(\U409_TRANSFER_ACK.N_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_12_8_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_12_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_12_8_0  (
            .in0(N__8204),
            .in1(N__8118),
            .in2(N__8186),
            .in3(N__8290),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_12_8_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_12_8_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_12_8_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_12_8_1  (
            .in0(N__8119),
            .in1(N__8184),
            .in2(_gnd_net_),
            .in3(N__8206),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__8090));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_12_8_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_12_8_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_12_8_2 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_12_8_2  (
            .in0(N__8205),
            .in1(N__8120),
            .in2(_gnd_net_),
            .in3(N__7849),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__8090));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_12_8_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_12_8_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_12_8_3  (
            .in0(N__8117),
            .in1(N__8289),
            .in2(N__8231),
            .in3(N__8244),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_12_8_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_12_8_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_12_8_4  (
            .in0(N__8312),
            .in1(N__8267),
            .in2(N__7823),
            .in3(N__8164),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_12_8_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_12_8_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_12_8_5  (
            .in0(N__8311),
            .in1(N__8288),
            .in2(N__8270),
            .in3(N__8245),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_12_8_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_12_8_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_12_8_6  (
            .in0(N__8126),
            .in1(N__8228),
            .in2(N__8210),
            .in3(N__8165),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_12_8_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_12_8_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_12_8_7  (
            .in0(_gnd_net_),
            .in1(N__8203),
            .in2(_gnd_net_),
            .in3(N__8180),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_12_9_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_12_9_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_12_9_1 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_12_9_1  (
            .in0(N__8495),
            .in1(N__8140),
            .in2(_gnd_net_),
            .in3(N__8155),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ),
            .ce(),
            .sr(N__8085));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_12_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_12_9_3 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_12_9_3 .LUT_INIT=16'b0001000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_12_9_3  (
            .in0(N__7997),
            .in1(N__8125),
            .in2(N__9872),
            .in3(N__8141),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ),
            .ce(),
            .sr(N__8085));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_2_LC_12_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_2_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_2_LC_12_10_0 .LUT_INIT=16'b0000000011101010;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_2_LC_12_10_0  (
            .in0(N__8054),
            .in1(N__7901),
            .in2(N__8033),
            .in3(N__8009),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_2 ),
            .ltout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_12_10_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_12_10_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_12_10_1 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_12_10_1  (
            .in0(N__9864),
            .in1(_gnd_net_),
            .in2(N__7955),
            .in3(N__8476),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .ce(),
            .sr(N__9731));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_11_LC_12_10_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_11_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_11_LC_12_10_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_11_LC_12_10_2  (
            .in0(N__7952),
            .in1(N__7928),
            .in2(N__9024),
            .in3(N__7919),
            .lcout(U409_ADDRESS_DECODE_AUTOVECTOR_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_12_10_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_12_10_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_12_10_3  (
            .in0(N__8483),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8983),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_12_10_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_12_10_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_12_10_4 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_12_10_4  (
            .in0(N__8477),
            .in1(N__9865),
            .in2(N__8468),
            .in3(N__9212),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .ce(),
            .sr(N__9731));
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_3.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_3.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_19_3 (
            .in0(N__8969),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_13_4_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_13_4_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_13_4_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_13_4_0  (
            .in0(N__8395),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8456),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS0n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNI692L_0_LC_13_4_7 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNI692L_0_LC_13_4_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNI692L_0_LC_13_4_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_CIA.VMA_RNI692L_0_LC_13_4_7  (
            .in0(N__8928),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8549),
            .lcout(CIA_ENABLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_13_5_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_13_5_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_13_5_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_13_5_1  (
            .in0(_gnd_net_),
            .in1(N__8396),
            .in2(_gnd_net_),
            .in3(N__8384),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS1n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_13_6_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_13_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_13_6_6 .LUT_INIT=16'b0111101000101010;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_1_LC_13_6_6  (
            .in0(N__9332),
            .in1(N__8321),
            .in2(N__8573),
            .in3(N__9338),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .ce(),
            .sr(N__9744));
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_13_7_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_13_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_13_7_3 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_0_LC_13_7_3  (
            .in0(N__8568),
            .in1(N__9272),
            .in2(_gnd_net_),
            .in3(N__9344),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(N__9737));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_13_7_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_13_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_13_7_4 .LUT_INIT=16'b0101111100001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_LC_13_7_4  (
            .in0(N__9331),
            .in1(N__9353),
            .in2(N__8572),
            .in3(N__8507),
            .lcout(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(N__9737));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_13_7_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_13_7_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_13_7_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_13_7_5  (
            .in0(N__8948),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8545),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(N__9737));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_13_7_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_13_7_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_13_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_13_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9293),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(N__9737));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_13_8_0 .C_ON=1'b1;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_13_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_13_8_0  (
            .in0(_gnd_net_),
            .in1(N__9437),
            .in2(N__9958),
            .in3(N__9949),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_13_8_0_),
            .carryout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_1_LC_13_8_1 .C_ON=1'b1;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_1_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_1_LC_13_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_1_LC_13_8_1  (
            .in0(_gnd_net_),
            .in1(N__9480),
            .in2(_gnd_net_),
            .in3(N__8528),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_0 ),
            .carryout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_2_LC_13_8_2 .C_ON=1'b1;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_2_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_2_LC_13_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_2_LC_13_8_2  (
            .in0(_gnd_net_),
            .in1(N__9244),
            .in2(_gnd_net_),
            .in3(N__8525),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_1 ),
            .carryout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_3_LC_13_8_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_3_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_3_LC_13_8_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_3_LC_13_8_3  (
            .in0(_gnd_net_),
            .in1(N__9256),
            .in2(_gnd_net_),
            .in3(N__8522),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_13_8_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_13_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_13_8_4 .LUT_INIT=16'b0000100010001000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_13_8_4  (
            .in0(N__8976),
            .in1(N__8519),
            .in2(N__9959),
            .in3(N__10036),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9825),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_13_8_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_13_8_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_13_8_5 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_13_8_5  (
            .in0(N__10035),
            .in1(N__8513),
            .in2(N__9021),
            .in3(N__9957),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9825),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_START_RNO_1_LC_13_8_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_START_RNO_1_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_START_RNO_1_LC_13_8_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.TACK_START_RNO_1_LC_13_8_6  (
            .in0(_gnd_net_),
            .in1(N__8506),
            .in2(_gnd_net_),
            .in3(N__8494),
            .lcout(\U409_TRANSFER_ACK.TACK_START_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_13_8_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_13_8_7 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_13_8_7  (
            .in0(N__10037),
            .in1(N__9956),
            .in2(N__9022),
            .in3(N__9230),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9825),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_START_LC_13_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_START_LC_13_9_5 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.TACK_START_LC_13_9_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_START_LC_13_9_5  (
            .in0(N__9224),
            .in1(N__9211),
            .in2(N__9192),
            .in3(N__9200),
            .lcout(\U409_TRANSFER_ACK.TACK_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9159),
            .ce(),
            .sr(N__8849));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_13_10_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_13_10_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_13_10_4 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_13_10_4  (
            .in0(N__10034),
            .in1(N__9131),
            .in2(N__9023),
            .in3(N__9936),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9819),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_START_RNO_0_LC_13_11_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_START_RNO_0_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_START_RNO_0_LC_13_11_1 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_START_RNO_0_LC_13_11_1  (
            .in0(N__9096),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8984),
            .lcout(\U409_TRANSFER_ACK.TACK_RST_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_14_6_0 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_14_6_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_0_LC_14_6_0  (
            .in0(N__8834),
            .in1(N__8807),
            .in2(N__8771),
            .in3(N__8741),
            .lcout(),
            .ltout(\U409_CIA.CLK_CIA6_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_LC_14_6_1 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_LC_14_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CLK_CIA_LC_14_6_1 .LUT_INIT=16'b1010101001101010;
    LogicCell40 \U409_CIA.CLK_CIA_LC_14_6_1  (
            .in0(N__9620),
            .in1(N__8579),
            .in2(N__8705),
            .in3(N__8702),
            .lcout(CLK_CIA_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11146),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_6_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_6_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_6_5  (
            .in0(N__9583),
            .in1(N__9656),
            .in2(N__9527),
            .in3(N__9566),
            .lcout(\U409_TICK.TICK503_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_14_6_7 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_14_6_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_14_6_7 .LUT_INIT=16'b0000000000011000;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_1_LC_14_6_7  (
            .in0(N__8666),
            .in1(N__8636),
            .in2(N__9627),
            .in3(N__8606),
            .lcout(\U409_CIA.CLK_CIA_r_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_14_7_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_14_7_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_14_7_0  (
            .in0(N__9870),
            .in1(N__9597),
            .in2(_gnd_net_),
            .in3(N__9265),
            .lcout(\U409_TRANSFER_ACK.N_17_mux ),
            .ltout(\U409_TRANSFER_ACK.N_17_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_14_7_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_14_7_1 .LUT_INIT=16'b0001101101011111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_14_7_1  (
            .in0(N__9329),
            .in1(N__9309),
            .in2(N__9347),
            .in3(N__9290),
            .lcout(\U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_14_7_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_14_7_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_14_7_2  (
            .in0(_gnd_net_),
            .in1(N__9598),
            .in2(_gnd_net_),
            .in3(N__9266),
            .lcout(\U409_TRANSFER_ACK.N_3_0 ),
            .ltout(\U409_TRANSFER_ACK.N_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_14_7_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_14_7_3 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_14_7_3  (
            .in0(N__9330),
            .in1(N__9310),
            .in2(N__9296),
            .in3(N__9291),
            .lcout(\U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_1_LC_14_7_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_1_LC_14_7_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_1_LC_14_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_TICK.COUNTER50_1_LC_14_7_5  (
            .in0(_gnd_net_),
            .in1(N__10169),
            .in2(_gnd_net_),
            .in3(N__9584),
            .lcout(\U409_TICK.COUNTER50Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10869),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_14_8_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_14_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_14_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_1_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9599),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .ce(),
            .sr(N__9738));
    defparam \U409_TRANSFER_ACK.ROM_TACK_STATE_ns_1_0__m6_LC_14_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_STATE_ns_1_0__m6_LC_14_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_STATE_ns_1_0__m6_LC_14_9_3 .LUT_INIT=16'b0001100000000001;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_STATE_ns_1_0__m6_LC_14_9_3  (
            .in0(N__9463),
            .in1(N__9481),
            .in2(N__9509),
            .in3(N__9435),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.N_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_STATE_ns_1_0__m10_LC_14_9_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_STATE_ns_1_0__m10_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_STATE_ns_1_0__m10_LC_14_9_4 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_STATE_ns_1_0__m10_LC_14_9_4  (
            .in0(N__9257),
            .in1(N__9245),
            .in2(N__9233),
            .in3(N__9419),
            .lcout(\U409_TRANSFER_ACK.N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_STATE_ns_1_0__m8_LC_14_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_STATE_ns_1_0__m8_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_STATE_ns_1_0__m8_LC_14_9_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_STATE_ns_1_0__m8_LC_14_9_5  (
            .in0(N__9508),
            .in1(N__9482),
            .in2(N__9467),
            .in3(N__9436),
            .lcout(\U409_TRANSFER_ACK.N_19_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_STATE_0_LC_14_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_STATE_0_LC_14_10_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_STATE_0_LC_14_10_5 .LUT_INIT=16'b0001000111111010;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_STATE_0_LC_14_10_5  (
            .in0(N__10015),
            .in1(N__10082),
            .in2(N__9982),
            .in3(N__9934),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9822),
            .ce(),
            .sr(N__9734));
    defparam \U409_TICK.TICK60_LC_15_5_0 .C_ON=1'b0;
    defparam \U409_TICK.TICK60_LC_15_5_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK60_LC_15_5_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \U409_TICK.TICK60_LC_15_5_0  (
            .in0(N__10320),
            .in1(N__9397),
            .in2(N__10262),
            .in3(N__10284),
            .lcout(TICK60_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10868),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_15_5_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_15_5_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_15_5_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER60_RNICDC71_14_LC_15_5_1  (
            .in0(N__10619),
            .in1(N__10640),
            .in2(N__10685),
            .in3(N__11090),
            .lcout(\U409_TICK.TICK603_9 ),
            .ltout(\U409_TICK.TICK603_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_6_LC_15_5_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_6_LC_15_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_6_LC_15_5_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_6_LC_15_5_2  (
            .in0(N__10319),
            .in1(N__10283),
            .in2(N__9386),
            .in3(N__10667),
            .lcout(\U409_TICK.COUNTER60Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10868),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK50_LC_15_5_3 .C_ON=1'b0;
    defparam \U409_TICK.TICK50_LC_15_5_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK50_LC_15_5_3 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \U409_TICK.TICK50_LC_15_5_3  (
            .in0(N__10987),
            .in1(N__11032),
            .in2(N__10946),
            .in3(N__9370),
            .lcout(TICK50_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10868),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_15_5_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_15_5_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_15_5_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_TICK.COUNTER60_RNIHJU51_4_LC_15_5_4  (
            .in0(N__10340),
            .in1(N__10366),
            .in2(_gnd_net_),
            .in3(N__10424),
            .lcout(),
            .ltout(\U409_TICK.TICK603_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_15_5_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_15_5_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_15_5_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER60_RNI335G2_11_LC_15_5_5  (
            .in0(N__9686),
            .in1(N__10580),
            .in2(N__9359),
            .in3(N__10388),
            .lcout(\U409_TICK.TICK603_14 ),
            .ltout(\U409_TICK.TICK603_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_4_LC_15_5_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_4_LC_15_5_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_4_LC_15_5_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_4_LC_15_5_6  (
            .in0(N__10318),
            .in1(N__10258),
            .in2(N__9356),
            .in3(N__10352),
            .lcout(\U409_TICK.COUNTER60Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10868),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_6_LC_15_5_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_6_LC_15_5_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_6_LC_15_5_7 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_6_LC_15_5_7  (
            .in0(N__10945),
            .in1(N__11031),
            .in2(N__9542),
            .in3(N__10993),
            .lcout(\U409_TICK.COUNTER50Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10868),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_15_6_0 .C_ON=1'b1;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_15_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_15_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_15_6_0  (
            .in0(_gnd_net_),
            .in1(N__9582),
            .in2(N__10164),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_6_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_2_LC_15_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_2_LC_15_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_2_LC_15_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_2_LC_15_6_1  (
            .in0(_gnd_net_),
            .in1(N__9565),
            .in2(_gnd_net_),
            .in3(N__9554),
            .lcout(\U409_TICK.COUNTER50Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .clk(N__10870),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_3_LC_15_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_3_LC_15_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_3_LC_15_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_3_LC_15_6_2  (
            .in0(_gnd_net_),
            .in1(N__10225),
            .in2(_gnd_net_),
            .in3(N__9551),
            .lcout(\U409_TICK.COUNTER50Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .clk(N__10870),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_4_LC_15_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_4_LC_15_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_4_LC_15_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_4_LC_15_6_3  (
            .in0(_gnd_net_),
            .in1(N__10492),
            .in2(_gnd_net_),
            .in3(N__9548),
            .lcout(\U409_TICK.COUNTER50Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .clk(N__10870),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_15_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_15_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_15_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_5_LC_15_6_4  (
            .in0(_gnd_net_),
            .in1(N__10519),
            .in2(_gnd_net_),
            .in3(N__9545),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_15_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_15_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_15_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_6_LC_15_6_5  (
            .in0(_gnd_net_),
            .in1(N__10102),
            .in2(_gnd_net_),
            .in3(N__9533),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_7_LC_15_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_7_LC_15_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_7_LC_15_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_7_LC_15_6_6  (
            .in0(_gnd_net_),
            .in1(N__10507),
            .in2(_gnd_net_),
            .in3(N__9530),
            .lcout(\U409_TICK.COUNTER50Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .clk(N__10870),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_8_LC_15_6_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_8_LC_15_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_8_LC_15_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_8_LC_15_6_7  (
            .in0(_gnd_net_),
            .in1(N__9523),
            .in2(_gnd_net_),
            .in3(N__9512),
            .lcout(\U409_TICK.COUNTER50Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .clk(N__10870),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_15_7_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_15_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_9_LC_15_7_0  (
            .in0(_gnd_net_),
            .in1(N__10117),
            .in2(_gnd_net_),
            .in3(N__9680),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_15_7_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_10_LC_15_7_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_10_LC_15_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_10_LC_15_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_10_LC_15_7_1  (
            .in0(_gnd_net_),
            .in1(N__10189),
            .in2(_gnd_net_),
            .in3(N__9677),
            .lcout(\U409_TICK.COUNTER50Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .clk(N__10872),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_15_7_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_15_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_15_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_11_LC_15_7_2  (
            .in0(_gnd_net_),
            .in1(N__10129),
            .in2(_gnd_net_),
            .in3(N__9674),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_12_LC_15_7_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_12_LC_15_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_12_LC_15_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_12_LC_15_7_3  (
            .in0(_gnd_net_),
            .in1(N__10204),
            .in2(_gnd_net_),
            .in3(N__9671),
            .lcout(\U409_TICK.COUNTER50Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .clk(N__10872),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_15_7_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_15_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_15_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_13_LC_15_7_4  (
            .in0(_gnd_net_),
            .in1(N__10892),
            .in2(_gnd_net_),
            .in3(N__9668),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_15_7_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_15_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_14_LC_15_7_5  (
            .in0(_gnd_net_),
            .in1(N__10480),
            .in2(_gnd_net_),
            .in3(N__9665),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_15_7_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_15_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_15_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_15_LC_15_7_6  (
            .in0(_gnd_net_),
            .in1(N__10459),
            .in2(_gnd_net_),
            .in3(N__9662),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_16_LC_15_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_16_LC_15_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_16_LC_15_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER50_16_LC_15_7_7  (
            .in0(_gnd_net_),
            .in1(N__9655),
            .in2(_gnd_net_),
            .in3(N__9659),
            .lcout(\U409_TICK.COUNTER50Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10872),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_15_8_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_15_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_15_8_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_0_LC_15_8_4  (
            .in0(N__9628),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .ce(),
            .sr(N__9745));
    defparam \U409_TRANSFER_ACK.ROM_TACK_STATE_1_LC_15_9_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_STATE_1_LC_15_9_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_STATE_1_LC_15_9_4 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_STATE_1_LC_15_9_4  (
            .in0(N__10011),
            .in1(N__10080),
            .in2(_gnd_net_),
            .in3(N__9932),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9832),
            .ce(),
            .sr(N__9739));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_15_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_15_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_15_9_6 .LUT_INIT=16'b1010111000001010;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_LC_15_9_6  (
            .in0(N__10058),
            .in1(N__10081),
            .in2(N__10023),
            .in3(N__9933),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9832),
            .ce(),
            .sr(N__9739));
    defparam \U409_TRANSFER_ACK.ROMENn_LC_15_10_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_15_10_6 .SEQ_MODE=4'b1001;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_15_10_6 .LUT_INIT=16'b1110111010001100;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_LC_15_10_6  (
            .in0(N__10016),
            .in1(N__9883),
            .in2(N__9986),
            .in3(N__9935),
            .lcout(ROMENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9826),
            .ce(),
            .sr(N__9735));
    defparam \U409_TICK.COUNTER60_0_LC_16_5_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_0_LC_16_5_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_0_LC_16_5_0 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U409_TICK.COUNTER60_0_LC_16_5_0  (
            .in0(N__10253),
            .in1(N__10285),
            .in2(N__10430),
            .in3(N__10310),
            .lcout(\U409_TICK.COUNTER60Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10871),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_15_LC_16_5_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_15_LC_16_5_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_15_LC_16_5_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_15_LC_16_5_1  (
            .in0(N__10287),
            .in1(N__10256),
            .in2(N__10321),
            .in3(N__11057),
            .lcout(\U409_TICK.COUNTER60Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10871),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_16_5_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_16_5_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_16_5_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER60_RNIDB4S_16_LC_16_5_2  (
            .in0(N__10559),
            .in1(N__10403),
            .in2(N__10448),
            .in3(N__11044),
            .lcout(\U409_TICK.TICK603_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_8_LC_16_5_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_8_LC_16_5_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_8_LC_16_5_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_8_LC_16_5_3  (
            .in0(N__10288),
            .in1(N__10257),
            .in2(N__10322),
            .in3(N__10628),
            .lcout(\U409_TICK.COUNTER60Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10871),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_9_LC_16_5_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_9_LC_16_5_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_9_LC_16_5_4 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_9_LC_16_5_4  (
            .in0(N__10254),
            .in1(N__10289),
            .in2(N__10607),
            .in3(N__10317),
            .lcout(\U409_TICK.COUNTER60Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10871),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_1_LC_16_5_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_1_LC_16_5_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_1_LC_16_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_TICK.COUNTER60_1_LC_16_5_5  (
            .in0(_gnd_net_),
            .in1(N__10425),
            .in2(_gnd_net_),
            .in3(N__10447),
            .lcout(\U409_TICK.COUNTER60Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10871),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_16_5_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_16_5_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_16_5_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U409_TICK.COUNTER60_RNI2USG_10_LC_16_5_6  (
            .in0(N__10595),
            .in1(N__11069),
            .in2(N__10544),
            .in3(N__10655),
            .lcout(\U409_TICK.TICK603_10 ),
            .ltout(\U409_TICK.TICK603_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_14_LC_16_5_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_14_LC_16_5_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_14_LC_16_5_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_14_LC_16_5_7  (
            .in0(N__10286),
            .in1(N__10255),
            .in2(N__10229),
            .in3(N__11078),
            .lcout(\U409_TICK.COUNTER60Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10871),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_16_6_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_16_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_16_6_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_TICK.COUNTER50_RNID6CP_3_LC_16_6_0  (
            .in0(N__10520),
            .in1(N__10226),
            .in2(_gnd_net_),
            .in3(N__10157),
            .lcout(),
            .ltout(\U409_TICK.TICK503_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_16_6_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_16_6_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_16_6_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER50_RNITU182_10_LC_16_6_1  (
            .in0(N__10214),
            .in1(N__10205),
            .in2(N__10193),
            .in3(N__10190),
            .lcout(\U409_TICK.TICK503_14 ),
            .ltout(\U409_TICK.TICK503_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_9_LC_16_6_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_9_LC_16_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_9_LC_16_6_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_9_LC_16_6_2  (
            .in0(N__11023),
            .in1(N__10932),
            .in2(N__10178),
            .in3(N__10175),
            .lcout(\U409_TICK.COUNTER50Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10873),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_0_LC_16_6_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_0_LC_16_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_0_LC_16_6_3 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U409_TICK.COUNTER50_0_LC_16_6_3  (
            .in0(N__10928),
            .in1(N__11024),
            .in2(N__10165),
            .in3(N__10983),
            .lcout(\U409_TICK.COUNTER50Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10873),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_11_LC_16_6_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_11_LC_16_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_11_LC_16_6_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_11_LC_16_6_4  (
            .in0(N__10981),
            .in1(N__10930),
            .in2(N__11033),
            .in3(N__10136),
            .lcout(\U409_TICK.COUNTER50Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10873),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_16_6_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_16_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_16_6_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNIH14V_11_LC_16_6_5  (
            .in0(N__10130),
            .in1(N__10118),
            .in2(N__10106),
            .in3(N__10891),
            .lcout(\U409_TICK.TICK503_9 ),
            .ltout(\U409_TICK.TICK503_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_14_LC_16_6_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_14_LC_16_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_14_LC_16_6_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_14_LC_16_6_6  (
            .in0(N__10982),
            .in1(N__10931),
            .in2(N__10091),
            .in3(N__10088),
            .lcout(\U409_TICK.COUNTER50Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10873),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_5_LC_16_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_5_LC_16_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_5_LC_16_6_7 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \U409_TICK.COUNTER50_5_LC_16_6_7  (
            .in0(N__10929),
            .in1(N__10526),
            .in2(N__10994),
            .in3(N__11028),
            .lcout(\U409_TICK.COUNTER50Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10873),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_16_7_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_16_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_16_7_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNII24V_14_LC_16_7_5  (
            .in0(N__10460),
            .in1(N__10508),
            .in2(N__10496),
            .in3(N__10481),
            .lcout(\U409_TICK.TICK503_10 ),
            .ltout(\U409_TICK.TICK503_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_15_LC_16_7_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_15_LC_16_7_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_15_LC_16_7_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_15_LC_16_7_6  (
            .in0(N__11029),
            .in1(N__10988),
            .in2(N__10469),
            .in3(N__10466),
            .lcout(\U409_TICK.COUNTER50Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10875),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_17_5_0 .C_ON=1'b1;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_17_5_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_17_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_17_5_0  (
            .in0(_gnd_net_),
            .in1(N__10443),
            .in2(N__10429),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_5_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_2_LC_17_5_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_2_LC_17_5_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_2_LC_17_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_2_LC_17_5_1  (
            .in0(_gnd_net_),
            .in1(N__10402),
            .in2(_gnd_net_),
            .in3(N__10391),
            .lcout(\U409_TICK.COUNTER60Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .clk(N__10874),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_3_LC_17_5_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_3_LC_17_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_3_LC_17_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_3_LC_17_5_2  (
            .in0(_gnd_net_),
            .in1(N__10384),
            .in2(_gnd_net_),
            .in3(N__10373),
            .lcout(\U409_TICK.COUNTER60Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .clk(N__10874),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_17_5_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_17_5_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_17_5_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_4_LC_17_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10370),
            .in3(N__10343),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_5_LC_17_5_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_5_LC_17_5_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_5_LC_17_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_5_LC_17_5_4  (
            .in0(_gnd_net_),
            .in1(N__10336),
            .in2(_gnd_net_),
            .in3(N__10325),
            .lcout(\U409_TICK.COUNTER60Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .clk(N__10874),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_17_5_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_17_5_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_17_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_6_LC_17_5_5  (
            .in0(_gnd_net_),
            .in1(N__10681),
            .in2(_gnd_net_),
            .in3(N__10658),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_7_LC_17_5_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_7_LC_17_5_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_7_LC_17_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_7_LC_17_5_6  (
            .in0(_gnd_net_),
            .in1(N__10654),
            .in2(_gnd_net_),
            .in3(N__10643),
            .lcout(\U409_TICK.COUNTER60Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .clk(N__10874),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_17_5_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_17_5_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_17_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_8_LC_17_5_7  (
            .in0(_gnd_net_),
            .in1(N__10639),
            .in2(_gnd_net_),
            .in3(N__10622),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_17_6_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_17_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_17_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_9_LC_17_6_0  (
            .in0(_gnd_net_),
            .in1(N__10618),
            .in2(_gnd_net_),
            .in3(N__10598),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_17_6_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_10_LC_17_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_10_LC_17_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_10_LC_17_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_10_LC_17_6_1  (
            .in0(_gnd_net_),
            .in1(N__10594),
            .in2(_gnd_net_),
            .in3(N__10583),
            .lcout(\U409_TICK.COUNTER60Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .clk(N__10876),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_11_LC_17_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_11_LC_17_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_11_LC_17_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_11_LC_17_6_2  (
            .in0(_gnd_net_),
            .in1(N__10573),
            .in2(_gnd_net_),
            .in3(N__10562),
            .lcout(\U409_TICK.COUNTER60Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .clk(N__10876),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_12_LC_17_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_12_LC_17_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_12_LC_17_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_12_LC_17_6_3  (
            .in0(_gnd_net_),
            .in1(N__10558),
            .in2(_gnd_net_),
            .in3(N__10547),
            .lcout(\U409_TICK.COUNTER60Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .clk(N__10876),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_13_LC_17_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_13_LC_17_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_13_LC_17_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_13_LC_17_6_4  (
            .in0(_gnd_net_),
            .in1(N__10540),
            .in2(_gnd_net_),
            .in3(N__10529),
            .lcout(\U409_TICK.COUNTER60Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .clk(N__10876),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_17_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_17_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_17_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_14_LC_17_6_5  (
            .in0(_gnd_net_),
            .in1(N__11089),
            .in2(_gnd_net_),
            .in3(N__11072),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_17_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_17_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_17_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_15_LC_17_6_6  (
            .in0(_gnd_net_),
            .in1(N__11068),
            .in2(_gnd_net_),
            .in3(N__11051),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_16_LC_17_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_16_LC_17_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_16_LC_17_6_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER60_16_LC_17_6_7  (
            .in0(_gnd_net_),
            .in1(N__11045),
            .in2(_gnd_net_),
            .in3(N__11048),
            .lcout(\U409_TICK.COUNTER60Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10876),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_13_LC_17_7_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_13_LC_17_7_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_13_LC_17_7_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_13_LC_17_7_6  (
            .in0(N__11030),
            .in1(N__10989),
            .in2(N__10941),
            .in3(N__10901),
            .lcout(\U409_TICK.COUNTER50Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10877),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PCS1_LC_20_2_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PCS1_LC_20_2_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PCS1_LC_20_2_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_ADDRESS_DECODE.PCS1_LC_20_2_4  (
            .in0(N__10804),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10766),
            .lcout(PCS1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.SCS0_LC_20_3_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.SCS0_LC_20_3_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.SCS0_LC_20_3_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U409_ADDRESS_DECODE.SCS0_LC_20_3_2  (
            .in0(_gnd_net_),
            .in1(N__10767),
            .in2(_gnd_net_),
            .in3(N__10720),
            .lcout(SCS0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PCS0_LC_22_2_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PCS0_LC_22_2_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PCS0_LC_22_2_0 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \U409_ADDRESS_DECODE.PCS0_LC_22_2_0  (
            .in0(N__10768),
            .in1(N__10805),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PCS0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.SCS1_LC_22_3_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.SCS1_LC_22_3_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.SCS1_LC_22_3_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_ADDRESS_DECODE.SCS1_LC_22_3_2  (
            .in0(_gnd_net_),
            .in1(N__10769),
            .in2(_gnd_net_),
            .in3(N__10721),
            .lcout(SCS1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_22_10_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_22_10_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_22_10_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_22_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam AGNUS_CLK_obuf_RNO_LC_24_14_2.C_ON=1'b0;
    defparam AGNUS_CLK_obuf_RNO_LC_24_14_2.SEQ_MODE=4'b0000;
    defparam AGNUS_CLK_obuf_RNO_LC_24_14_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 AGNUS_CLK_obuf_RNO_LC_24_14_2 (
            .in0(N__11153),
            .in1(N__11126),
            .in2(_gnd_net_),
            .in3(N__11114),
            .lcout(AGNUS_CLK_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U409_TOP

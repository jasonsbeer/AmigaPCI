// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Dec 13 2024 16:29:06

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U409_TOP" view "INTERFACE"

module U409_TOP (
    A,
    RnW,
    TT1,
    TICK50,
    nROMEN,
    nCIACS1,
    TT0,
    TICK60,
    LBENn,
    CLKCIA,
    CLK6,
    CLK40_IN,
    CLK28_IN,
    TSn,
    nBUFEN,
    nREGSPACE,
    nRAMSPACE,
    RESETn,
    OVL,
    TACKn,
    nCIACS0,
    PORTSIZE);

    input [31:1] A;
    input RnW;
    input TT1;
    output TICK50;
    output nROMEN;
    output nCIACS1;
    input TT0;
    output TICK60;
    input LBENn;
    output CLKCIA;
    input CLK6;
    input CLK40_IN;
    input CLK28_IN;
    input TSn;
    output nBUFEN;
    output nREGSPACE;
    output nRAMSPACE;
    input RESETn;
    input OVL;
    inout TACKn;
    output nCIACS0;
    output PORTSIZE;

    wire N__6036;
    wire N__6035;
    wire N__6034;
    wire N__6026;
    wire N__6025;
    wire N__6024;
    wire N__6015;
    wire N__6014;
    wire N__6013;
    wire N__6006;
    wire N__6005;
    wire N__6004;
    wire N__5997;
    wire N__5996;
    wire N__5995;
    wire N__5988;
    wire N__5987;
    wire N__5986;
    wire N__5979;
    wire N__5978;
    wire N__5977;
    wire N__5970;
    wire N__5969;
    wire N__5968;
    wire N__5961;
    wire N__5960;
    wire N__5959;
    wire N__5952;
    wire N__5951;
    wire N__5950;
    wire N__5943;
    wire N__5942;
    wire N__5941;
    wire N__5934;
    wire N__5933;
    wire N__5932;
    wire N__5925;
    wire N__5924;
    wire N__5923;
    wire N__5916;
    wire N__5915;
    wire N__5914;
    wire N__5907;
    wire N__5906;
    wire N__5905;
    wire N__5898;
    wire N__5897;
    wire N__5896;
    wire N__5889;
    wire N__5888;
    wire N__5887;
    wire N__5880;
    wire N__5879;
    wire N__5878;
    wire N__5871;
    wire N__5870;
    wire N__5869;
    wire N__5862;
    wire N__5861;
    wire N__5860;
    wire N__5853;
    wire N__5852;
    wire N__5851;
    wire N__5844;
    wire N__5843;
    wire N__5842;
    wire N__5835;
    wire N__5834;
    wire N__5833;
    wire N__5826;
    wire N__5825;
    wire N__5824;
    wire N__5817;
    wire N__5816;
    wire N__5815;
    wire N__5808;
    wire N__5807;
    wire N__5806;
    wire N__5799;
    wire N__5798;
    wire N__5797;
    wire N__5790;
    wire N__5789;
    wire N__5788;
    wire N__5781;
    wire N__5780;
    wire N__5779;
    wire N__5772;
    wire N__5771;
    wire N__5770;
    wire N__5763;
    wire N__5762;
    wire N__5761;
    wire N__5754;
    wire N__5753;
    wire N__5752;
    wire N__5745;
    wire N__5744;
    wire N__5743;
    wire N__5736;
    wire N__5735;
    wire N__5734;
    wire N__5727;
    wire N__5726;
    wire N__5725;
    wire N__5708;
    wire N__5707;
    wire N__5702;
    wire N__5699;
    wire N__5696;
    wire N__5695;
    wire N__5694;
    wire N__5693;
    wire N__5692;
    wire N__5689;
    wire N__5684;
    wire N__5679;
    wire N__5672;
    wire N__5671;
    wire N__5670;
    wire N__5669;
    wire N__5668;
    wire N__5667;
    wire N__5666;
    wire N__5661;
    wire N__5658;
    wire N__5649;
    wire N__5642;
    wire N__5641;
    wire N__5640;
    wire N__5637;
    wire N__5636;
    wire N__5633;
    wire N__5630;
    wire N__5625;
    wire N__5618;
    wire N__5615;
    wire N__5612;
    wire N__5611;
    wire N__5608;
    wire N__5605;
    wire N__5604;
    wire N__5601;
    wire N__5600;
    wire N__5599;
    wire N__5596;
    wire N__5593;
    wire N__5592;
    wire N__5591;
    wire N__5590;
    wire N__5587;
    wire N__5584;
    wire N__5583;
    wire N__5580;
    wire N__5579;
    wire N__5578;
    wire N__5577;
    wire N__5576;
    wire N__5573;
    wire N__5570;
    wire N__5563;
    wire N__5562;
    wire N__5559;
    wire N__5554;
    wire N__5549;
    wire N__5546;
    wire N__5543;
    wire N__5542;
    wire N__5541;
    wire N__5538;
    wire N__5537;
    wire N__5536;
    wire N__5535;
    wire N__5532;
    wire N__5527;
    wire N__5524;
    wire N__5523;
    wire N__5520;
    wire N__5517;
    wire N__5514;
    wire N__5509;
    wire N__5504;
    wire N__5497;
    wire N__5494;
    wire N__5487;
    wire N__5484;
    wire N__5469;
    wire N__5466;
    wire N__5463;
    wire N__5460;
    wire N__5455;
    wire N__5450;
    wire N__5447;
    wire N__5444;
    wire N__5441;
    wire N__5438;
    wire N__5435;
    wire N__5432;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5419;
    wire N__5418;
    wire N__5415;
    wire N__5412;
    wire N__5409;
    wire N__5406;
    wire N__5403;
    wire N__5400;
    wire N__5397;
    wire N__5394;
    wire N__5391;
    wire N__5384;
    wire N__5381;
    wire N__5378;
    wire N__5375;
    wire N__5372;
    wire N__5369;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5354;
    wire N__5351;
    wire N__5350;
    wire N__5349;
    wire N__5346;
    wire N__5345;
    wire N__5342;
    wire N__5339;
    wire N__5336;
    wire N__5335;
    wire N__5332;
    wire N__5327;
    wire N__5326;
    wire N__5323;
    wire N__5322;
    wire N__5319;
    wire N__5316;
    wire N__5313;
    wire N__5310;
    wire N__5307;
    wire N__5304;
    wire N__5301;
    wire N__5298;
    wire N__5293;
    wire N__5288;
    wire N__5285;
    wire N__5282;
    wire N__5279;
    wire N__5276;
    wire N__5267;
    wire N__5266;
    wire N__5263;
    wire N__5260;
    wire N__5257;
    wire N__5254;
    wire N__5251;
    wire N__5248;
    wire N__5243;
    wire N__5240;
    wire N__5237;
    wire N__5234;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5222;
    wire N__5219;
    wire N__5216;
    wire N__5213;
    wire N__5210;
    wire N__5207;
    wire N__5206;
    wire N__5205;
    wire N__5198;
    wire N__5195;
    wire N__5194;
    wire N__5193;
    wire N__5192;
    wire N__5189;
    wire N__5188;
    wire N__5185;
    wire N__5178;
    wire N__5175;
    wire N__5168;
    wire N__5165;
    wire N__5164;
    wire N__5161;
    wire N__5158;
    wire N__5155;
    wire N__5150;
    wire N__5149;
    wire N__5148;
    wire N__5147;
    wire N__5146;
    wire N__5139;
    wire N__5136;
    wire N__5133;
    wire N__5126;
    wire N__5125;
    wire N__5124;
    wire N__5121;
    wire N__5120;
    wire N__5117;
    wire N__5114;
    wire N__5109;
    wire N__5102;
    wire N__5101;
    wire N__5100;
    wire N__5099;
    wire N__5096;
    wire N__5093;
    wire N__5090;
    wire N__5085;
    wire N__5078;
    wire N__5077;
    wire N__5076;
    wire N__5073;
    wire N__5068;
    wire N__5063;
    wire N__5062;
    wire N__5061;
    wire N__5060;
    wire N__5057;
    wire N__5052;
    wire N__5047;
    wire N__5042;
    wire N__5039;
    wire N__5038;
    wire N__5037;
    wire N__5032;
    wire N__5029;
    wire N__5024;
    wire N__5021;
    wire N__5018;
    wire N__5015;
    wire N__5012;
    wire N__5009;
    wire N__5008;
    wire N__5005;
    wire N__5004;
    wire N__5001;
    wire N__4998;
    wire N__4995;
    wire N__4992;
    wire N__4987;
    wire N__4984;
    wire N__4981;
    wire N__4978;
    wire N__4975;
    wire N__4970;
    wire N__4969;
    wire N__4968;
    wire N__4967;
    wire N__4966;
    wire N__4965;
    wire N__4962;
    wire N__4959;
    wire N__4956;
    wire N__4953;
    wire N__4950;
    wire N__4947;
    wire N__4944;
    wire N__4939;
    wire N__4936;
    wire N__4933;
    wire N__4930;
    wire N__4927;
    wire N__4924;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4908;
    wire N__4905;
    wire N__4900;
    wire N__4897;
    wire N__4894;
    wire N__4891;
    wire N__4888;
    wire N__4883;
    wire N__4882;
    wire N__4879;
    wire N__4876;
    wire N__4871;
    wire N__4868;
    wire N__4867;
    wire N__4864;
    wire N__4861;
    wire N__4860;
    wire N__4857;
    wire N__4854;
    wire N__4851;
    wire N__4846;
    wire N__4843;
    wire N__4840;
    wire N__4837;
    wire N__4832;
    wire N__4829;
    wire N__4826;
    wire N__4825;
    wire N__4822;
    wire N__4819;
    wire N__4818;
    wire N__4815;
    wire N__4812;
    wire N__4809;
    wire N__4802;
    wire N__4799;
    wire N__4796;
    wire N__4793;
    wire N__4790;
    wire N__4787;
    wire N__4784;
    wire N__4781;
    wire N__4778;
    wire N__4777;
    wire N__4774;
    wire N__4771;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4756;
    wire N__4755;
    wire N__4754;
    wire N__4753;
    wire N__4752;
    wire N__4751;
    wire N__4742;
    wire N__4735;
    wire N__4730;
    wire N__4727;
    wire N__4724;
    wire N__4721;
    wire N__4720;
    wire N__4719;
    wire N__4718;
    wire N__4717;
    wire N__4716;
    wire N__4715;
    wire N__4714;
    wire N__4711;
    wire N__4708;
    wire N__4699;
    wire N__4692;
    wire N__4685;
    wire N__4682;
    wire N__4681;
    wire N__4680;
    wire N__4679;
    wire N__4678;
    wire N__4677;
    wire N__4668;
    wire N__4663;
    wire N__4658;
    wire N__4655;
    wire N__4652;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4642;
    wire N__4641;
    wire N__4638;
    wire N__4635;
    wire N__4632;
    wire N__4625;
    wire N__4624;
    wire N__4623;
    wire N__4622;
    wire N__4613;
    wire N__4610;
    wire N__4607;
    wire N__4606;
    wire N__4603;
    wire N__4602;
    wire N__4599;
    wire N__4598;
    wire N__4593;
    wire N__4588;
    wire N__4583;
    wire N__4582;
    wire N__4581;
    wire N__4580;
    wire N__4577;
    wire N__4572;
    wire N__4569;
    wire N__4562;
    wire N__4561;
    wire N__4560;
    wire N__4559;
    wire N__4554;
    wire N__4549;
    wire N__4544;
    wire N__4543;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4523;
    wire N__4520;
    wire N__4517;
    wire N__4514;
    wire N__4511;
    wire N__4508;
    wire N__4507;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4492;
    wire N__4491;
    wire N__4488;
    wire N__4483;
    wire N__4480;
    wire N__4479;
    wire N__4476;
    wire N__4473;
    wire N__4470;
    wire N__4467;
    wire N__4460;
    wire N__4459;
    wire N__4458;
    wire N__4457;
    wire N__4452;
    wire N__4447;
    wire N__4442;
    wire N__4439;
    wire N__4438;
    wire N__4437;
    wire N__4434;
    wire N__4431;
    wire N__4428;
    wire N__4421;
    wire N__4420;
    wire N__4417;
    wire N__4414;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4400;
    wire N__4397;
    wire N__4394;
    wire N__4391;
    wire N__4388;
    wire N__4385;
    wire N__4384;
    wire N__4381;
    wire N__4378;
    wire N__4373;
    wire N__4372;
    wire N__4371;
    wire N__4368;
    wire N__4361;
    wire N__4358;
    wire N__4357;
    wire N__4356;
    wire N__4349;
    wire N__4346;
    wire N__4343;
    wire N__4340;
    wire N__4337;
    wire N__4334;
    wire N__4331;
    wire N__4330;
    wire N__4327;
    wire N__4324;
    wire N__4319;
    wire N__4318;
    wire N__4317;
    wire N__4316;
    wire N__4315;
    wire N__4312;
    wire N__4309;
    wire N__4308;
    wire N__4307;
    wire N__4306;
    wire N__4303;
    wire N__4300;
    wire N__4291;
    wire N__4286;
    wire N__4277;
    wire N__4276;
    wire N__4275;
    wire N__4274;
    wire N__4273;
    wire N__4272;
    wire N__4271;
    wire N__4270;
    wire N__4267;
    wire N__4264;
    wire N__4255;
    wire N__4250;
    wire N__4241;
    wire N__4240;
    wire N__4237;
    wire N__4234;
    wire N__4233;
    wire N__4232;
    wire N__4231;
    wire N__4230;
    wire N__4229;
    wire N__4228;
    wire N__4225;
    wire N__4222;
    wire N__4215;
    wire N__4208;
    wire N__4199;
    wire N__4196;
    wire N__4193;
    wire N__4190;
    wire N__4189;
    wire N__4186;
    wire N__4183;
    wire N__4180;
    wire N__4175;
    wire N__4174;
    wire N__4173;
    wire N__4172;
    wire N__4171;
    wire N__4170;
    wire N__4169;
    wire N__4168;
    wire N__4167;
    wire N__4166;
    wire N__4165;
    wire N__4142;
    wire N__4139;
    wire N__4136;
    wire N__4135;
    wire N__4130;
    wire N__4127;
    wire N__4126;
    wire N__4125;
    wire N__4118;
    wire N__4115;
    wire N__4112;
    wire N__4109;
    wire N__4106;
    wire N__4103;
    wire N__4100;
    wire N__4097;
    wire N__4096;
    wire N__4093;
    wire N__4090;
    wire N__4085;
    wire N__4082;
    wire N__4079;
    wire N__4076;
    wire N__4073;
    wire N__4070;
    wire N__4069;
    wire N__4068;
    wire N__4067;
    wire N__4066;
    wire N__4063;
    wire N__4054;
    wire N__4049;
    wire N__4048;
    wire N__4047;
    wire N__4044;
    wire N__4041;
    wire N__4040;
    wire N__4037;
    wire N__4032;
    wire N__4029;
    wire N__4026;
    wire N__4021;
    wire N__4016;
    wire N__4013;
    wire N__4012;
    wire N__4009;
    wire N__4006;
    wire N__4001;
    wire N__4000;
    wire N__3997;
    wire N__3994;
    wire N__3989;
    wire N__3986;
    wire N__3983;
    wire N__3980;
    wire N__3979;
    wire N__3976;
    wire N__3973;
    wire N__3968;
    wire N__3965;
    wire N__3962;
    wire N__3961;
    wire N__3958;
    wire N__3955;
    wire N__3950;
    wire N__3947;
    wire N__3944;
    wire N__3941;
    wire N__3940;
    wire N__3937;
    wire N__3934;
    wire N__3929;
    wire N__3926;
    wire N__3925;
    wire N__3922;
    wire N__3919;
    wire N__3914;
    wire N__3913;
    wire N__3910;
    wire N__3907;
    wire N__3902;
    wire N__3899;
    wire N__3898;
    wire N__3895;
    wire N__3892;
    wire N__3887;
    wire N__3884;
    wire N__3883;
    wire N__3882;
    wire N__3881;
    wire N__3878;
    wire N__3871;
    wire N__3868;
    wire N__3863;
    wire N__3862;
    wire N__3859;
    wire N__3856;
    wire N__3851;
    wire N__3848;
    wire N__3847;
    wire N__3844;
    wire N__3841;
    wire N__3836;
    wire N__3833;
    wire N__3830;
    wire N__3827;
    wire N__3826;
    wire N__3823;
    wire N__3820;
    wire N__3815;
    wire N__3814;
    wire N__3811;
    wire N__3808;
    wire N__3803;
    wire N__3802;
    wire N__3799;
    wire N__3796;
    wire N__3791;
    wire N__3790;
    wire N__3787;
    wire N__3782;
    wire N__3781;
    wire N__3778;
    wire N__3775;
    wire N__3770;
    wire N__3769;
    wire N__3766;
    wire N__3763;
    wire N__3758;
    wire N__3755;
    wire N__3752;
    wire N__3749;
    wire N__3746;
    wire N__3743;
    wire N__3740;
    wire N__3737;
    wire N__3736;
    wire N__3731;
    wire N__3728;
    wire N__3725;
    wire N__3722;
    wire N__3721;
    wire N__3720;
    wire N__3717;
    wire N__3712;
    wire N__3707;
    wire N__3706;
    wire N__3701;
    wire N__3698;
    wire N__3697;
    wire N__3694;
    wire N__3691;
    wire N__3686;
    wire N__3683;
    wire N__3682;
    wire N__3679;
    wire N__3676;
    wire N__3671;
    wire N__3670;
    wire N__3667;
    wire N__3664;
    wire N__3659;
    wire N__3656;
    wire N__3653;
    wire N__3650;
    wire N__3647;
    wire N__3644;
    wire N__3641;
    wire N__3638;
    wire N__3635;
    wire N__3632;
    wire N__3631;
    wire N__3630;
    wire N__3629;
    wire N__3624;
    wire N__3619;
    wire N__3614;
    wire N__3613;
    wire N__3612;
    wire N__3611;
    wire N__3610;
    wire N__3599;
    wire N__3596;
    wire N__3595;
    wire N__3590;
    wire N__3587;
    wire N__3584;
    wire N__3581;
    wire N__3578;
    wire N__3575;
    wire N__3572;
    wire N__3571;
    wire N__3568;
    wire N__3565;
    wire N__3560;
    wire N__3557;
    wire N__3554;
    wire N__3551;
    wire N__3550;
    wire N__3547;
    wire N__3544;
    wire N__3539;
    wire N__3538;
    wire N__3535;
    wire N__3532;
    wire N__3527;
    wire N__3524;
    wire N__3521;
    wire N__3518;
    wire N__3515;
    wire N__3512;
    wire N__3509;
    wire N__3506;
    wire N__3505;
    wire N__3502;
    wire N__3499;
    wire N__3494;
    wire N__3493;
    wire N__3490;
    wire N__3487;
    wire N__3482;
    wire N__3481;
    wire N__3478;
    wire N__3475;
    wire N__3470;
    wire N__3467;
    wire N__3466;
    wire N__3463;
    wire N__3460;
    wire N__3455;
    wire N__3454;
    wire N__3451;
    wire N__3448;
    wire N__3443;
    wire N__3442;
    wire N__3441;
    wire N__3434;
    wire N__3433;
    wire N__3432;
    wire N__3431;
    wire N__3430;
    wire N__3427;
    wire N__3420;
    wire N__3417;
    wire N__3410;
    wire N__3409;
    wire N__3408;
    wire N__3407;
    wire N__3406;
    wire N__3405;
    wire N__3404;
    wire N__3395;
    wire N__3392;
    wire N__3387;
    wire N__3380;
    wire N__3379;
    wire N__3378;
    wire N__3375;
    wire N__3374;
    wire N__3373;
    wire N__3372;
    wire N__3371;
    wire N__3368;
    wire N__3365;
    wire N__3362;
    wire N__3355;
    wire N__3348;
    wire N__3341;
    wire N__3338;
    wire N__3335;
    wire N__3332;
    wire N__3331;
    wire N__3328;
    wire N__3325;
    wire N__3320;
    wire N__3317;
    wire N__3314;
    wire N__3311;
    wire N__3308;
    wire N__3305;
    wire N__3302;
    wire N__3299;
    wire N__3296;
    wire N__3293;
    wire N__3290;
    wire N__3287;
    wire N__3284;
    wire N__3281;
    wire N__3278;
    wire N__3275;
    wire N__3272;
    wire N__3269;
    wire N__3266;
    wire N__3263;
    wire N__3260;
    wire N__3257;
    wire N__3254;
    wire N__3251;
    wire N__3248;
    wire N__3245;
    wire N__3242;
    wire N__3239;
    wire N__3236;
    wire N__3233;
    wire N__3230;
    wire N__3227;
    wire N__3224;
    wire N__3221;
    wire N__3218;
    wire N__3215;
    wire N__3212;
    wire N__3209;
    wire N__3206;
    wire N__3203;
    wire N__3200;
    wire N__3197;
    wire N__3194;
    wire N__3191;
    wire N__3190;
    wire N__3187;
    wire N__3184;
    wire N__3179;
    wire N__3176;
    wire N__3173;
    wire N__3172;
    wire N__3169;
    wire N__3166;
    wire N__3161;
    wire N__3158;
    wire N__3155;
    wire N__3152;
    wire N__3149;
    wire N__3146;
    wire N__3143;
    wire N__3142;
    wire N__3139;
    wire N__3136;
    wire N__3133;
    wire N__3128;
    wire N__3125;
    wire N__3124;
    wire N__3121;
    wire N__3118;
    wire N__3113;
    wire N__3110;
    wire N__3107;
    wire N__3104;
    wire N__3101;
    wire N__3098;
    wire N__3095;
    wire N__3092;
    wire N__3089;
    wire N__3088;
    wire N__3085;
    wire N__3082;
    wire N__3081;
    wire N__3076;
    wire N__3073;
    wire N__3068;
    wire N__3067;
    wire N__3066;
    wire N__3065;
    wire N__3062;
    wire N__3055;
    wire N__3052;
    wire N__3047;
    wire N__3046;
    wire N__3043;
    wire N__3040;
    wire N__3035;
    wire N__3032;
    wire N__3031;
    wire N__3028;
    wire N__3025;
    wire N__3020;
    wire N__3017;
    wire N__3016;
    wire N__3013;
    wire N__3010;
    wire N__3005;
    wire N__3002;
    wire N__2999;
    wire N__2996;
    wire N__2995;
    wire N__2992;
    wire N__2989;
    wire N__2984;
    wire N__2981;
    wire N__2978;
    wire N__2975;
    wire N__2972;
    wire N__2969;
    wire N__2966;
    wire N__2965;
    wire N__2962;
    wire N__2959;
    wire N__2954;
    wire N__2953;
    wire N__2952;
    wire N__2951;
    wire N__2950;
    wire N__2949;
    wire N__2944;
    wire N__2941;
    wire N__2936;
    wire N__2933;
    wire N__2928;
    wire N__2925;
    wire N__2922;
    wire N__2919;
    wire N__2916;
    wire N__2913;
    wire N__2910;
    wire N__2907;
    wire N__2904;
    wire N__2897;
    wire N__2894;
    wire N__2891;
    wire N__2888;
    wire N__2885;
    wire N__2882;
    wire N__2879;
    wire N__2876;
    wire N__2873;
    wire N__2870;
    wire N__2867;
    wire N__2864;
    wire N__2861;
    wire N__2858;
    wire N__2855;
    wire N__2852;
    wire N__2851;
    wire N__2846;
    wire N__2843;
    wire N__2840;
    wire N__2837;
    wire N__2834;
    wire N__2831;
    wire N__2828;
    wire N__2827;
    wire N__2822;
    wire N__2819;
    wire N__2816;
    wire N__2813;
    wire N__2810;
    wire N__2809;
    wire N__2804;
    wire N__2801;
    wire N__2798;
    wire N__2795;
    wire N__2792;
    wire N__2789;
    wire N__2786;
    wire N__2785;
    wire N__2784;
    wire N__2783;
    wire N__2780;
    wire N__2773;
    wire N__2770;
    wire N__2767;
    wire N__2764;
    wire N__2761;
    wire N__2758;
    wire N__2753;
    wire N__2750;
    wire N__2747;
    wire N__2746;
    wire N__2745;
    wire N__2742;
    wire N__2737;
    wire N__2732;
    wire N__2729;
    wire N__2726;
    wire N__2725;
    wire N__2720;
    wire N__2717;
    wire N__2714;
    wire N__2711;
    wire N__2710;
    wire N__2709;
    wire N__2706;
    wire N__2701;
    wire N__2698;
    wire N__2695;
    wire N__2692;
    wire N__2689;
    wire N__2686;
    wire N__2683;
    wire N__2680;
    wire N__2677;
    wire N__2674;
    wire N__2671;
    wire N__2666;
    wire N__2665;
    wire N__2664;
    wire N__2661;
    wire N__2660;
    wire N__2657;
    wire N__2656;
    wire N__2653;
    wire N__2644;
    wire N__2641;
    wire N__2636;
    wire N__2633;
    wire N__2630;
    wire N__2627;
    wire N__2624;
    wire N__2621;
    wire N__2618;
    wire N__2615;
    wire N__2612;
    wire N__2609;
    wire N__2606;
    wire N__2603;
    wire N__2600;
    wire N__2597;
    wire N__2594;
    wire N__2593;
    wire N__2588;
    wire N__2585;
    wire N__2582;
    wire N__2579;
    wire N__2576;
    wire N__2575;
    wire N__2572;
    wire N__2567;
    wire N__2564;
    wire N__2561;
    wire N__2558;
    wire N__2555;
    wire N__2552;
    wire N__2549;
    wire N__2548;
    wire N__2543;
    wire N__2540;
    wire N__2537;
    wire N__2534;
    wire N__2531;
    wire N__2528;
    wire N__2525;
    wire N__2522;
    wire N__2519;
    wire N__2516;
    wire N__2515;
    wire N__2512;
    wire N__2509;
    wire N__2506;
    wire N__2503;
    wire N__2498;
    wire N__2495;
    wire N__2492;
    wire N__2489;
    wire N__2488;
    wire N__2483;
    wire N__2480;
    wire N__2477;
    wire N__2474;
    wire N__2471;
    wire N__2468;
    wire N__2467;
    wire N__2462;
    wire N__2459;
    wire N__2456;
    wire N__2453;
    wire N__2450;
    wire N__2449;
    wire N__2446;
    wire N__2443;
    wire N__2440;
    wire N__2435;
    wire N__2432;
    wire N__2429;
    wire N__2426;
    wire N__2423;
    wire N__2422;
    wire N__2417;
    wire N__2414;
    wire N__2411;
    wire N__2408;
    wire N__2405;
    wire N__2402;
    wire N__2399;
    wire N__2398;
    wire N__2397;
    wire N__2396;
    wire N__2395;
    wire N__2394;
    wire N__2393;
    wire N__2392;
    wire N__2391;
    wire N__2390;
    wire N__2369;
    wire CLK80_OUT;
    wire GNDG0;
    wire VCCG0;
    wire A_c_18;
    wire A_c_16;
    wire A_c_17;
    wire \U409_CIA.g0Z0Z_11_cascade_ ;
    wire \U409_CIA.g0Z0Z_8 ;
    wire A_c_25;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_ ;
    wire A_c_27;
    wire A_c_24;
    wire A_c_26;
    wire A_c_28;
    wire \U409_CIA.g0Z0Z_10_cascade_ ;
    wire A_c_29;
    wire \U409_CIA.g0Z0Z_2 ;
    wire A_c_31;
    wire A_c_30;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3 ;
    wire A_c_21;
    wire A_c_20;
    wire \U409_ADDRESS_DECODE.CIA_SPACEm_6 ;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2_cascade_ ;
    wire A_c_19;
    wire A_c_22;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2 ;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3 ;
    wire PORTSIZE_0_i;
    wire \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3 ;
    wire A_c_23;
    wire U409_ADDRESS_DECODE_un1_nREGSPACE_i;
    wire \U409_ADDRESS_DECODE.un10_ROMENZ0 ;
    wire \U409_TICK.TICK603_8 ;
    wire \U409_TICK.TICK603_11_cascade_ ;
    wire \U409_TICK.TICK603_14_cascade_ ;
    wire \U409_TICK.COUNTER60Z0Z_1 ;
    wire \U409_TICK.COUNTER60Z0Z_0 ;
    wire bfn_8_8_0_;
    wire \U409_TICK.COUNTER60Z0Z_2 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_1 ;
    wire \U409_TICK.COUNTER60Z0Z_3 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_2 ;
    wire \U409_TICK.COUNTER60Z0Z_4 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_4 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_3 ;
    wire \U409_TICK.COUNTER60Z0Z_5 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_4 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_6 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_5 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_6 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_8 ;
    wire bfn_8_9_0_;
    wire \U409_TICK.un3_COUNTER60_1_cry_9 ;
    wire \U409_TICK.COUNTER60Z0Z_11 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_10 ;
    wire \U409_TICK.COUNTER60Z0Z_12 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_11 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_12 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_13 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_15 ;
    wire \U409_TICK.COUNTER60Z0Z_16 ;
    wire \U409_ADDRESS_DECODE.un1_nREGSPACEZ0 ;
    wire nBUFEN_c;
    wire A_c_13;
    wire U409_ADDRESS_DECODE_un1_nCIACS1_i;
    wire A_c_12;
    wire U409_ADDRESS_DECODE_un1_nCIACS0_i;
    wire bfn_9_5_0_;
    wire \U409_TICK.un2_COUNTER50_1_cry_1 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_3 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_4 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_5 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_6 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_8 ;
    wire bfn_9_6_0_;
    wire \U409_TICK.un2_COUNTER50_1_cry_9 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_10 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_11 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_12 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_13 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_15 ;
    wire TICK60_c;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_9 ;
    wire \U409_TICK.COUNTER60Z0Z_9 ;
    wire \U409_TICK.COUNTER60Z0Z_6 ;
    wire \U409_TICK.TICK603_9_cascade_ ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_15 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_8 ;
    wire \U409_TICK.COUNTER60Z0Z_8 ;
    wire \U409_TICK.COUNTER60Z0Z_13 ;
    wire \U409_TICK.COUNTER60Z0Z_10 ;
    wire \U409_TICK.COUNTER60Z0Z_7 ;
    wire \U409_TICK.COUNTER60Z0Z_15 ;
    wire \U409_TICK.TICK603_10 ;
    wire \U409_TICK.TICK603_14 ;
    wire \U409_TICK.TICK603_9 ;
    wire \U409_TICK.TICK603_10_cascade_ ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_14 ;
    wire \U409_TICK.COUNTER60Z0Z_14 ;
    wire CIA_ENABLEm;
    wire \U409_CIA.CIA_HOLDZ0 ;
    wire \U409_CIA.g0Z0Z_14 ;
    wire \U409_CIA.g0Z0Z_13 ;
    wire \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ;
    wire \U409_TRANSFER_ACK.RESETn_c_i ;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_3_0_cascade_ ;
    wire \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa_cascade_ ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0 ;
    wire \U409_TICK.COUNTER50Z0Z_3 ;
    wire \U409_TICK.COUNTER50Z0Z_12 ;
    wire \U409_TICK.TICK503_8_cascade_ ;
    wire \U409_TICK.COUNTER50Z0Z_10 ;
    wire \U409_TICK.TICK503_14_cascade_ ;
    wire \U409_TICK.COUNTER50Z0Z_0 ;
    wire \U409_TICK.COUNTER50Z0Z_4 ;
    wire \U409_TICK.COUNTER50Z0Z_7 ;
    wire \U409_TICK.TICK503_10_cascade_ ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_5 ;
    wire \U409_TICK.COUNTER50Z0Z_5 ;
    wire \U409_TICK.COUNTER50Z0Z_8 ;
    wire \U409_TICK.COUNTER50Z0Z_2 ;
    wire \U409_TICK.COUNTER50Z0Z_1 ;
    wire \U409_TICK.COUNTER50Z0Z_16 ;
    wire \U409_TICK.TICK503_11 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_6 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_13 ;
    wire \U409_TICK.COUNTER50Z0Z_6 ;
    wire \U409_TICK.COUNTER50Z0Z_13 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_11 ;
    wire \U409_TICK.TICK503_9_cascade_ ;
    wire \U409_TICK.COUNTER50Z0Z_11 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_14 ;
    wire \U409_TICK.COUNTER50Z0Z_14 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_15 ;
    wire \U409_TICK.COUNTER50Z0Z_15 ;
    wire \INVU409_TRANSFER_ACK.LASTCLK_0C_net ;
    wire \U409_TRANSFER_ACK.N_97_cascade_ ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_1 ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_0 ;
    wire \U409_TRANSFER_ACK.N_4_cascade_ ;
    wire \U409_TRANSFER_ACK.N_97 ;
    wire \U409_TRANSFER_ACK.CIA_TACK_EN_0_cascade_ ;
    wire \U409_TRANSFER_ACK.i6_mux_0 ;
    wire \INVU409_TRANSFER_ACK.LASTCLK_1C_net ;
    wire \U409_TRANSFER_ACK.CIA_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.N_4 ;
    wire \U409_TRANSFER_ACK.m9_bm ;
    wire \U409_TRANSFER_ACK.m9_am_cascade_ ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_0C_net ;
    wire \U409_TRANSFER_ACK.ROM_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER5_0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_ ;
    wire TACK_OUTn;
    wire \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ;
    wire TICK50_c;
    wire \U409_TICK.TICK503_10 ;
    wire \U409_TICK.TICK503_14 ;
    wire \U409_TICK.TICK503_9 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_9 ;
    wire \U409_TICK.COUNTER50Z0Z_9 ;
    wire CLK6_c_g;
    wire bfn_11_7_0_;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_1 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_3 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4 ;
    wire \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_ ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ;
    wire \U409_CIA.CIA_CLK_COUNT11_0_a2_2 ;
    wire \U409_CIA.N_9_cascade_ ;
    wire \U409_CIA.VMAZ0 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_3 ;
    wire \U409_CIA.N_20_cascade_ ;
    wire \U409_CIA.CLKCIA6_0_a2_1 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_0 ;
    wire \U409_CIA.CLKCIAZ0_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_1 ;
    wire CLKCIA_c;
    wire CLK28_IN_c_g;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_5 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_4 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_2 ;
    wire \U409_CIA.CLKCIA8_0_a2_0 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ;
    wire TSn_c;
    wire CLK40_IN_c;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ;
    wire OVL_c;
    wire \U409_ADDRESS_DECODE.un6_ROMENZ0 ;
    wire U409_ADDRESS_DECODE_un1_nRAMSPACE_i;
    wire \U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ;
    wire \INVU409_TRANSFER_ACK.TACK_EN_iC_net ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0 ;
    wire U409_ADDRESS_DECODE_Z2_SPACE;
    wire U409_ADDRESS_DECODE_un1_ROMEN_0;
    wire ROMENm_i;
    wire CONSTANT_ONE_NET;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0 ;
    wire RESETn_c;
    wire TACKn_in;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ;
    wire TACK_EN_i;
    wire N_347_i;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="SIMPLE";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0001111;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE pll (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__4970),
            .RESETB(N__5222),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(CLK80_OUT));
    PRE_IO_GBUF CLK28_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__6034),
            .GLOBALBUFFEROUTPUT(CLK28_IN_c_g));
    IO_PAD CLK28_IN_ibuf_gb_io_iopad (
            .OE(N__6036),
            .DIN(N__6035),
            .DOUT(N__6034),
            .PACKAGEPIN(CLK28_IN));
    defparam CLK28_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK28_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK28_IN_ibuf_gb_io_preio (
            .PADOEN(N__6036),
            .PADOUT(N__6035),
            .PADIN(N__6034),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK6_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__6024),
            .GLOBALBUFFEROUTPUT(CLK6_c_g));
    IO_PAD CLK6_ibuf_gb_io_iopad (
            .OE(N__6026),
            .DIN(N__6025),
            .DOUT(N__6024),
            .PACKAGEPIN(CLK6));
    defparam CLK6_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK6_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK6_ibuf_gb_io_preio (
            .PADOEN(N__6026),
            .PADOUT(N__6025),
            .PADIN(N__6024),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKCIA_obuf_iopad (
            .OE(N__6015),
            .DIN(N__6014),
            .DOUT(N__6013),
            .PACKAGEPIN(CLKCIA));
    defparam CLKCIA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKCIA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKCIA_obuf_preio (
            .PADOEN(N__6015),
            .PADOUT(N__6014),
            .PADIN(N__6013),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4658),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_23_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_23_iopad (
            .OE(N__6006),
            .DIN(N__6005),
            .DOUT(N__6004),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__6006),
            .PADOUT(N__6005),
            .PADIN(N__6004),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_24_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_24_iopad (
            .OE(N__5997),
            .DIN(N__5996),
            .DOUT(N__5995),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__5997),
            .PADOUT(N__5996),
            .PADIN(N__5995),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nCIACS0_obuf_iopad (
            .OE(N__5988),
            .DIN(N__5987),
            .DOUT(N__5986),
            .PACKAGEPIN(nCIACS0));
    defparam nCIACS0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nCIACS0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nCIACS0_obuf_preio (
            .PADOEN(N__5988),
            .PADOUT(N__5987),
            .PADIN(N__5986),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3239),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nCIACS1_obuf_iopad (
            .OE(N__5979),
            .DIN(N__5978),
            .DOUT(N__5977),
            .PACKAGEPIN(nCIACS1));
    defparam nCIACS1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nCIACS1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nCIACS1_obuf_preio (
            .PADOEN(N__5979),
            .PADOUT(N__5978),
            .PADIN(N__5977),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3275),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_31_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_31_iopad (
            .OE(N__5970),
            .DIN(N__5969),
            .DOUT(N__5968),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__5970),
            .PADOUT(N__5969),
            .PADIN(N__5968),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_17_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_17_iopad (
            .OE(N__5961),
            .DIN(N__5960),
            .DOUT(N__5959),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__5961),
            .PADOUT(N__5960),
            .PADIN(N__5959),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_21_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_21_iopad (
            .OE(N__5952),
            .DIN(N__5951),
            .DOUT(N__5950),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__5952),
            .PADOUT(N__5951),
            .PADIN(N__5950),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TACKn_iobuf_iopad.PULLUP=1'b1;
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__5943),
            .DIN(N__5942),
            .DOUT(N__5941),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__5943),
            .PADOUT(N__5942),
            .PADIN(N__5941),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5372),
            .DIN0(TACKn_in),
            .DOUT0(N__4400),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_12_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_12_iopad (
            .OE(N__5934),
            .DIN(N__5933),
            .DOUT(N__5932),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__5934),
            .PADOUT(N__5933),
            .PADIN(N__5932),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__5925),
            .DIN(N__5924),
            .DOUT(N__5923),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__5925),
            .PADOUT(N__5924),
            .PADIN(N__5923),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam PORTSIZE_obuf_iopad.PULLUP=1'b1;
    IO_PAD PORTSIZE_obuf_iopad (
            .OE(N__5916),
            .DIN(N__5915),
            .DOUT(N__5914),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PORTSIZE_obuf_preio (
            .PADOEN(N__5916),
            .PADOUT(N__5915),
            .PADIN(N__5914),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2618),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nRAMSPACE_obuf_iopad (
            .OE(N__5907),
            .DIN(N__5906),
            .DOUT(N__5905),
            .PACKAGEPIN(nRAMSPACE));
    defparam nRAMSPACE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nRAMSPACE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nRAMSPACE_obuf_preio (
            .PADOEN(N__5907),
            .PADOUT(N__5906),
            .PADIN(N__5905),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4799),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nROMEN_obuf_iopad (
            .OE(N__5898),
            .DIN(N__5897),
            .DOUT(N__5896),
            .PACKAGEPIN(nROMEN));
    defparam nROMEN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nROMEN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nROMEN_obuf_preio (
            .PADOEN(N__5898),
            .PADOUT(N__5897),
            .PADIN(N__5896),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5243),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_18_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_18_iopad (
            .OE(N__5889),
            .DIN(N__5888),
            .DOUT(N__5887),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__5889),
            .PADOUT(N__5888),
            .PADIN(N__5887),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_29_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_29_iopad (
            .OE(N__5880),
            .DIN(N__5879),
            .DOUT(N__5878),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__5880),
            .PADOUT(N__5879),
            .PADIN(N__5878),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nBUFEN_obuf_iopad (
            .OE(N__5871),
            .DIN(N__5870),
            .DOUT(N__5869),
            .PACKAGEPIN(nBUFEN));
    defparam nBUFEN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nBUFEN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nBUFEN_obuf_preio (
            .PADOEN(N__5871),
            .PADOUT(N__5870),
            .PADIN(N__5869),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3113),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_22_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_22_iopad (
            .OE(N__5862),
            .DIN(N__5861),
            .DOUT(N__5860),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__5862),
            .PADOUT(N__5861),
            .PADIN(N__5860),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_27_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_27_iopad (
            .OE(N__5853),
            .DIN(N__5852),
            .DOUT(N__5851),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__5853),
            .PADOUT(N__5852),
            .PADIN(N__5851),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__5844),
            .DIN(N__5843),
            .DOUT(N__5842),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__5844),
            .PADOUT(N__5843),
            .PADIN(N__5842),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__5835),
            .DIN(N__5834),
            .DOUT(N__5833),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__5835),
            .PADOUT(N__5834),
            .PADIN(N__5833),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_20_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_20_iopad (
            .OE(N__5826),
            .DIN(N__5825),
            .DOUT(N__5824),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__5826),
            .PADOUT(N__5825),
            .PADIN(N__5824),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_13_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_13_iopad (
            .OE(N__5817),
            .DIN(N__5816),
            .DOUT(N__5815),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__5817),
            .PADOUT(N__5816),
            .PADIN(N__5815),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_25_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_25_iopad (
            .OE(N__5808),
            .DIN(N__5807),
            .DOUT(N__5806),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__5808),
            .PADOUT(N__5807),
            .PADIN(N__5806),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nREGSPACE_obuf_iopad (
            .OE(N__5799),
            .DIN(N__5798),
            .DOUT(N__5797),
            .PACKAGEPIN(nREGSPACE));
    defparam nREGSPACE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nREGSPACE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nREGSPACE_obuf_preio (
            .PADOEN(N__5799),
            .PADOUT(N__5798),
            .PADIN(N__5797),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2897),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK50_obuf_iopad (
            .OE(N__5790),
            .DIN(N__5789),
            .DOUT(N__5788),
            .PACKAGEPIN(TICK50));
    defparam TICK50_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK50_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK50_obuf_preio (
            .PADOEN(N__5790),
            .PADOUT(N__5789),
            .PADIN(N__5788),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4346),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_19_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_19_iopad (
            .OE(N__5781),
            .DIN(N__5780),
            .DOUT(N__5779),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__5781),
            .PADOUT(N__5780),
            .PADIN(N__5779),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_28_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_28_iopad (
            .OE(N__5772),
            .DIN(N__5771),
            .DOUT(N__5770),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__5772),
            .PADOUT(N__5771),
            .PADIN(N__5770),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_30_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_30_iopad (
            .OE(N__5763),
            .DIN(N__5762),
            .DOUT(N__5761),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__5763),
            .PADOUT(N__5762),
            .PADIN(N__5761),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD OVL_ibuf_iopad (
            .OE(N__5754),
            .DIN(N__5753),
            .DOUT(N__5752),
            .PACKAGEPIN(OVL));
    defparam OVL_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam OVL_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO OVL_ibuf_preio (
            .PADOEN(N__5754),
            .PADOUT(N__5753),
            .PADIN(N__5752),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(OVL_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_16_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_16_iopad (
            .OE(N__5745),
            .DIN(N__5744),
            .DOUT(N__5743),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__5745),
            .PADOUT(N__5744),
            .PADIN(N__5743),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK60_obuf_iopad (
            .OE(N__5736),
            .DIN(N__5735),
            .DOUT(N__5734),
            .PACKAGEPIN(TICK60));
    defparam TICK60_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK60_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK60_obuf_preio (
            .PADOEN(N__5736),
            .PADOUT(N__5735),
            .PADIN(N__5734),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3587),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_26_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_26_iopad (
            .OE(N__5727),
            .DIN(N__5726),
            .DOUT(N__5725),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__5727),
            .PADOUT(N__5726),
            .PADIN(N__5725),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1319 (
            .O(N__5708),
            .I(N__5702));
    InMux I__1318 (
            .O(N__5707),
            .I(N__5702));
    LocalMux I__1317 (
            .O(N__5702),
            .I(N__5699));
    Odrv4 I__1316 (
            .O(N__5699),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ));
    InMux I__1315 (
            .O(N__5696),
            .I(N__5689));
    InMux I__1314 (
            .O(N__5695),
            .I(N__5684));
    InMux I__1313 (
            .O(N__5694),
            .I(N__5684));
    InMux I__1312 (
            .O(N__5693),
            .I(N__5679));
    InMux I__1311 (
            .O(N__5692),
            .I(N__5679));
    LocalMux I__1310 (
            .O(N__5689),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1309 (
            .O(N__5684),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1308 (
            .O(N__5679),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    InMux I__1307 (
            .O(N__5672),
            .I(N__5661));
    InMux I__1306 (
            .O(N__5671),
            .I(N__5661));
    InMux I__1305 (
            .O(N__5670),
            .I(N__5658));
    InMux I__1304 (
            .O(N__5669),
            .I(N__5649));
    InMux I__1303 (
            .O(N__5668),
            .I(N__5649));
    InMux I__1302 (
            .O(N__5667),
            .I(N__5649));
    InMux I__1301 (
            .O(N__5666),
            .I(N__5649));
    LocalMux I__1300 (
            .O(N__5661),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1299 (
            .O(N__5658),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1298 (
            .O(N__5649),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    CascadeMux I__1297 (
            .O(N__5642),
            .I(N__5637));
    InMux I__1296 (
            .O(N__5641),
            .I(N__5633));
    InMux I__1295 (
            .O(N__5640),
            .I(N__5630));
    InMux I__1294 (
            .O(N__5637),
            .I(N__5625));
    InMux I__1293 (
            .O(N__5636),
            .I(N__5625));
    LocalMux I__1292 (
            .O(N__5633),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1291 (
            .O(N__5630),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1290 (
            .O(N__5625),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    InMux I__1289 (
            .O(N__5618),
            .I(N__5615));
    LocalMux I__1288 (
            .O(N__5615),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0 ));
    CascadeMux I__1287 (
            .O(N__5612),
            .I(N__5608));
    InMux I__1286 (
            .O(N__5611),
            .I(N__5605));
    InMux I__1285 (
            .O(N__5608),
            .I(N__5601));
    LocalMux I__1284 (
            .O(N__5605),
            .I(N__5596));
    CascadeMux I__1283 (
            .O(N__5604),
            .I(N__5593));
    LocalMux I__1282 (
            .O(N__5601),
            .I(N__5587));
    CascadeMux I__1281 (
            .O(N__5600),
            .I(N__5584));
    CascadeMux I__1280 (
            .O(N__5599),
            .I(N__5580));
    Span4Mux_v I__1279 (
            .O(N__5596),
            .I(N__5573));
    InMux I__1278 (
            .O(N__5593),
            .I(N__5570));
    InMux I__1277 (
            .O(N__5592),
            .I(N__5563));
    InMux I__1276 (
            .O(N__5591),
            .I(N__5563));
    InMux I__1275 (
            .O(N__5590),
            .I(N__5563));
    Span4Mux_v I__1274 (
            .O(N__5587),
            .I(N__5559));
    InMux I__1273 (
            .O(N__5584),
            .I(N__5554));
    InMux I__1272 (
            .O(N__5583),
            .I(N__5554));
    InMux I__1271 (
            .O(N__5580),
            .I(N__5549));
    InMux I__1270 (
            .O(N__5579),
            .I(N__5549));
    InMux I__1269 (
            .O(N__5578),
            .I(N__5546));
    InMux I__1268 (
            .O(N__5577),
            .I(N__5543));
    CascadeMux I__1267 (
            .O(N__5576),
            .I(N__5538));
    Span4Mux_h I__1266 (
            .O(N__5573),
            .I(N__5532));
    LocalMux I__1265 (
            .O(N__5570),
            .I(N__5527));
    LocalMux I__1264 (
            .O(N__5563),
            .I(N__5527));
    InMux I__1263 (
            .O(N__5562),
            .I(N__5524));
    Span4Mux_h I__1262 (
            .O(N__5559),
            .I(N__5520));
    LocalMux I__1261 (
            .O(N__5554),
            .I(N__5517));
    LocalMux I__1260 (
            .O(N__5549),
            .I(N__5514));
    LocalMux I__1259 (
            .O(N__5546),
            .I(N__5509));
    LocalMux I__1258 (
            .O(N__5543),
            .I(N__5509));
    InMux I__1257 (
            .O(N__5542),
            .I(N__5504));
    InMux I__1256 (
            .O(N__5541),
            .I(N__5504));
    InMux I__1255 (
            .O(N__5538),
            .I(N__5497));
    InMux I__1254 (
            .O(N__5537),
            .I(N__5497));
    InMux I__1253 (
            .O(N__5536),
            .I(N__5497));
    InMux I__1252 (
            .O(N__5535),
            .I(N__5494));
    Span4Mux_h I__1251 (
            .O(N__5532),
            .I(N__5487));
    Span4Mux_v I__1250 (
            .O(N__5527),
            .I(N__5487));
    LocalMux I__1249 (
            .O(N__5524),
            .I(N__5487));
    InMux I__1248 (
            .O(N__5523),
            .I(N__5484));
    Span4Mux_h I__1247 (
            .O(N__5520),
            .I(N__5469));
    Span4Mux_v I__1246 (
            .O(N__5517),
            .I(N__5469));
    Span4Mux_v I__1245 (
            .O(N__5514),
            .I(N__5469));
    Span4Mux_v I__1244 (
            .O(N__5509),
            .I(N__5469));
    LocalMux I__1243 (
            .O(N__5504),
            .I(N__5469));
    LocalMux I__1242 (
            .O(N__5497),
            .I(N__5469));
    LocalMux I__1241 (
            .O(N__5494),
            .I(N__5469));
    Span4Mux_v I__1240 (
            .O(N__5487),
            .I(N__5466));
    LocalMux I__1239 (
            .O(N__5484),
            .I(N__5463));
    Span4Mux_v I__1238 (
            .O(N__5469),
            .I(N__5460));
    Span4Mux_h I__1237 (
            .O(N__5466),
            .I(N__5455));
    Span4Mux_v I__1236 (
            .O(N__5463),
            .I(N__5455));
    Sp12to4 I__1235 (
            .O(N__5460),
            .I(N__5450));
    Sp12to4 I__1234 (
            .O(N__5455),
            .I(N__5450));
    Span12Mux_h I__1233 (
            .O(N__5450),
            .I(N__5447));
    Span12Mux_v I__1232 (
            .O(N__5447),
            .I(N__5444));
    Odrv12 I__1231 (
            .O(N__5444),
            .I(RESETn_c));
    InMux I__1230 (
            .O(N__5441),
            .I(N__5438));
    LocalMux I__1229 (
            .O(N__5438),
            .I(N__5435));
    Span4Mux_v I__1228 (
            .O(N__5435),
            .I(N__5432));
    Sp12to4 I__1227 (
            .O(N__5432),
            .I(N__5429));
    Span12Mux_h I__1226 (
            .O(N__5429),
            .I(N__5426));
    Span12Mux_v I__1225 (
            .O(N__5426),
            .I(N__5423));
    Odrv12 I__1224 (
            .O(N__5423),
            .I(TACKn_in));
    SRMux I__1223 (
            .O(N__5420),
            .I(N__5415));
    SRMux I__1222 (
            .O(N__5419),
            .I(N__5412));
    SRMux I__1221 (
            .O(N__5418),
            .I(N__5409));
    LocalMux I__1220 (
            .O(N__5415),
            .I(N__5406));
    LocalMux I__1219 (
            .O(N__5412),
            .I(N__5403));
    LocalMux I__1218 (
            .O(N__5409),
            .I(N__5400));
    Span12Mux_h I__1217 (
            .O(N__5406),
            .I(N__5397));
    Span4Mux_h I__1216 (
            .O(N__5403),
            .I(N__5394));
    Span4Mux_h I__1215 (
            .O(N__5400),
            .I(N__5391));
    Odrv12 I__1214 (
            .O(N__5397),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    Odrv4 I__1213 (
            .O(N__5394),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    Odrv4 I__1212 (
            .O(N__5391),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    InMux I__1211 (
            .O(N__5384),
            .I(N__5381));
    LocalMux I__1210 (
            .O(N__5381),
            .I(N__5378));
    Span4Mux_v I__1209 (
            .O(N__5378),
            .I(N__5375));
    Odrv4 I__1208 (
            .O(N__5375),
            .I(TACK_EN_i));
    IoInMux I__1207 (
            .O(N__5372),
            .I(N__5369));
    LocalMux I__1206 (
            .O(N__5369),
            .I(N__5366));
    IoSpan4Mux I__1205 (
            .O(N__5366),
            .I(N__5363));
    Sp12to4 I__1204 (
            .O(N__5363),
            .I(N__5360));
    Span12Mux_v I__1203 (
            .O(N__5360),
            .I(N__5357));
    Span12Mux_h I__1202 (
            .O(N__5357),
            .I(N__5354));
    Odrv12 I__1201 (
            .O(N__5354),
            .I(N_347_i));
    InMux I__1200 (
            .O(N__5351),
            .I(N__5346));
    InMux I__1199 (
            .O(N__5350),
            .I(N__5342));
    InMux I__1198 (
            .O(N__5349),
            .I(N__5339));
    LocalMux I__1197 (
            .O(N__5346),
            .I(N__5336));
    InMux I__1196 (
            .O(N__5345),
            .I(N__5332));
    LocalMux I__1195 (
            .O(N__5342),
            .I(N__5327));
    LocalMux I__1194 (
            .O(N__5339),
            .I(N__5327));
    Span4Mux_h I__1193 (
            .O(N__5336),
            .I(N__5323));
    InMux I__1192 (
            .O(N__5335),
            .I(N__5319));
    LocalMux I__1191 (
            .O(N__5332),
            .I(N__5316));
    Span4Mux_h I__1190 (
            .O(N__5327),
            .I(N__5313));
    InMux I__1189 (
            .O(N__5326),
            .I(N__5310));
    Span4Mux_h I__1188 (
            .O(N__5323),
            .I(N__5307));
    InMux I__1187 (
            .O(N__5322),
            .I(N__5304));
    LocalMux I__1186 (
            .O(N__5319),
            .I(N__5301));
    Span4Mux_v I__1185 (
            .O(N__5316),
            .I(N__5298));
    Span4Mux_h I__1184 (
            .O(N__5313),
            .I(N__5293));
    LocalMux I__1183 (
            .O(N__5310),
            .I(N__5293));
    Span4Mux_h I__1182 (
            .O(N__5307),
            .I(N__5288));
    LocalMux I__1181 (
            .O(N__5304),
            .I(N__5288));
    Span12Mux_v I__1180 (
            .O(N__5301),
            .I(N__5285));
    Span4Mux_v I__1179 (
            .O(N__5298),
            .I(N__5282));
    Span4Mux_h I__1178 (
            .O(N__5293),
            .I(N__5279));
    Span4Mux_v I__1177 (
            .O(N__5288),
            .I(N__5276));
    Odrv12 I__1176 (
            .O(N__5285),
            .I(U409_ADDRESS_DECODE_Z2_SPACE));
    Odrv4 I__1175 (
            .O(N__5282),
            .I(U409_ADDRESS_DECODE_Z2_SPACE));
    Odrv4 I__1174 (
            .O(N__5279),
            .I(U409_ADDRESS_DECODE_Z2_SPACE));
    Odrv4 I__1173 (
            .O(N__5276),
            .I(U409_ADDRESS_DECODE_Z2_SPACE));
    InMux I__1172 (
            .O(N__5267),
            .I(N__5263));
    InMux I__1171 (
            .O(N__5266),
            .I(N__5260));
    LocalMux I__1170 (
            .O(N__5263),
            .I(N__5257));
    LocalMux I__1169 (
            .O(N__5260),
            .I(N__5254));
    Span4Mux_v I__1168 (
            .O(N__5257),
            .I(N__5251));
    Span4Mux_v I__1167 (
            .O(N__5254),
            .I(N__5248));
    Odrv4 I__1166 (
            .O(N__5251),
            .I(U409_ADDRESS_DECODE_un1_ROMEN_0));
    Odrv4 I__1165 (
            .O(N__5248),
            .I(U409_ADDRESS_DECODE_un1_ROMEN_0));
    IoInMux I__1164 (
            .O(N__5243),
            .I(N__5240));
    LocalMux I__1163 (
            .O(N__5240),
            .I(N__5237));
    Span4Mux_s1_v I__1162 (
            .O(N__5237),
            .I(N__5234));
    Sp12to4 I__1161 (
            .O(N__5234),
            .I(N__5231));
    Span12Mux_h I__1160 (
            .O(N__5231),
            .I(N__5228));
    Span12Mux_v I__1159 (
            .O(N__5228),
            .I(N__5225));
    Odrv12 I__1158 (
            .O(N__5225),
            .I(ROMENm_i));
    IoInMux I__1157 (
            .O(N__5222),
            .I(N__5219));
    LocalMux I__1156 (
            .O(N__5219),
            .I(N__5216));
    Span4Mux_s2_v I__1155 (
            .O(N__5216),
            .I(N__5213));
    Span4Mux_v I__1154 (
            .O(N__5213),
            .I(N__5210));
    Odrv4 I__1153 (
            .O(N__5210),
            .I(CONSTANT_ONE_NET));
    InMux I__1152 (
            .O(N__5207),
            .I(N__5198));
    InMux I__1151 (
            .O(N__5206),
            .I(N__5198));
    InMux I__1150 (
            .O(N__5205),
            .I(N__5198));
    LocalMux I__1149 (
            .O(N__5198),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ));
    CascadeMux I__1148 (
            .O(N__5195),
            .I(N__5189));
    InMux I__1147 (
            .O(N__5194),
            .I(N__5185));
    InMux I__1146 (
            .O(N__5193),
            .I(N__5178));
    InMux I__1145 (
            .O(N__5192),
            .I(N__5178));
    InMux I__1144 (
            .O(N__5189),
            .I(N__5178));
    InMux I__1143 (
            .O(N__5188),
            .I(N__5175));
    LocalMux I__1142 (
            .O(N__5185),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__1141 (
            .O(N__5178),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__1140 (
            .O(N__5175),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    CascadeMux I__1139 (
            .O(N__5168),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_ ));
    CascadeMux I__1138 (
            .O(N__5165),
            .I(N__5161));
    InMux I__1137 (
            .O(N__5164),
            .I(N__5158));
    InMux I__1136 (
            .O(N__5161),
            .I(N__5155));
    LocalMux I__1135 (
            .O(N__5158),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ));
    LocalMux I__1134 (
            .O(N__5155),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ));
    InMux I__1133 (
            .O(N__5150),
            .I(N__5139));
    InMux I__1132 (
            .O(N__5149),
            .I(N__5139));
    InMux I__1131 (
            .O(N__5148),
            .I(N__5139));
    InMux I__1130 (
            .O(N__5147),
            .I(N__5136));
    InMux I__1129 (
            .O(N__5146),
            .I(N__5133));
    LocalMux I__1128 (
            .O(N__5139),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__1127 (
            .O(N__5136),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__1126 (
            .O(N__5133),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    CascadeMux I__1125 (
            .O(N__5126),
            .I(N__5121));
    InMux I__1124 (
            .O(N__5125),
            .I(N__5117));
    InMux I__1123 (
            .O(N__5124),
            .I(N__5114));
    InMux I__1122 (
            .O(N__5121),
            .I(N__5109));
    InMux I__1121 (
            .O(N__5120),
            .I(N__5109));
    LocalMux I__1120 (
            .O(N__5117),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1119 (
            .O(N__5114),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1118 (
            .O(N__5109),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    CascadeMux I__1117 (
            .O(N__5102),
            .I(N__5096));
    InMux I__1116 (
            .O(N__5101),
            .I(N__5093));
    InMux I__1115 (
            .O(N__5100),
            .I(N__5090));
    InMux I__1114 (
            .O(N__5099),
            .I(N__5085));
    InMux I__1113 (
            .O(N__5096),
            .I(N__5085));
    LocalMux I__1112 (
            .O(N__5093),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__1111 (
            .O(N__5090),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__1110 (
            .O(N__5085),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    InMux I__1109 (
            .O(N__5078),
            .I(N__5073));
    InMux I__1108 (
            .O(N__5077),
            .I(N__5068));
    InMux I__1107 (
            .O(N__5076),
            .I(N__5068));
    LocalMux I__1106 (
            .O(N__5073),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    LocalMux I__1105 (
            .O(N__5068),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    CascadeMux I__1104 (
            .O(N__5063),
            .I(N__5057));
    InMux I__1103 (
            .O(N__5062),
            .I(N__5052));
    InMux I__1102 (
            .O(N__5061),
            .I(N__5052));
    InMux I__1101 (
            .O(N__5060),
            .I(N__5047));
    InMux I__1100 (
            .O(N__5057),
            .I(N__5047));
    LocalMux I__1099 (
            .O(N__5052),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__1098 (
            .O(N__5047),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    CascadeMux I__1097 (
            .O(N__5042),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_ ));
    InMux I__1096 (
            .O(N__5039),
            .I(N__5032));
    InMux I__1095 (
            .O(N__5038),
            .I(N__5032));
    InMux I__1094 (
            .O(N__5037),
            .I(N__5029));
    LocalMux I__1093 (
            .O(N__5032),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    LocalMux I__1092 (
            .O(N__5029),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    CascadeMux I__1091 (
            .O(N__5024),
            .I(N__5021));
    InMux I__1090 (
            .O(N__5021),
            .I(N__5018));
    LocalMux I__1089 (
            .O(N__5018),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ));
    CascadeMux I__1088 (
            .O(N__5015),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ));
    InMux I__1087 (
            .O(N__5012),
            .I(N__5009));
    LocalMux I__1086 (
            .O(N__5009),
            .I(N__5005));
    InMux I__1085 (
            .O(N__5008),
            .I(N__5001));
    Span4Mux_v I__1084 (
            .O(N__5005),
            .I(N__4998));
    InMux I__1083 (
            .O(N__5004),
            .I(N__4995));
    LocalMux I__1082 (
            .O(N__5001),
            .I(N__4992));
    Sp12to4 I__1081 (
            .O(N__4998),
            .I(N__4987));
    LocalMux I__1080 (
            .O(N__4995),
            .I(N__4987));
    Span12Mux_h I__1079 (
            .O(N__4992),
            .I(N__4984));
    Span12Mux_h I__1078 (
            .O(N__4987),
            .I(N__4981));
    Span12Mux_v I__1077 (
            .O(N__4984),
            .I(N__4978));
    Span12Mux_v I__1076 (
            .O(N__4981),
            .I(N__4975));
    Odrv12 I__1075 (
            .O(N__4978),
            .I(TSn_c));
    Odrv12 I__1074 (
            .O(N__4975),
            .I(TSn_c));
    IoInMux I__1073 (
            .O(N__4970),
            .I(N__4962));
    CascadeMux I__1072 (
            .O(N__4969),
            .I(N__4959));
    CascadeMux I__1071 (
            .O(N__4968),
            .I(N__4956));
    InMux I__1070 (
            .O(N__4967),
            .I(N__4953));
    CascadeMux I__1069 (
            .O(N__4966),
            .I(N__4950));
    CascadeMux I__1068 (
            .O(N__4965),
            .I(N__4947));
    LocalMux I__1067 (
            .O(N__4962),
            .I(N__4944));
    InMux I__1066 (
            .O(N__4959),
            .I(N__4939));
    InMux I__1065 (
            .O(N__4956),
            .I(N__4939));
    LocalMux I__1064 (
            .O(N__4953),
            .I(N__4936));
    InMux I__1063 (
            .O(N__4950),
            .I(N__4933));
    InMux I__1062 (
            .O(N__4947),
            .I(N__4930));
    IoSpan4Mux I__1061 (
            .O(N__4944),
            .I(N__4927));
    LocalMux I__1060 (
            .O(N__4939),
            .I(N__4924));
    Span4Mux_h I__1059 (
            .O(N__4936),
            .I(N__4917));
    LocalMux I__1058 (
            .O(N__4933),
            .I(N__4917));
    LocalMux I__1057 (
            .O(N__4930),
            .I(N__4917));
    Span4Mux_s0_v I__1056 (
            .O(N__4927),
            .I(N__4914));
    Span4Mux_v I__1055 (
            .O(N__4924),
            .I(N__4911));
    Span4Mux_v I__1054 (
            .O(N__4917),
            .I(N__4908));
    Sp12to4 I__1053 (
            .O(N__4914),
            .I(N__4905));
    Sp12to4 I__1052 (
            .O(N__4911),
            .I(N__4900));
    Sp12to4 I__1051 (
            .O(N__4908),
            .I(N__4900));
    Span12Mux_v I__1050 (
            .O(N__4905),
            .I(N__4897));
    Span12Mux_h I__1049 (
            .O(N__4900),
            .I(N__4894));
    Span12Mux_v I__1048 (
            .O(N__4897),
            .I(N__4891));
    Span12Mux_v I__1047 (
            .O(N__4894),
            .I(N__4888));
    Odrv12 I__1046 (
            .O(N__4891),
            .I(CLK40_IN_c));
    Odrv12 I__1045 (
            .O(N__4888),
            .I(CLK40_IN_c));
    InMux I__1044 (
            .O(N__4883),
            .I(N__4879));
    InMux I__1043 (
            .O(N__4882),
            .I(N__4876));
    LocalMux I__1042 (
            .O(N__4879),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    LocalMux I__1041 (
            .O(N__4876),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    InMux I__1040 (
            .O(N__4871),
            .I(N__4868));
    LocalMux I__1039 (
            .O(N__4868),
            .I(N__4864));
    InMux I__1038 (
            .O(N__4867),
            .I(N__4861));
    Span4Mux_v I__1037 (
            .O(N__4864),
            .I(N__4857));
    LocalMux I__1036 (
            .O(N__4861),
            .I(N__4854));
    InMux I__1035 (
            .O(N__4860),
            .I(N__4851));
    Sp12to4 I__1034 (
            .O(N__4857),
            .I(N__4846));
    Span12Mux_v I__1033 (
            .O(N__4854),
            .I(N__4846));
    LocalMux I__1032 (
            .O(N__4851),
            .I(N__4843));
    Span12Mux_v I__1031 (
            .O(N__4846),
            .I(N__4840));
    Span12Mux_h I__1030 (
            .O(N__4843),
            .I(N__4837));
    Span12Mux_h I__1029 (
            .O(N__4840),
            .I(N__4832));
    Span12Mux_v I__1028 (
            .O(N__4837),
            .I(N__4832));
    Odrv12 I__1027 (
            .O(N__4832),
            .I(OVL_c));
    InMux I__1026 (
            .O(N__4829),
            .I(N__4826));
    LocalMux I__1025 (
            .O(N__4826),
            .I(N__4822));
    CascadeMux I__1024 (
            .O(N__4825),
            .I(N__4819));
    Span4Mux_v I__1023 (
            .O(N__4822),
            .I(N__4815));
    InMux I__1022 (
            .O(N__4819),
            .I(N__4812));
    InMux I__1021 (
            .O(N__4818),
            .I(N__4809));
    Sp12to4 I__1020 (
            .O(N__4815),
            .I(N__4802));
    LocalMux I__1019 (
            .O(N__4812),
            .I(N__4802));
    LocalMux I__1018 (
            .O(N__4809),
            .I(N__4802));
    Odrv12 I__1017 (
            .O(N__4802),
            .I(\U409_ADDRESS_DECODE.un6_ROMENZ0 ));
    IoInMux I__1016 (
            .O(N__4799),
            .I(N__4796));
    LocalMux I__1015 (
            .O(N__4796),
            .I(N__4793));
    IoSpan4Mux I__1014 (
            .O(N__4793),
            .I(N__4790));
    Span4Mux_s2_v I__1013 (
            .O(N__4790),
            .I(N__4787));
    Sp12to4 I__1012 (
            .O(N__4787),
            .I(N__4784));
    Span12Mux_v I__1011 (
            .O(N__4784),
            .I(N__4781));
    Odrv12 I__1010 (
            .O(N__4781),
            .I(U409_ADDRESS_DECODE_un1_nRAMSPACE_i));
    InMux I__1009 (
            .O(N__4778),
            .I(N__4774));
    InMux I__1008 (
            .O(N__4777),
            .I(N__4771));
    LocalMux I__1007 (
            .O(N__4774),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ));
    LocalMux I__1006 (
            .O(N__4771),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ));
    CEMux I__1005 (
            .O(N__4766),
            .I(N__4763));
    LocalMux I__1004 (
            .O(N__4763),
            .I(N__4760));
    Odrv4 I__1003 (
            .O(N__4760),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0 ));
    InMux I__1002 (
            .O(N__4757),
            .I(N__4742));
    InMux I__1001 (
            .O(N__4756),
            .I(N__4742));
    InMux I__1000 (
            .O(N__4755),
            .I(N__4742));
    InMux I__999 (
            .O(N__4754),
            .I(N__4742));
    InMux I__998 (
            .O(N__4753),
            .I(N__4735));
    InMux I__997 (
            .O(N__4752),
            .I(N__4735));
    InMux I__996 (
            .O(N__4751),
            .I(N__4735));
    LocalMux I__995 (
            .O(N__4742),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__994 (
            .O(N__4735),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    CascadeMux I__993 (
            .O(N__4730),
            .I(\U409_CIA.N_20_cascade_ ));
    InMux I__992 (
            .O(N__4727),
            .I(N__4724));
    LocalMux I__991 (
            .O(N__4724),
            .I(\U409_CIA.CLKCIA6_0_a2_1 ));
    CascadeMux I__990 (
            .O(N__4721),
            .I(N__4711));
    InMux I__989 (
            .O(N__4720),
            .I(N__4708));
    InMux I__988 (
            .O(N__4719),
            .I(N__4699));
    InMux I__987 (
            .O(N__4718),
            .I(N__4699));
    InMux I__986 (
            .O(N__4717),
            .I(N__4699));
    InMux I__985 (
            .O(N__4716),
            .I(N__4699));
    InMux I__984 (
            .O(N__4715),
            .I(N__4692));
    InMux I__983 (
            .O(N__4714),
            .I(N__4692));
    InMux I__982 (
            .O(N__4711),
            .I(N__4692));
    LocalMux I__981 (
            .O(N__4708),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__980 (
            .O(N__4699),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__979 (
            .O(N__4692),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    CascadeMux I__978 (
            .O(N__4685),
            .I(\U409_CIA.CLKCIAZ0_cascade_ ));
    InMux I__977 (
            .O(N__4682),
            .I(N__4668));
    InMux I__976 (
            .O(N__4681),
            .I(N__4668));
    InMux I__975 (
            .O(N__4680),
            .I(N__4668));
    InMux I__974 (
            .O(N__4679),
            .I(N__4668));
    InMux I__973 (
            .O(N__4678),
            .I(N__4663));
    InMux I__972 (
            .O(N__4677),
            .I(N__4663));
    LocalMux I__971 (
            .O(N__4668),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__970 (
            .O(N__4663),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    IoInMux I__969 (
            .O(N__4658),
            .I(N__4655));
    LocalMux I__968 (
            .O(N__4655),
            .I(N__4652));
    Span4Mux_s0_v I__967 (
            .O(N__4652),
            .I(N__4649));
    Sp12to4 I__966 (
            .O(N__4649),
            .I(N__4646));
    Span12Mux_h I__965 (
            .O(N__4646),
            .I(N__4643));
    Span12Mux_v I__964 (
            .O(N__4643),
            .I(N__4638));
    InMux I__963 (
            .O(N__4642),
            .I(N__4635));
    InMux I__962 (
            .O(N__4641),
            .I(N__4632));
    Odrv12 I__961 (
            .O(N__4638),
            .I(CLKCIA_c));
    LocalMux I__960 (
            .O(N__4635),
            .I(CLKCIA_c));
    LocalMux I__959 (
            .O(N__4632),
            .I(CLKCIA_c));
    ClkMux I__958 (
            .O(N__4625),
            .I(N__4613));
    ClkMux I__957 (
            .O(N__4624),
            .I(N__4613));
    ClkMux I__956 (
            .O(N__4623),
            .I(N__4613));
    ClkMux I__955 (
            .O(N__4622),
            .I(N__4613));
    GlobalMux I__954 (
            .O(N__4613),
            .I(N__4610));
    gio2CtrlBuf I__953 (
            .O(N__4610),
            .I(CLK28_IN_c_g));
    CascadeMux I__952 (
            .O(N__4607),
            .I(N__4603));
    CascadeMux I__951 (
            .O(N__4606),
            .I(N__4599));
    InMux I__950 (
            .O(N__4603),
            .I(N__4593));
    InMux I__949 (
            .O(N__4602),
            .I(N__4593));
    InMux I__948 (
            .O(N__4599),
            .I(N__4588));
    InMux I__947 (
            .O(N__4598),
            .I(N__4588));
    LocalMux I__946 (
            .O(N__4593),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__945 (
            .O(N__4588),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    InMux I__944 (
            .O(N__4583),
            .I(N__4577));
    InMux I__943 (
            .O(N__4582),
            .I(N__4572));
    InMux I__942 (
            .O(N__4581),
            .I(N__4572));
    InMux I__941 (
            .O(N__4580),
            .I(N__4569));
    LocalMux I__940 (
            .O(N__4577),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__939 (
            .O(N__4572),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__938 (
            .O(N__4569),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    InMux I__937 (
            .O(N__4562),
            .I(N__4554));
    InMux I__936 (
            .O(N__4561),
            .I(N__4554));
    InMux I__935 (
            .O(N__4560),
            .I(N__4549));
    InMux I__934 (
            .O(N__4559),
            .I(N__4549));
    LocalMux I__933 (
            .O(N__4554),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__932 (
            .O(N__4549),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    InMux I__931 (
            .O(N__4544),
            .I(N__4538));
    InMux I__930 (
            .O(N__4543),
            .I(N__4538));
    LocalMux I__929 (
            .O(N__4538),
            .I(\U409_CIA.CLKCIA8_0_a2_0 ));
    CascadeMux I__928 (
            .O(N__4535),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_ ));
    InMux I__927 (
            .O(N__4532),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ));
    InMux I__926 (
            .O(N__4529),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ));
    InMux I__925 (
            .O(N__4526),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ));
    InMux I__924 (
            .O(N__4523),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ));
    CascadeMux I__923 (
            .O(N__4520),
            .I(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_ ));
    InMux I__922 (
            .O(N__4517),
            .I(N__4514));
    LocalMux I__921 (
            .O(N__4514),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ));
    CascadeMux I__920 (
            .O(N__4511),
            .I(N__4508));
    InMux I__919 (
            .O(N__4508),
            .I(N__4502));
    InMux I__918 (
            .O(N__4507),
            .I(N__4502));
    LocalMux I__917 (
            .O(N__4502),
            .I(\U409_CIA.CIA_CLK_COUNT11_0_a2_2 ));
    CascadeMux I__916 (
            .O(N__4499),
            .I(\U409_CIA.N_9_cascade_ ));
    CascadeMux I__915 (
            .O(N__4496),
            .I(N__4493));
    InMux I__914 (
            .O(N__4493),
            .I(N__4488));
    InMux I__913 (
            .O(N__4492),
            .I(N__4483));
    InMux I__912 (
            .O(N__4491),
            .I(N__4483));
    LocalMux I__911 (
            .O(N__4488),
            .I(N__4480));
    LocalMux I__910 (
            .O(N__4483),
            .I(N__4476));
    Span4Mux_v I__909 (
            .O(N__4480),
            .I(N__4473));
    InMux I__908 (
            .O(N__4479),
            .I(N__4470));
    Span4Mux_h I__907 (
            .O(N__4476),
            .I(N__4467));
    Odrv4 I__906 (
            .O(N__4473),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__905 (
            .O(N__4470),
            .I(\U409_CIA.VMAZ0 ));
    Odrv4 I__904 (
            .O(N__4467),
            .I(\U409_CIA.VMAZ0 ));
    InMux I__903 (
            .O(N__4460),
            .I(N__4452));
    InMux I__902 (
            .O(N__4459),
            .I(N__4452));
    InMux I__901 (
            .O(N__4458),
            .I(N__4447));
    InMux I__900 (
            .O(N__4457),
            .I(N__4447));
    LocalMux I__899 (
            .O(N__4452),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__898 (
            .O(N__4447),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    InMux I__897 (
            .O(N__4442),
            .I(N__4439));
    LocalMux I__896 (
            .O(N__4439),
            .I(N__4434));
    InMux I__895 (
            .O(N__4438),
            .I(N__4431));
    InMux I__894 (
            .O(N__4437),
            .I(N__4428));
    Odrv4 I__893 (
            .O(N__4434),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    LocalMux I__892 (
            .O(N__4431),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    LocalMux I__891 (
            .O(N__4428),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    InMux I__890 (
            .O(N__4421),
            .I(N__4417));
    InMux I__889 (
            .O(N__4420),
            .I(N__4414));
    LocalMux I__888 (
            .O(N__4417),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    LocalMux I__887 (
            .O(N__4414),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    InMux I__886 (
            .O(N__4409),
            .I(N__4406));
    LocalMux I__885 (
            .O(N__4406),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER5_0 ));
    CascadeMux I__884 (
            .O(N__4403),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_ ));
    IoInMux I__883 (
            .O(N__4400),
            .I(N__4397));
    LocalMux I__882 (
            .O(N__4397),
            .I(N__4394));
    IoSpan4Mux I__881 (
            .O(N__4394),
            .I(N__4391));
    Span4Mux_s1_v I__880 (
            .O(N__4391),
            .I(N__4388));
    Sp12to4 I__879 (
            .O(N__4388),
            .I(N__4385));
    Span12Mux_v I__878 (
            .O(N__4385),
            .I(N__4381));
    InMux I__877 (
            .O(N__4384),
            .I(N__4378));
    Odrv12 I__876 (
            .O(N__4381),
            .I(TACK_OUTn));
    LocalMux I__875 (
            .O(N__4378),
            .I(TACK_OUTn));
    CascadeMux I__874 (
            .O(N__4373),
            .I(N__4368));
    InMux I__873 (
            .O(N__4372),
            .I(N__4361));
    InMux I__872 (
            .O(N__4371),
            .I(N__4361));
    InMux I__871 (
            .O(N__4368),
            .I(N__4361));
    LocalMux I__870 (
            .O(N__4361),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    InMux I__869 (
            .O(N__4358),
            .I(N__4349));
    InMux I__868 (
            .O(N__4357),
            .I(N__4349));
    InMux I__867 (
            .O(N__4356),
            .I(N__4349));
    LocalMux I__866 (
            .O(N__4349),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    IoInMux I__865 (
            .O(N__4346),
            .I(N__4343));
    LocalMux I__864 (
            .O(N__4343),
            .I(N__4340));
    Span4Mux_s2_v I__863 (
            .O(N__4340),
            .I(N__4337));
    Span4Mux_v I__862 (
            .O(N__4337),
            .I(N__4334));
    Span4Mux_v I__861 (
            .O(N__4334),
            .I(N__4331));
    Sp12to4 I__860 (
            .O(N__4331),
            .I(N__4327));
    InMux I__859 (
            .O(N__4330),
            .I(N__4324));
    Odrv12 I__858 (
            .O(N__4327),
            .I(TICK50_c));
    LocalMux I__857 (
            .O(N__4324),
            .I(TICK50_c));
    CascadeMux I__856 (
            .O(N__4319),
            .I(N__4312));
    CascadeMux I__855 (
            .O(N__4318),
            .I(N__4309));
    InMux I__854 (
            .O(N__4317),
            .I(N__4303));
    InMux I__853 (
            .O(N__4316),
            .I(N__4300));
    InMux I__852 (
            .O(N__4315),
            .I(N__4291));
    InMux I__851 (
            .O(N__4312),
            .I(N__4291));
    InMux I__850 (
            .O(N__4309),
            .I(N__4291));
    InMux I__849 (
            .O(N__4308),
            .I(N__4291));
    InMux I__848 (
            .O(N__4307),
            .I(N__4286));
    InMux I__847 (
            .O(N__4306),
            .I(N__4286));
    LocalMux I__846 (
            .O(N__4303),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__845 (
            .O(N__4300),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__844 (
            .O(N__4291),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__843 (
            .O(N__4286),
            .I(\U409_TICK.TICK503_10 ));
    InMux I__842 (
            .O(N__4277),
            .I(N__4267));
    InMux I__841 (
            .O(N__4276),
            .I(N__4264));
    InMux I__840 (
            .O(N__4275),
            .I(N__4255));
    InMux I__839 (
            .O(N__4274),
            .I(N__4255));
    InMux I__838 (
            .O(N__4273),
            .I(N__4255));
    InMux I__837 (
            .O(N__4272),
            .I(N__4255));
    InMux I__836 (
            .O(N__4271),
            .I(N__4250));
    InMux I__835 (
            .O(N__4270),
            .I(N__4250));
    LocalMux I__834 (
            .O(N__4267),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__833 (
            .O(N__4264),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__832 (
            .O(N__4255),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__831 (
            .O(N__4250),
            .I(\U409_TICK.TICK503_14 ));
    CascadeMux I__830 (
            .O(N__4241),
            .I(N__4237));
    CascadeMux I__829 (
            .O(N__4240),
            .I(N__4234));
    InMux I__828 (
            .O(N__4237),
            .I(N__4225));
    InMux I__827 (
            .O(N__4234),
            .I(N__4222));
    InMux I__826 (
            .O(N__4233),
            .I(N__4215));
    InMux I__825 (
            .O(N__4232),
            .I(N__4215));
    InMux I__824 (
            .O(N__4231),
            .I(N__4215));
    InMux I__823 (
            .O(N__4230),
            .I(N__4208));
    InMux I__822 (
            .O(N__4229),
            .I(N__4208));
    InMux I__821 (
            .O(N__4228),
            .I(N__4208));
    LocalMux I__820 (
            .O(N__4225),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__819 (
            .O(N__4222),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__818 (
            .O(N__4215),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__817 (
            .O(N__4208),
            .I(\U409_TICK.TICK503_9 ));
    InMux I__816 (
            .O(N__4199),
            .I(N__4196));
    LocalMux I__815 (
            .O(N__4196),
            .I(N__4193));
    Odrv4 I__814 (
            .O(N__4193),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ));
    InMux I__813 (
            .O(N__4190),
            .I(N__4186));
    InMux I__812 (
            .O(N__4189),
            .I(N__4183));
    LocalMux I__811 (
            .O(N__4186),
            .I(N__4180));
    LocalMux I__810 (
            .O(N__4183),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    Odrv4 I__809 (
            .O(N__4180),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    ClkMux I__808 (
            .O(N__4175),
            .I(N__4142));
    ClkMux I__807 (
            .O(N__4174),
            .I(N__4142));
    ClkMux I__806 (
            .O(N__4173),
            .I(N__4142));
    ClkMux I__805 (
            .O(N__4172),
            .I(N__4142));
    ClkMux I__804 (
            .O(N__4171),
            .I(N__4142));
    ClkMux I__803 (
            .O(N__4170),
            .I(N__4142));
    ClkMux I__802 (
            .O(N__4169),
            .I(N__4142));
    ClkMux I__801 (
            .O(N__4168),
            .I(N__4142));
    ClkMux I__800 (
            .O(N__4167),
            .I(N__4142));
    ClkMux I__799 (
            .O(N__4166),
            .I(N__4142));
    ClkMux I__798 (
            .O(N__4165),
            .I(N__4142));
    GlobalMux I__797 (
            .O(N__4142),
            .I(N__4139));
    gio2CtrlBuf I__796 (
            .O(N__4139),
            .I(CLK6_c_g));
    InMux I__795 (
            .O(N__4136),
            .I(N__4130));
    InMux I__794 (
            .O(N__4135),
            .I(N__4130));
    LocalMux I__793 (
            .O(N__4130),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    InMux I__792 (
            .O(N__4127),
            .I(N__4118));
    InMux I__791 (
            .O(N__4126),
            .I(N__4118));
    InMux I__790 (
            .O(N__4125),
            .I(N__4118));
    LocalMux I__789 (
            .O(N__4118),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    CascadeMux I__788 (
            .O(N__4115),
            .I(\U409_TRANSFER_ACK.N_4_cascade_ ));
    InMux I__787 (
            .O(N__4112),
            .I(N__4109));
    LocalMux I__786 (
            .O(N__4109),
            .I(\U409_TRANSFER_ACK.N_97 ));
    CascadeMux I__785 (
            .O(N__4106),
            .I(\U409_TRANSFER_ACK.CIA_TACK_EN_0_cascade_ ));
    InMux I__784 (
            .O(N__4103),
            .I(N__4100));
    LocalMux I__783 (
            .O(N__4100),
            .I(\U409_TRANSFER_ACK.i6_mux_0 ));
    InMux I__782 (
            .O(N__4097),
            .I(N__4093));
    InMux I__781 (
            .O(N__4096),
            .I(N__4090));
    LocalMux I__780 (
            .O(N__4093),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    LocalMux I__779 (
            .O(N__4090),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    InMux I__778 (
            .O(N__4085),
            .I(N__4082));
    LocalMux I__777 (
            .O(N__4082),
            .I(\U409_TRANSFER_ACK.N_4 ));
    InMux I__776 (
            .O(N__4079),
            .I(N__4076));
    LocalMux I__775 (
            .O(N__4076),
            .I(\U409_TRANSFER_ACK.m9_bm ));
    CascadeMux I__774 (
            .O(N__4073),
            .I(\U409_TRANSFER_ACK.m9_am_cascade_ ));
    InMux I__773 (
            .O(N__4070),
            .I(N__4063));
    InMux I__772 (
            .O(N__4069),
            .I(N__4054));
    InMux I__771 (
            .O(N__4068),
            .I(N__4054));
    InMux I__770 (
            .O(N__4067),
            .I(N__4054));
    InMux I__769 (
            .O(N__4066),
            .I(N__4054));
    LocalMux I__768 (
            .O(N__4063),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__767 (
            .O(N__4054),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    CascadeMux I__766 (
            .O(N__4049),
            .I(N__4044));
    CascadeMux I__765 (
            .O(N__4048),
            .I(N__4041));
    CascadeMux I__764 (
            .O(N__4047),
            .I(N__4037));
    InMux I__763 (
            .O(N__4044),
            .I(N__4032));
    InMux I__762 (
            .O(N__4041),
            .I(N__4032));
    InMux I__761 (
            .O(N__4040),
            .I(N__4029));
    InMux I__760 (
            .O(N__4037),
            .I(N__4026));
    LocalMux I__759 (
            .O(N__4032),
            .I(N__4021));
    LocalMux I__758 (
            .O(N__4029),
            .I(N__4021));
    LocalMux I__757 (
            .O(N__4026),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    Odrv4 I__756 (
            .O(N__4021),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    CascadeMux I__755 (
            .O(N__4016),
            .I(N__4013));
    InMux I__754 (
            .O(N__4013),
            .I(N__4009));
    InMux I__753 (
            .O(N__4012),
            .I(N__4006));
    LocalMux I__752 (
            .O(N__4009),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    LocalMux I__751 (
            .O(N__4006),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    InMux I__750 (
            .O(N__4001),
            .I(N__3997));
    InMux I__749 (
            .O(N__4000),
            .I(N__3994));
    LocalMux I__748 (
            .O(N__3997),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    LocalMux I__747 (
            .O(N__3994),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    InMux I__746 (
            .O(N__3989),
            .I(N__3986));
    LocalMux I__745 (
            .O(N__3986),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ));
    CascadeMux I__744 (
            .O(N__3983),
            .I(\U409_TICK.TICK503_9_cascade_ ));
    InMux I__743 (
            .O(N__3980),
            .I(N__3976));
    InMux I__742 (
            .O(N__3979),
            .I(N__3973));
    LocalMux I__741 (
            .O(N__3976),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    LocalMux I__740 (
            .O(N__3973),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    InMux I__739 (
            .O(N__3968),
            .I(N__3965));
    LocalMux I__738 (
            .O(N__3965),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ));
    InMux I__737 (
            .O(N__3962),
            .I(N__3958));
    InMux I__736 (
            .O(N__3961),
            .I(N__3955));
    LocalMux I__735 (
            .O(N__3958),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    LocalMux I__734 (
            .O(N__3955),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    CascadeMux I__733 (
            .O(N__3950),
            .I(N__3947));
    InMux I__732 (
            .O(N__3947),
            .I(N__3944));
    LocalMux I__731 (
            .O(N__3944),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ));
    InMux I__730 (
            .O(N__3941),
            .I(N__3937));
    InMux I__729 (
            .O(N__3940),
            .I(N__3934));
    LocalMux I__728 (
            .O(N__3937),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    LocalMux I__727 (
            .O(N__3934),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    CascadeMux I__726 (
            .O(N__3929),
            .I(\U409_TRANSFER_ACK.N_97_cascade_ ));
    InMux I__725 (
            .O(N__3926),
            .I(N__3922));
    InMux I__724 (
            .O(N__3925),
            .I(N__3919));
    LocalMux I__723 (
            .O(N__3922),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    LocalMux I__722 (
            .O(N__3919),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    InMux I__721 (
            .O(N__3914),
            .I(N__3910));
    InMux I__720 (
            .O(N__3913),
            .I(N__3907));
    LocalMux I__719 (
            .O(N__3910),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    LocalMux I__718 (
            .O(N__3907),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    CascadeMux I__717 (
            .O(N__3902),
            .I(\U409_TICK.TICK503_8_cascade_ ));
    InMux I__716 (
            .O(N__3899),
            .I(N__3895));
    InMux I__715 (
            .O(N__3898),
            .I(N__3892));
    LocalMux I__714 (
            .O(N__3895),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    LocalMux I__713 (
            .O(N__3892),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    CascadeMux I__712 (
            .O(N__3887),
            .I(\U409_TICK.TICK503_14_cascade_ ));
    CascadeMux I__711 (
            .O(N__3884),
            .I(N__3878));
    InMux I__710 (
            .O(N__3883),
            .I(N__3871));
    InMux I__709 (
            .O(N__3882),
            .I(N__3871));
    InMux I__708 (
            .O(N__3881),
            .I(N__3871));
    InMux I__707 (
            .O(N__3878),
            .I(N__3868));
    LocalMux I__706 (
            .O(N__3871),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__705 (
            .O(N__3868),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    InMux I__704 (
            .O(N__3863),
            .I(N__3859));
    InMux I__703 (
            .O(N__3862),
            .I(N__3856));
    LocalMux I__702 (
            .O(N__3859),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    LocalMux I__701 (
            .O(N__3856),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    CascadeMux I__700 (
            .O(N__3851),
            .I(N__3848));
    InMux I__699 (
            .O(N__3848),
            .I(N__3844));
    InMux I__698 (
            .O(N__3847),
            .I(N__3841));
    LocalMux I__697 (
            .O(N__3844),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    LocalMux I__696 (
            .O(N__3841),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    CascadeMux I__695 (
            .O(N__3836),
            .I(\U409_TICK.TICK503_10_cascade_ ));
    InMux I__694 (
            .O(N__3833),
            .I(N__3830));
    LocalMux I__693 (
            .O(N__3830),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ));
    InMux I__692 (
            .O(N__3827),
            .I(N__3823));
    InMux I__691 (
            .O(N__3826),
            .I(N__3820));
    LocalMux I__690 (
            .O(N__3823),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    LocalMux I__689 (
            .O(N__3820),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    InMux I__688 (
            .O(N__3815),
            .I(N__3811));
    InMux I__687 (
            .O(N__3814),
            .I(N__3808));
    LocalMux I__686 (
            .O(N__3811),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    LocalMux I__685 (
            .O(N__3808),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    InMux I__684 (
            .O(N__3803),
            .I(N__3799));
    InMux I__683 (
            .O(N__3802),
            .I(N__3796));
    LocalMux I__682 (
            .O(N__3799),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    LocalMux I__681 (
            .O(N__3796),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    CascadeMux I__680 (
            .O(N__3791),
            .I(N__3787));
    InMux I__679 (
            .O(N__3790),
            .I(N__3782));
    InMux I__678 (
            .O(N__3787),
            .I(N__3782));
    LocalMux I__677 (
            .O(N__3782),
            .I(N__3778));
    InMux I__676 (
            .O(N__3781),
            .I(N__3775));
    Odrv4 I__675 (
            .O(N__3778),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    LocalMux I__674 (
            .O(N__3775),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    InMux I__673 (
            .O(N__3770),
            .I(N__3766));
    InMux I__672 (
            .O(N__3769),
            .I(N__3763));
    LocalMux I__671 (
            .O(N__3766),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    LocalMux I__670 (
            .O(N__3763),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    InMux I__669 (
            .O(N__3758),
            .I(N__3755));
    LocalMux I__668 (
            .O(N__3755),
            .I(\U409_TICK.TICK503_11 ));
    CascadeMux I__667 (
            .O(N__3752),
            .I(N__3749));
    InMux I__666 (
            .O(N__3749),
            .I(N__3746));
    LocalMux I__665 (
            .O(N__3746),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ));
    InMux I__664 (
            .O(N__3743),
            .I(N__3740));
    LocalMux I__663 (
            .O(N__3740),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ));
    InMux I__662 (
            .O(N__3737),
            .I(N__3731));
    InMux I__661 (
            .O(N__3736),
            .I(N__3731));
    LocalMux I__660 (
            .O(N__3731),
            .I(N__3728));
    Odrv12 I__659 (
            .O(N__3728),
            .I(CIA_ENABLEm));
    InMux I__658 (
            .O(N__3725),
            .I(N__3722));
    LocalMux I__657 (
            .O(N__3722),
            .I(N__3717));
    InMux I__656 (
            .O(N__3721),
            .I(N__3712));
    InMux I__655 (
            .O(N__3720),
            .I(N__3712));
    Odrv4 I__654 (
            .O(N__3717),
            .I(\U409_CIA.CIA_HOLDZ0 ));
    LocalMux I__653 (
            .O(N__3712),
            .I(\U409_CIA.CIA_HOLDZ0 ));
    InMux I__652 (
            .O(N__3707),
            .I(N__3701));
    InMux I__651 (
            .O(N__3706),
            .I(N__3701));
    LocalMux I__650 (
            .O(N__3701),
            .I(N__3698));
    Span4Mux_v I__649 (
            .O(N__3698),
            .I(N__3694));
    InMux I__648 (
            .O(N__3697),
            .I(N__3691));
    Sp12to4 I__647 (
            .O(N__3694),
            .I(N__3686));
    LocalMux I__646 (
            .O(N__3691),
            .I(N__3686));
    Odrv12 I__645 (
            .O(N__3686),
            .I(\U409_CIA.g0Z0Z_14 ));
    CascadeMux I__644 (
            .O(N__3683),
            .I(N__3679));
    CascadeMux I__643 (
            .O(N__3682),
            .I(N__3676));
    InMux I__642 (
            .O(N__3679),
            .I(N__3671));
    InMux I__641 (
            .O(N__3676),
            .I(N__3671));
    LocalMux I__640 (
            .O(N__3671),
            .I(N__3667));
    InMux I__639 (
            .O(N__3670),
            .I(N__3664));
    Span4Mux_h I__638 (
            .O(N__3667),
            .I(N__3659));
    LocalMux I__637 (
            .O(N__3664),
            .I(N__3659));
    Span4Mux_v I__636 (
            .O(N__3659),
            .I(N__3656));
    Span4Mux_v I__635 (
            .O(N__3656),
            .I(N__3653));
    Span4Mux_h I__634 (
            .O(N__3653),
            .I(N__3650));
    Odrv4 I__633 (
            .O(N__3650),
            .I(\U409_CIA.g0Z0Z_13 ));
    SRMux I__632 (
            .O(N__3647),
            .I(N__3644));
    LocalMux I__631 (
            .O(N__3644),
            .I(N__3641));
    Odrv4 I__630 (
            .O(N__3641),
            .I(\U409_TRANSFER_ACK.RESETn_c_i ));
    CascadeMux I__629 (
            .O(N__3638),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_3_0_cascade_ ));
    CascadeMux I__628 (
            .O(N__3635),
            .I(\U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa_cascade_ ));
    InMux I__627 (
            .O(N__3632),
            .I(N__3624));
    InMux I__626 (
            .O(N__3631),
            .I(N__3624));
    InMux I__625 (
            .O(N__3630),
            .I(N__3619));
    InMux I__624 (
            .O(N__3629),
            .I(N__3619));
    LocalMux I__623 (
            .O(N__3624),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__622 (
            .O(N__3619),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    InMux I__621 (
            .O(N__3614),
            .I(N__3599));
    InMux I__620 (
            .O(N__3613),
            .I(N__3599));
    InMux I__619 (
            .O(N__3612),
            .I(N__3599));
    InMux I__618 (
            .O(N__3611),
            .I(N__3599));
    InMux I__617 (
            .O(N__3610),
            .I(N__3599));
    LocalMux I__616 (
            .O(N__3599),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    InMux I__615 (
            .O(N__3596),
            .I(N__3590));
    InMux I__614 (
            .O(N__3595),
            .I(N__3590));
    LocalMux I__613 (
            .O(N__3590),
            .I(\U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0 ));
    IoInMux I__612 (
            .O(N__3587),
            .I(N__3584));
    LocalMux I__611 (
            .O(N__3584),
            .I(N__3581));
    Span4Mux_s0_v I__610 (
            .O(N__3581),
            .I(N__3578));
    Sp12to4 I__609 (
            .O(N__3578),
            .I(N__3575));
    Span12Mux_h I__608 (
            .O(N__3575),
            .I(N__3572));
    Span12Mux_v I__607 (
            .O(N__3572),
            .I(N__3568));
    InMux I__606 (
            .O(N__3571),
            .I(N__3565));
    Odrv12 I__605 (
            .O(N__3568),
            .I(TICK60_c));
    LocalMux I__604 (
            .O(N__3565),
            .I(TICK60_c));
    CascadeMux I__603 (
            .O(N__3560),
            .I(N__3557));
    InMux I__602 (
            .O(N__3557),
            .I(N__3554));
    LocalMux I__601 (
            .O(N__3554),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ));
    InMux I__600 (
            .O(N__3551),
            .I(N__3547));
    InMux I__599 (
            .O(N__3550),
            .I(N__3544));
    LocalMux I__598 (
            .O(N__3547),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    LocalMux I__597 (
            .O(N__3544),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    InMux I__596 (
            .O(N__3539),
            .I(N__3535));
    InMux I__595 (
            .O(N__3538),
            .I(N__3532));
    LocalMux I__594 (
            .O(N__3535),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    LocalMux I__593 (
            .O(N__3532),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    CascadeMux I__592 (
            .O(N__3527),
            .I(\U409_TICK.TICK603_9_cascade_ ));
    InMux I__591 (
            .O(N__3524),
            .I(N__3521));
    LocalMux I__590 (
            .O(N__3521),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ));
    CascadeMux I__589 (
            .O(N__3518),
            .I(N__3515));
    InMux I__588 (
            .O(N__3515),
            .I(N__3512));
    LocalMux I__587 (
            .O(N__3512),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ));
    CascadeMux I__586 (
            .O(N__3509),
            .I(N__3506));
    InMux I__585 (
            .O(N__3506),
            .I(N__3502));
    InMux I__584 (
            .O(N__3505),
            .I(N__3499));
    LocalMux I__583 (
            .O(N__3502),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    LocalMux I__582 (
            .O(N__3499),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    InMux I__581 (
            .O(N__3494),
            .I(N__3490));
    InMux I__580 (
            .O(N__3493),
            .I(N__3487));
    LocalMux I__579 (
            .O(N__3490),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    LocalMux I__578 (
            .O(N__3487),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    InMux I__577 (
            .O(N__3482),
            .I(N__3478));
    InMux I__576 (
            .O(N__3481),
            .I(N__3475));
    LocalMux I__575 (
            .O(N__3478),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    LocalMux I__574 (
            .O(N__3475),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    CascadeMux I__573 (
            .O(N__3470),
            .I(N__3467));
    InMux I__572 (
            .O(N__3467),
            .I(N__3463));
    InMux I__571 (
            .O(N__3466),
            .I(N__3460));
    LocalMux I__570 (
            .O(N__3463),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    LocalMux I__569 (
            .O(N__3460),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    InMux I__568 (
            .O(N__3455),
            .I(N__3451));
    InMux I__567 (
            .O(N__3454),
            .I(N__3448));
    LocalMux I__566 (
            .O(N__3451),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    LocalMux I__565 (
            .O(N__3448),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    InMux I__564 (
            .O(N__3443),
            .I(N__3434));
    InMux I__563 (
            .O(N__3442),
            .I(N__3434));
    InMux I__562 (
            .O(N__3441),
            .I(N__3434));
    LocalMux I__561 (
            .O(N__3434),
            .I(N__3427));
    InMux I__560 (
            .O(N__3433),
            .I(N__3420));
    InMux I__559 (
            .O(N__3432),
            .I(N__3420));
    InMux I__558 (
            .O(N__3431),
            .I(N__3420));
    InMux I__557 (
            .O(N__3430),
            .I(N__3417));
    Odrv4 I__556 (
            .O(N__3427),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__555 (
            .O(N__3420),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__554 (
            .O(N__3417),
            .I(\U409_TICK.TICK603_10 ));
    InMux I__553 (
            .O(N__3410),
            .I(N__3395));
    InMux I__552 (
            .O(N__3409),
            .I(N__3395));
    InMux I__551 (
            .O(N__3408),
            .I(N__3395));
    InMux I__550 (
            .O(N__3407),
            .I(N__3395));
    InMux I__549 (
            .O(N__3406),
            .I(N__3392));
    InMux I__548 (
            .O(N__3405),
            .I(N__3387));
    InMux I__547 (
            .O(N__3404),
            .I(N__3387));
    LocalMux I__546 (
            .O(N__3395),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__545 (
            .O(N__3392),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__544 (
            .O(N__3387),
            .I(\U409_TICK.TICK603_14 ));
    CascadeMux I__543 (
            .O(N__3380),
            .I(N__3375));
    CascadeMux I__542 (
            .O(N__3379),
            .I(N__3368));
    CascadeMux I__541 (
            .O(N__3378),
            .I(N__3365));
    InMux I__540 (
            .O(N__3375),
            .I(N__3362));
    InMux I__539 (
            .O(N__3374),
            .I(N__3355));
    InMux I__538 (
            .O(N__3373),
            .I(N__3355));
    InMux I__537 (
            .O(N__3372),
            .I(N__3355));
    InMux I__536 (
            .O(N__3371),
            .I(N__3348));
    InMux I__535 (
            .O(N__3368),
            .I(N__3348));
    InMux I__534 (
            .O(N__3365),
            .I(N__3348));
    LocalMux I__533 (
            .O(N__3362),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__532 (
            .O(N__3355),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__531 (
            .O(N__3348),
            .I(\U409_TICK.TICK603_9 ));
    CascadeMux I__530 (
            .O(N__3341),
            .I(\U409_TICK.TICK603_10_cascade_ ));
    InMux I__529 (
            .O(N__3338),
            .I(N__3335));
    LocalMux I__528 (
            .O(N__3335),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ));
    InMux I__527 (
            .O(N__3332),
            .I(N__3328));
    InMux I__526 (
            .O(N__3331),
            .I(N__3325));
    LocalMux I__525 (
            .O(N__3328),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    LocalMux I__524 (
            .O(N__3325),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    InMux I__523 (
            .O(N__3320),
            .I(\U409_TICK.un2_COUNTER50_1_cry_7 ));
    InMux I__522 (
            .O(N__3317),
            .I(bfn_9_6_0_));
    InMux I__521 (
            .O(N__3314),
            .I(\U409_TICK.un2_COUNTER50_1_cry_9 ));
    InMux I__520 (
            .O(N__3311),
            .I(\U409_TICK.un2_COUNTER50_1_cry_10 ));
    InMux I__519 (
            .O(N__3308),
            .I(\U409_TICK.un2_COUNTER50_1_cry_11 ));
    InMux I__518 (
            .O(N__3305),
            .I(\U409_TICK.un2_COUNTER50_1_cry_12 ));
    InMux I__517 (
            .O(N__3302),
            .I(\U409_TICK.un2_COUNTER50_1_cry_13 ));
    InMux I__516 (
            .O(N__3299),
            .I(\U409_TICK.un2_COUNTER50_1_cry_14 ));
    InMux I__515 (
            .O(N__3296),
            .I(\U409_TICK.un2_COUNTER50_1_cry_15 ));
    InMux I__514 (
            .O(N__3293),
            .I(N__3290));
    LocalMux I__513 (
            .O(N__3290),
            .I(N__3287));
    Span4Mux_v I__512 (
            .O(N__3287),
            .I(N__3284));
    Sp12to4 I__511 (
            .O(N__3284),
            .I(N__3281));
    Span12Mux_h I__510 (
            .O(N__3281),
            .I(N__3278));
    Odrv12 I__509 (
            .O(N__3278),
            .I(A_c_13));
    IoInMux I__508 (
            .O(N__3275),
            .I(N__3272));
    LocalMux I__507 (
            .O(N__3272),
            .I(N__3269));
    Span4Mux_s1_h I__506 (
            .O(N__3269),
            .I(N__3266));
    Sp12to4 I__505 (
            .O(N__3266),
            .I(N__3263));
    Span12Mux_s9_v I__504 (
            .O(N__3263),
            .I(N__3260));
    Span12Mux_h I__503 (
            .O(N__3260),
            .I(N__3257));
    Odrv12 I__502 (
            .O(N__3257),
            .I(U409_ADDRESS_DECODE_un1_nCIACS1_i));
    InMux I__501 (
            .O(N__3254),
            .I(N__3251));
    LocalMux I__500 (
            .O(N__3251),
            .I(N__3248));
    Span4Mux_v I__499 (
            .O(N__3248),
            .I(N__3245));
    Sp12to4 I__498 (
            .O(N__3245),
            .I(N__3242));
    Odrv12 I__497 (
            .O(N__3242),
            .I(A_c_12));
    IoInMux I__496 (
            .O(N__3239),
            .I(N__3236));
    LocalMux I__495 (
            .O(N__3236),
            .I(N__3233));
    Span4Mux_s2_h I__494 (
            .O(N__3233),
            .I(N__3230));
    Sp12to4 I__493 (
            .O(N__3230),
            .I(N__3227));
    Span12Mux_s9_v I__492 (
            .O(N__3227),
            .I(N__3224));
    Span12Mux_h I__491 (
            .O(N__3224),
            .I(N__3221));
    Odrv12 I__490 (
            .O(N__3221),
            .I(U409_ADDRESS_DECODE_un1_nCIACS0_i));
    InMux I__489 (
            .O(N__3218),
            .I(\U409_TICK.un2_COUNTER50_1_cry_1 ));
    InMux I__488 (
            .O(N__3215),
            .I(\U409_TICK.un2_COUNTER50_1_cry_2 ));
    InMux I__487 (
            .O(N__3212),
            .I(\U409_TICK.un2_COUNTER50_1_cry_3 ));
    InMux I__486 (
            .O(N__3209),
            .I(\U409_TICK.un2_COUNTER50_1_cry_4 ));
    InMux I__485 (
            .O(N__3206),
            .I(\U409_TICK.un2_COUNTER50_1_cry_5 ));
    InMux I__484 (
            .O(N__3203),
            .I(\U409_TICK.un2_COUNTER50_1_cry_6 ));
    InMux I__483 (
            .O(N__3200),
            .I(bfn_8_9_0_));
    InMux I__482 (
            .O(N__3197),
            .I(\U409_TICK.un3_COUNTER60_1_cry_9 ));
    InMux I__481 (
            .O(N__3194),
            .I(N__3191));
    LocalMux I__480 (
            .O(N__3191),
            .I(N__3187));
    InMux I__479 (
            .O(N__3190),
            .I(N__3184));
    Odrv4 I__478 (
            .O(N__3187),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    LocalMux I__477 (
            .O(N__3184),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    InMux I__476 (
            .O(N__3179),
            .I(\U409_TICK.un3_COUNTER60_1_cry_10 ));
    InMux I__475 (
            .O(N__3176),
            .I(N__3173));
    LocalMux I__474 (
            .O(N__3173),
            .I(N__3169));
    InMux I__473 (
            .O(N__3172),
            .I(N__3166));
    Odrv4 I__472 (
            .O(N__3169),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    LocalMux I__471 (
            .O(N__3166),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    InMux I__470 (
            .O(N__3161),
            .I(\U409_TICK.un3_COUNTER60_1_cry_11 ));
    InMux I__469 (
            .O(N__3158),
            .I(\U409_TICK.un3_COUNTER60_1_cry_12 ));
    InMux I__468 (
            .O(N__3155),
            .I(\U409_TICK.un3_COUNTER60_1_cry_13 ));
    InMux I__467 (
            .O(N__3152),
            .I(\U409_TICK.un3_COUNTER60_1_cry_14 ));
    InMux I__466 (
            .O(N__3149),
            .I(\U409_TICK.un3_COUNTER60_1_cry_15 ));
    InMux I__465 (
            .O(N__3146),
            .I(N__3143));
    LocalMux I__464 (
            .O(N__3143),
            .I(N__3139));
    InMux I__463 (
            .O(N__3142),
            .I(N__3136));
    Span4Mux_h I__462 (
            .O(N__3139),
            .I(N__3133));
    LocalMux I__461 (
            .O(N__3136),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    Odrv4 I__460 (
            .O(N__3133),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    InMux I__459 (
            .O(N__3128),
            .I(N__3125));
    LocalMux I__458 (
            .O(N__3125),
            .I(N__3121));
    InMux I__457 (
            .O(N__3124),
            .I(N__3118));
    Odrv12 I__456 (
            .O(N__3121),
            .I(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0 ));
    LocalMux I__455 (
            .O(N__3118),
            .I(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0 ));
    IoInMux I__454 (
            .O(N__3113),
            .I(N__3110));
    LocalMux I__453 (
            .O(N__3110),
            .I(N__3107));
    IoSpan4Mux I__452 (
            .O(N__3107),
            .I(N__3104));
    IoSpan4Mux I__451 (
            .O(N__3104),
            .I(N__3101));
    Span4Mux_s2_v I__450 (
            .O(N__3101),
            .I(N__3098));
    Sp12to4 I__449 (
            .O(N__3098),
            .I(N__3095));
    Span12Mux_v I__448 (
            .O(N__3095),
            .I(N__3092));
    Odrv12 I__447 (
            .O(N__3092),
            .I(nBUFEN_c));
    CascadeMux I__446 (
            .O(N__3089),
            .I(N__3085));
    CascadeMux I__445 (
            .O(N__3088),
            .I(N__3082));
    InMux I__444 (
            .O(N__3085),
            .I(N__3076));
    InMux I__443 (
            .O(N__3082),
            .I(N__3076));
    InMux I__442 (
            .O(N__3081),
            .I(N__3073));
    LocalMux I__441 (
            .O(N__3076),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__440 (
            .O(N__3073),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    CascadeMux I__439 (
            .O(N__3068),
            .I(N__3062));
    InMux I__438 (
            .O(N__3067),
            .I(N__3055));
    InMux I__437 (
            .O(N__3066),
            .I(N__3055));
    InMux I__436 (
            .O(N__3065),
            .I(N__3055));
    InMux I__435 (
            .O(N__3062),
            .I(N__3052));
    LocalMux I__434 (
            .O(N__3055),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__433 (
            .O(N__3052),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    InMux I__432 (
            .O(N__3047),
            .I(N__3043));
    InMux I__431 (
            .O(N__3046),
            .I(N__3040));
    LocalMux I__430 (
            .O(N__3043),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    LocalMux I__429 (
            .O(N__3040),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    InMux I__428 (
            .O(N__3035),
            .I(\U409_TICK.un3_COUNTER60_1_cry_1 ));
    InMux I__427 (
            .O(N__3032),
            .I(N__3028));
    InMux I__426 (
            .O(N__3031),
            .I(N__3025));
    LocalMux I__425 (
            .O(N__3028),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    LocalMux I__424 (
            .O(N__3025),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    InMux I__423 (
            .O(N__3020),
            .I(\U409_TICK.un3_COUNTER60_1_cry_2 ));
    InMux I__422 (
            .O(N__3017),
            .I(N__3013));
    InMux I__421 (
            .O(N__3016),
            .I(N__3010));
    LocalMux I__420 (
            .O(N__3013),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    LocalMux I__419 (
            .O(N__3010),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    InMux I__418 (
            .O(N__3005),
            .I(N__3002));
    LocalMux I__417 (
            .O(N__3002),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ));
    InMux I__416 (
            .O(N__2999),
            .I(\U409_TICK.un3_COUNTER60_1_cry_3 ));
    InMux I__415 (
            .O(N__2996),
            .I(N__2992));
    InMux I__414 (
            .O(N__2995),
            .I(N__2989));
    LocalMux I__413 (
            .O(N__2992),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    LocalMux I__412 (
            .O(N__2989),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    InMux I__411 (
            .O(N__2984),
            .I(\U409_TICK.un3_COUNTER60_1_cry_4 ));
    InMux I__410 (
            .O(N__2981),
            .I(N__2978));
    LocalMux I__409 (
            .O(N__2978),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ));
    InMux I__408 (
            .O(N__2975),
            .I(\U409_TICK.un3_COUNTER60_1_cry_5 ));
    InMux I__407 (
            .O(N__2972),
            .I(\U409_TICK.un3_COUNTER60_1_cry_6 ));
    InMux I__406 (
            .O(N__2969),
            .I(\U409_TICK.un3_COUNTER60_1_cry_7 ));
    InMux I__405 (
            .O(N__2966),
            .I(N__2962));
    InMux I__404 (
            .O(N__2965),
            .I(N__2959));
    LocalMux I__403 (
            .O(N__2962),
            .I(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3 ));
    LocalMux I__402 (
            .O(N__2959),
            .I(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3 ));
    InMux I__401 (
            .O(N__2954),
            .I(N__2944));
    InMux I__400 (
            .O(N__2953),
            .I(N__2944));
    InMux I__399 (
            .O(N__2952),
            .I(N__2941));
    InMux I__398 (
            .O(N__2951),
            .I(N__2936));
    InMux I__397 (
            .O(N__2950),
            .I(N__2936));
    InMux I__396 (
            .O(N__2949),
            .I(N__2933));
    LocalMux I__395 (
            .O(N__2944),
            .I(N__2928));
    LocalMux I__394 (
            .O(N__2941),
            .I(N__2928));
    LocalMux I__393 (
            .O(N__2936),
            .I(N__2925));
    LocalMux I__392 (
            .O(N__2933),
            .I(N__2922));
    Span4Mux_v I__391 (
            .O(N__2928),
            .I(N__2919));
    Span4Mux_v I__390 (
            .O(N__2925),
            .I(N__2916));
    Span4Mux_v I__389 (
            .O(N__2922),
            .I(N__2913));
    Sp12to4 I__388 (
            .O(N__2919),
            .I(N__2910));
    Span4Mux_h I__387 (
            .O(N__2916),
            .I(N__2907));
    Span4Mux_h I__386 (
            .O(N__2913),
            .I(N__2904));
    Odrv12 I__385 (
            .O(N__2910),
            .I(A_c_23));
    Odrv4 I__384 (
            .O(N__2907),
            .I(A_c_23));
    Odrv4 I__383 (
            .O(N__2904),
            .I(A_c_23));
    IoInMux I__382 (
            .O(N__2897),
            .I(N__2894));
    LocalMux I__381 (
            .O(N__2894),
            .I(N__2891));
    IoSpan4Mux I__380 (
            .O(N__2891),
            .I(N__2888));
    Span4Mux_s2_v I__379 (
            .O(N__2888),
            .I(N__2885));
    Sp12to4 I__378 (
            .O(N__2885),
            .I(N__2882));
    Span12Mux_v I__377 (
            .O(N__2882),
            .I(N__2879));
    Span12Mux_h I__376 (
            .O(N__2879),
            .I(N__2876));
    Odrv12 I__375 (
            .O(N__2876),
            .I(U409_ADDRESS_DECODE_un1_nREGSPACE_i));
    InMux I__374 (
            .O(N__2873),
            .I(N__2870));
    LocalMux I__373 (
            .O(N__2870),
            .I(N__2867));
    Odrv12 I__372 (
            .O(N__2867),
            .I(\U409_ADDRESS_DECODE.un10_ROMENZ0 ));
    InMux I__371 (
            .O(N__2864),
            .I(N__2861));
    LocalMux I__370 (
            .O(N__2861),
            .I(\U409_TICK.TICK603_8 ));
    CascadeMux I__369 (
            .O(N__2858),
            .I(\U409_TICK.TICK603_11_cascade_ ));
    CascadeMux I__368 (
            .O(N__2855),
            .I(\U409_TICK.TICK603_14_cascade_ ));
    InMux I__367 (
            .O(N__2852),
            .I(N__2846));
    InMux I__366 (
            .O(N__2851),
            .I(N__2846));
    LocalMux I__365 (
            .O(N__2846),
            .I(N__2843));
    Span4Mux_h I__364 (
            .O(N__2843),
            .I(N__2840));
    Span4Mux_v I__363 (
            .O(N__2840),
            .I(N__2837));
    Odrv4 I__362 (
            .O(N__2837),
            .I(A_c_29));
    InMux I__361 (
            .O(N__2834),
            .I(N__2831));
    LocalMux I__360 (
            .O(N__2831),
            .I(\U409_CIA.g0Z0Z_2 ));
    InMux I__359 (
            .O(N__2828),
            .I(N__2822));
    InMux I__358 (
            .O(N__2827),
            .I(N__2822));
    LocalMux I__357 (
            .O(N__2822),
            .I(N__2819));
    Span4Mux_v I__356 (
            .O(N__2819),
            .I(N__2816));
    Sp12to4 I__355 (
            .O(N__2816),
            .I(N__2813));
    Odrv12 I__354 (
            .O(N__2813),
            .I(A_c_31));
    InMux I__353 (
            .O(N__2810),
            .I(N__2804));
    InMux I__352 (
            .O(N__2809),
            .I(N__2804));
    LocalMux I__351 (
            .O(N__2804),
            .I(N__2801));
    Span4Mux_v I__350 (
            .O(N__2801),
            .I(N__2798));
    Sp12to4 I__349 (
            .O(N__2798),
            .I(N__2795));
    Odrv12 I__348 (
            .O(N__2795),
            .I(A_c_30));
    InMux I__347 (
            .O(N__2792),
            .I(N__2789));
    LocalMux I__346 (
            .O(N__2789),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3 ));
    InMux I__345 (
            .O(N__2786),
            .I(N__2780));
    InMux I__344 (
            .O(N__2785),
            .I(N__2773));
    InMux I__343 (
            .O(N__2784),
            .I(N__2773));
    InMux I__342 (
            .O(N__2783),
            .I(N__2773));
    LocalMux I__341 (
            .O(N__2780),
            .I(N__2770));
    LocalMux I__340 (
            .O(N__2773),
            .I(N__2767));
    Span4Mux_v I__339 (
            .O(N__2770),
            .I(N__2764));
    Span12Mux_v I__338 (
            .O(N__2767),
            .I(N__2761));
    Sp12to4 I__337 (
            .O(N__2764),
            .I(N__2758));
    Odrv12 I__336 (
            .O(N__2761),
            .I(A_c_21));
    Odrv12 I__335 (
            .O(N__2758),
            .I(A_c_21));
    InMux I__334 (
            .O(N__2753),
            .I(N__2750));
    LocalMux I__333 (
            .O(N__2750),
            .I(N__2747));
    Span4Mux_v I__332 (
            .O(N__2747),
            .I(N__2742));
    InMux I__331 (
            .O(N__2746),
            .I(N__2737));
    InMux I__330 (
            .O(N__2745),
            .I(N__2737));
    Sp12to4 I__329 (
            .O(N__2742),
            .I(N__2732));
    LocalMux I__328 (
            .O(N__2737),
            .I(N__2732));
    Odrv12 I__327 (
            .O(N__2732),
            .I(A_c_20));
    CascadeMux I__326 (
            .O(N__2729),
            .I(N__2726));
    InMux I__325 (
            .O(N__2726),
            .I(N__2720));
    InMux I__324 (
            .O(N__2725),
            .I(N__2720));
    LocalMux I__323 (
            .O(N__2720),
            .I(N__2717));
    Odrv4 I__322 (
            .O(N__2717),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEm_6 ));
    CascadeMux I__321 (
            .O(N__2714),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2_cascade_ ));
    InMux I__320 (
            .O(N__2711),
            .I(N__2706));
    InMux I__319 (
            .O(N__2710),
            .I(N__2701));
    InMux I__318 (
            .O(N__2709),
            .I(N__2701));
    LocalMux I__317 (
            .O(N__2706),
            .I(N__2698));
    LocalMux I__316 (
            .O(N__2701),
            .I(N__2695));
    Span4Mux_v I__315 (
            .O(N__2698),
            .I(N__2692));
    Span4Mux_h I__314 (
            .O(N__2695),
            .I(N__2689));
    Sp12to4 I__313 (
            .O(N__2692),
            .I(N__2686));
    Span4Mux_v I__312 (
            .O(N__2689),
            .I(N__2683));
    Span12Mux_h I__311 (
            .O(N__2686),
            .I(N__2680));
    Span4Mux_v I__310 (
            .O(N__2683),
            .I(N__2677));
    Span12Mux_v I__309 (
            .O(N__2680),
            .I(N__2674));
    Span4Mux_v I__308 (
            .O(N__2677),
            .I(N__2671));
    Odrv12 I__307 (
            .O(N__2674),
            .I(A_c_19));
    Odrv4 I__306 (
            .O(N__2671),
            .I(A_c_19));
    CascadeMux I__305 (
            .O(N__2666),
            .I(N__2661));
    CascadeMux I__304 (
            .O(N__2665),
            .I(N__2657));
    InMux I__303 (
            .O(N__2664),
            .I(N__2653));
    InMux I__302 (
            .O(N__2661),
            .I(N__2644));
    InMux I__301 (
            .O(N__2660),
            .I(N__2644));
    InMux I__300 (
            .O(N__2657),
            .I(N__2644));
    InMux I__299 (
            .O(N__2656),
            .I(N__2644));
    LocalMux I__298 (
            .O(N__2653),
            .I(N__2641));
    LocalMux I__297 (
            .O(N__2644),
            .I(N__2636));
    Sp12to4 I__296 (
            .O(N__2641),
            .I(N__2636));
    Span12Mux_v I__295 (
            .O(N__2636),
            .I(N__2633));
    Odrv12 I__294 (
            .O(N__2633),
            .I(A_c_22));
    InMux I__293 (
            .O(N__2630),
            .I(N__2627));
    LocalMux I__292 (
            .O(N__2627),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2 ));
    InMux I__291 (
            .O(N__2624),
            .I(N__2621));
    LocalMux I__290 (
            .O(N__2621),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3 ));
    IoInMux I__289 (
            .O(N__2618),
            .I(N__2615));
    LocalMux I__288 (
            .O(N__2615),
            .I(N__2612));
    Span4Mux_s0_v I__287 (
            .O(N__2612),
            .I(N__2609));
    Span4Mux_v I__286 (
            .O(N__2609),
            .I(N__2606));
    Span4Mux_v I__285 (
            .O(N__2606),
            .I(N__2603));
    Span4Mux_v I__284 (
            .O(N__2603),
            .I(N__2600));
    Odrv4 I__283 (
            .O(N__2600),
            .I(PORTSIZE_0_i));
    CascadeMux I__282 (
            .O(N__2597),
            .I(N__2594));
    InMux I__281 (
            .O(N__2594),
            .I(N__2588));
    InMux I__280 (
            .O(N__2593),
            .I(N__2588));
    LocalMux I__279 (
            .O(N__2588),
            .I(N__2585));
    Span12Mux_h I__278 (
            .O(N__2585),
            .I(N__2582));
    Span12Mux_v I__277 (
            .O(N__2582),
            .I(N__2579));
    Odrv12 I__276 (
            .O(N__2579),
            .I(A_c_18));
    CascadeMux I__275 (
            .O(N__2576),
            .I(N__2572));
    InMux I__274 (
            .O(N__2575),
            .I(N__2567));
    InMux I__273 (
            .O(N__2572),
            .I(N__2567));
    LocalMux I__272 (
            .O(N__2567),
            .I(N__2564));
    Span4Mux_v I__271 (
            .O(N__2564),
            .I(N__2561));
    Span4Mux_h I__270 (
            .O(N__2561),
            .I(N__2558));
    Span4Mux_v I__269 (
            .O(N__2558),
            .I(N__2555));
    Span4Mux_v I__268 (
            .O(N__2555),
            .I(N__2552));
    Odrv4 I__267 (
            .O(N__2552),
            .I(A_c_16));
    InMux I__266 (
            .O(N__2549),
            .I(N__2543));
    InMux I__265 (
            .O(N__2548),
            .I(N__2543));
    LocalMux I__264 (
            .O(N__2543),
            .I(N__2540));
    Span12Mux_s5_h I__263 (
            .O(N__2540),
            .I(N__2537));
    Span12Mux_v I__262 (
            .O(N__2537),
            .I(N__2534));
    Odrv12 I__261 (
            .O(N__2534),
            .I(A_c_17));
    CascadeMux I__260 (
            .O(N__2531),
            .I(\U409_CIA.g0Z0Z_11_cascade_ ));
    InMux I__259 (
            .O(N__2528),
            .I(N__2525));
    LocalMux I__258 (
            .O(N__2525),
            .I(N__2522));
    Odrv4 I__257 (
            .O(N__2522),
            .I(\U409_CIA.g0Z0Z_8 ));
    InMux I__256 (
            .O(N__2519),
            .I(N__2516));
    LocalMux I__255 (
            .O(N__2516),
            .I(N__2512));
    InMux I__254 (
            .O(N__2515),
            .I(N__2509));
    Span4Mux_v I__253 (
            .O(N__2512),
            .I(N__2506));
    LocalMux I__252 (
            .O(N__2509),
            .I(N__2503));
    Span4Mux_v I__251 (
            .O(N__2506),
            .I(N__2498));
    Span4Mux_v I__250 (
            .O(N__2503),
            .I(N__2498));
    Sp12to4 I__249 (
            .O(N__2498),
            .I(N__2495));
    Odrv12 I__248 (
            .O(N__2495),
            .I(A_c_25));
    CascadeMux I__247 (
            .O(N__2492),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_ ));
    InMux I__246 (
            .O(N__2489),
            .I(N__2483));
    InMux I__245 (
            .O(N__2488),
            .I(N__2483));
    LocalMux I__244 (
            .O(N__2483),
            .I(N__2480));
    Span4Mux_v I__243 (
            .O(N__2480),
            .I(N__2477));
    Sp12to4 I__242 (
            .O(N__2477),
            .I(N__2474));
    Odrv12 I__241 (
            .O(N__2474),
            .I(A_c_27));
    CascadeMux I__240 (
            .O(N__2471),
            .I(N__2468));
    InMux I__239 (
            .O(N__2468),
            .I(N__2462));
    InMux I__238 (
            .O(N__2467),
            .I(N__2462));
    LocalMux I__237 (
            .O(N__2462),
            .I(N__2459));
    Span4Mux_h I__236 (
            .O(N__2459),
            .I(N__2456));
    Span4Mux_v I__235 (
            .O(N__2456),
            .I(N__2453));
    Odrv4 I__234 (
            .O(N__2453),
            .I(A_c_24));
    CascadeMux I__233 (
            .O(N__2450),
            .I(N__2446));
    InMux I__232 (
            .O(N__2449),
            .I(N__2443));
    InMux I__231 (
            .O(N__2446),
            .I(N__2440));
    LocalMux I__230 (
            .O(N__2443),
            .I(N__2435));
    LocalMux I__229 (
            .O(N__2440),
            .I(N__2435));
    Span4Mux_v I__228 (
            .O(N__2435),
            .I(N__2432));
    Span4Mux_v I__227 (
            .O(N__2432),
            .I(N__2429));
    Span4Mux_h I__226 (
            .O(N__2429),
            .I(N__2426));
    Odrv4 I__225 (
            .O(N__2426),
            .I(A_c_26));
    InMux I__224 (
            .O(N__2423),
            .I(N__2417));
    InMux I__223 (
            .O(N__2422),
            .I(N__2417));
    LocalMux I__222 (
            .O(N__2417),
            .I(N__2414));
    Span4Mux_v I__221 (
            .O(N__2414),
            .I(N__2411));
    Span4Mux_v I__220 (
            .O(N__2411),
            .I(N__2408));
    Sp12to4 I__219 (
            .O(N__2408),
            .I(N__2405));
    Odrv12 I__218 (
            .O(N__2405),
            .I(A_c_28));
    CascadeMux I__217 (
            .O(N__2402),
            .I(\U409_CIA.g0Z0Z_10_cascade_ ));
    ClkMux I__216 (
            .O(N__2399),
            .I(N__2369));
    ClkMux I__215 (
            .O(N__2398),
            .I(N__2369));
    ClkMux I__214 (
            .O(N__2397),
            .I(N__2369));
    ClkMux I__213 (
            .O(N__2396),
            .I(N__2369));
    ClkMux I__212 (
            .O(N__2395),
            .I(N__2369));
    ClkMux I__211 (
            .O(N__2394),
            .I(N__2369));
    ClkMux I__210 (
            .O(N__2393),
            .I(N__2369));
    ClkMux I__209 (
            .O(N__2392),
            .I(N__2369));
    ClkMux I__208 (
            .O(N__2391),
            .I(N__2369));
    ClkMux I__207 (
            .O(N__2390),
            .I(N__2369));
    GlobalMux I__206 (
            .O(N__2369),
            .I(CLK80_OUT));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .I(N__2390));
    INV \INVU409_TRANSFER_ACK.TACK_EN_iC  (
            .O(\INVU409_TRANSFER_ACK.TACK_EN_iC_net ),
            .I(N__2397));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .I(N__2393));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .I(N__2391));
    INV \INVU409_TRANSFER_ACK.TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .I(N__2398));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .I(N__2396));
    INV \INVU409_TRANSFER_ACK.LASTCLK_1C  (
            .O(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .I(N__2394));
    INV \INVU409_TRANSFER_ACK.LASTCLK_0C  (
            .O(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .I(N__2392));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ),
            .I(N__2399));
    INV \INVU409_TRANSFER_ACK.CIA_ENABLED_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .I(N__2395));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_9_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_5_0_));
    defparam IN_MUX_bfv_9_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_6_0_ (
            .carryinitin(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .carryinitout(bfn_9_6_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_7_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_1_10_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_1_10_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_1_10_0  (
            .in0(N__2709),
            .in1(N__2593),
            .in2(N__2576),
            .in3(N__2548),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEm_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_11_LC_1_10_3 .C_ON=1'b0;
    defparam \U409_CIA.g0_11_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_11_LC_1_10_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_CIA.g0_11_LC_1_10_3  (
            .in0(N__2519),
            .in1(N__2710),
            .in2(N__2597),
            .in3(N__2575),
            .lcout(),
            .ltout(\U409_CIA.g0Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_14_LC_1_10_4 .C_ON=1'b0;
    defparam \U409_CIA.g0_14_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_14_LC_1_10_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_CIA.g0_14_LC_1_10_4  (
            .in0(N__2753),
            .in1(N__2549),
            .in2(N__2531),
            .in3(N__2528),
            .lcout(\U409_CIA.g0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_8_LC_1_12_3 .C_ON=1'b0;
    defparam \U409_CIA.g0_8_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_8_LC_1_12_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_CIA.g0_8_LC_1_12_3  (
            .in0(N__5611),
            .in1(N__2949),
            .in2(_gnd_net_),
            .in3(N__2786),
            .lcout(\U409_CIA.g0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_0  (
            .in0(N__2467),
            .in1(N__2488),
            .in2(N__2450),
            .in3(N__2515),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_1  (
            .in0(N__2851),
            .in1(N__2422),
            .in2(N__2492),
            .in3(N__2792),
            .lcout(U409_ADDRESS_DECODE_Z2_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_10_LC_1_17_2 .C_ON=1'b0;
    defparam \U409_CIA.g0_10_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_10_LC_1_17_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_CIA.g0_10_LC_1_17_2  (
            .in0(N__2828),
            .in1(N__2489),
            .in2(N__2471),
            .in3(N__2449),
            .lcout(),
            .ltout(\U409_CIA.g0Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_13_LC_1_17_3 .C_ON=1'b0;
    defparam \U409_CIA.g0_13_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_13_LC_1_17_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_CIA.g0_13_LC_1_17_3  (
            .in0(N__2664),
            .in1(N__2423),
            .in2(N__2402),
            .in3(N__2834),
            .lcout(\U409_CIA.g0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_2_LC_1_17_4 .C_ON=1'b0;
    defparam \U409_CIA.g0_2_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_2_LC_1_17_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_CIA.g0_2_LC_1_17_4  (
            .in0(N__2810),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2852),
            .lcout(\U409_CIA.g0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_17_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_17_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_17_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_17_7  (
            .in0(_gnd_net_),
            .in1(N__2827),
            .in2(_gnd_net_),
            .in3(N__2809),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_2_12_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_2_12_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_2_12_0  (
            .in0(N__2784),
            .in1(N__2660),
            .in2(N__2729),
            .in3(N__2746),
            .lcout(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un6_ROMEN_LC_2_12_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un6_ROMEN_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un6_ROMEN_LC_2_12_1 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \U409_ADDRESS_DECODE.un6_ROMEN_LC_2_12_1  (
            .in0(N__2951),
            .in1(_gnd_net_),
            .in2(N__2666),
            .in3(N__2785),
            .lcout(\U409_ADDRESS_DECODE.un6_ROMENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_2_12_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_2_12_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_2_12_4  (
            .in0(N__2783),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2745),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2 ),
            .ltout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_2_12_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_2_12_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_2_12_5  (
            .in0(N__2656),
            .in1(N__2725),
            .in2(N__2714),
            .in3(N__5322),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un10_ROMEN_LC_2_12_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un10_ROMEN_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un10_ROMEN_LC_2_12_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un10_ROMEN_LC_2_12_7  (
            .in0(N__2950),
            .in1(N__2711),
            .in2(N__2665),
            .in3(N__2630),
            .lcout(\U409_ADDRESS_DECODE.un10_ROMENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_3_12_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_3_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_3_12_0 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_3_12_0  (
            .in0(N__2953),
            .in1(N__3124),
            .in2(N__5612),
            .in3(N__2624),
            .lcout(PORTSIZE_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_3_12_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_3_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_3_12_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_3_12_7  (
            .in0(N__2965),
            .in1(N__2954),
            .in2(_gnd_net_),
            .in3(N__5345),
            .lcout(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_3_13_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_3_13_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_3_13_7 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_3_13_7  (
            .in0(N__2966),
            .in1(N__2952),
            .in2(_gnd_net_),
            .in3(N__5326),
            .lcout(U409_ADDRESS_DECODE_un1_nREGSPACE_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_ROMEN_LC_7_12_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_ROMEN_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_ROMEN_LC_7_12_2 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \U409_ADDRESS_DECODE.un1_ROMEN_LC_7_12_2  (
            .in0(N__4871),
            .in1(N__2873),
            .in2(_gnd_net_),
            .in3(N__4818),
            .lcout(U409_ADDRESS_DECODE_un1_ROMEN_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_8_7_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_8_7_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_TICK.COUNTER60_RNIHJU51_4_LC_8_7_0  (
            .in0(N__2996),
            .in1(N__3017),
            .in2(_gnd_net_),
            .in3(N__3065),
            .lcout(\U409_TICK.TICK603_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_4_LC_8_7_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_4_LC_8_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_4_LC_8_7_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_4_LC_8_7_2  (
            .in0(N__3431),
            .in1(N__3404),
            .in2(N__3378),
            .in3(N__3005),
            .lcout(\U409_TICK.COUNTER60Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4172),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_1_LC_8_7_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_1_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_1_LC_8_7_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER60_1_LC_8_7_3  (
            .in0(N__3067),
            .in1(_gnd_net_),
            .in2(N__3089),
            .in3(_gnd_net_),
            .lcout(\U409_TICK.COUNTER60Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4172),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_6_LC_8_7_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_6_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_6_LC_8_7_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_6_LC_8_7_4  (
            .in0(N__3432),
            .in1(N__3405),
            .in2(N__3379),
            .in3(N__2981),
            .lcout(\U409_TICK.COUNTER60Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4172),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_8_7_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_8_7_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER60_RNIDB4S_16_LC_8_7_5  (
            .in0(N__3176),
            .in1(N__3047),
            .in2(N__3088),
            .in3(N__3146),
            .lcout(),
            .ltout(\U409_TICK.TICK603_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_8_7_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_8_7_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER60_RNI335G2_11_LC_8_7_6  (
            .in0(N__2864),
            .in1(N__3194),
            .in2(N__2858),
            .in3(N__3032),
            .lcout(\U409_TICK.TICK603_14 ),
            .ltout(\U409_TICK.TICK603_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_0_LC_8_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_0_LC_8_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_0_LC_8_7_7 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \U409_TICK.COUNTER60_0_LC_8_7_7  (
            .in0(N__3066),
            .in1(N__3433),
            .in2(N__2855),
            .in3(N__3371),
            .lcout(\U409_TICK.COUNTER60Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4172),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_8_8_0 .C_ON=1'b1;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_8_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__3081),
            .in2(N__3068),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_2_LC_8_8_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_2_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_2_LC_8_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_2_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(N__3046),
            .in2(_gnd_net_),
            .in3(N__3035),
            .lcout(\U409_TICK.COUNTER60Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .clk(N__4174),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_3_LC_8_8_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_3_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_3_LC_8_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_3_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__3031),
            .in2(_gnd_net_),
            .in3(N__3020),
            .lcout(\U409_TICK.COUNTER60Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .clk(N__4174),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_8_8_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_8_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_4_LC_8_8_3  (
            .in0(_gnd_net_),
            .in1(N__3016),
            .in2(_gnd_net_),
            .in3(N__2999),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_5_LC_8_8_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_5_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_5_LC_8_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_5_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(N__2995),
            .in2(_gnd_net_),
            .in3(N__2984),
            .lcout(\U409_TICK.COUNTER60Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .clk(N__4174),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_8_8_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_8_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_6_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(N__3538),
            .in2(_gnd_net_),
            .in3(N__2975),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_7_LC_8_8_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_7_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_7_LC_8_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_7_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(N__3466),
            .in2(_gnd_net_),
            .in3(N__2972),
            .lcout(\U409_TICK.COUNTER60Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .clk(N__4174),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_8_8_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_8_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_8_LC_8_8_7  (
            .in0(_gnd_net_),
            .in1(N__3505),
            .in2(_gnd_net_),
            .in3(N__2969),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_8_9_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_8_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_9_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__3550),
            .in2(_gnd_net_),
            .in3(N__3200),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_10_LC_8_9_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_10_LC_8_9_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_10_LC_8_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_10_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__3481),
            .in2(_gnd_net_),
            .in3(N__3197),
            .lcout(\U409_TICK.COUNTER60Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .clk(N__4175),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_11_LC_8_9_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_11_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_11_LC_8_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_11_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__3190),
            .in2(_gnd_net_),
            .in3(N__3179),
            .lcout(\U409_TICK.COUNTER60Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .clk(N__4175),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_12_LC_8_9_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_12_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_12_LC_8_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_12_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__3172),
            .in2(_gnd_net_),
            .in3(N__3161),
            .lcout(\U409_TICK.COUNTER60Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .clk(N__4175),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_13_LC_8_9_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_13_LC_8_9_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_13_LC_8_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_13_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__3493),
            .in2(_gnd_net_),
            .in3(N__3158),
            .lcout(\U409_TICK.COUNTER60Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .clk(N__4175),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_8_9_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_8_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_14_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(N__3331),
            .in2(_gnd_net_),
            .in3(N__3155),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_8_9_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_8_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_15_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__3454),
            .in2(_gnd_net_),
            .in3(N__3152),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_16_LC_8_9_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_16_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_16_LC_8_9_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER60_16_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(N__3142),
            .in2(_gnd_net_),
            .in3(N__3149),
            .lcout(\U409_TICK.COUNTER60Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4175),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_8_12_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_8_12_0 .LUT_INIT=16'b0011001100010011;
    LogicCell40 \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_8_12_0  (
            .in0(N__5335),
            .in1(N__3128),
            .in2(N__4825),
            .in3(N__4867),
            .lcout(nBUFEN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_9_4_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_9_4_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_9_4_2  (
            .in0(_gnd_net_),
            .in1(N__3293),
            .in2(_gnd_net_),
            .in3(N__3737),
            .lcout(U409_ADDRESS_DECODE_un1_nCIACS1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_9_4_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_9_4_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_9_4_3  (
            .in0(N__3736),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3254),
            .lcout(U409_ADDRESS_DECODE_un1_nCIACS0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_9_5_0 .C_ON=1'b1;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_9_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_9_5_0  (
            .in0(_gnd_net_),
            .in1(N__3781),
            .in2(N__3884),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_5_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_2_LC_9_5_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_2_LC_9_5_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_2_LC_9_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_2_LC_9_5_1  (
            .in0(_gnd_net_),
            .in1(N__3802),
            .in2(_gnd_net_),
            .in3(N__3218),
            .lcout(\U409_TICK.COUNTER50Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .clk(N__4168),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_3_LC_9_5_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_3_LC_9_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_3_LC_9_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_3_LC_9_5_2  (
            .in0(_gnd_net_),
            .in1(N__3925),
            .in2(_gnd_net_),
            .in3(N__3215),
            .lcout(\U409_TICK.COUNTER50Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .clk(N__4168),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_4_LC_9_5_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_4_LC_9_5_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_4_LC_9_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_4_LC_9_5_3  (
            .in0(_gnd_net_),
            .in1(N__3862),
            .in2(_gnd_net_),
            .in3(N__3212),
            .lcout(\U409_TICK.COUNTER50Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .clk(N__4168),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_9_5_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_9_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_5_LC_9_5_4  (
            .in0(_gnd_net_),
            .in1(N__3826),
            .in2(_gnd_net_),
            .in3(N__3209),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_9_5_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_9_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_6_LC_9_5_5  (
            .in0(_gnd_net_),
            .in1(N__4012),
            .in2(_gnd_net_),
            .in3(N__3206),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_7_LC_9_5_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_7_LC_9_5_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_7_LC_9_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_7_LC_9_5_6  (
            .in0(_gnd_net_),
            .in1(N__3847),
            .in2(_gnd_net_),
            .in3(N__3203),
            .lcout(\U409_TICK.COUNTER50Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .clk(N__4168),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_8_LC_9_5_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_8_LC_9_5_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_8_LC_9_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_8_LC_9_5_7  (
            .in0(_gnd_net_),
            .in1(N__3814),
            .in2(_gnd_net_),
            .in3(N__3320),
            .lcout(\U409_TICK.COUNTER50Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .clk(N__4168),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_9_6_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_9_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_9_LC_9_6_0  (
            .in0(_gnd_net_),
            .in1(N__4190),
            .in2(_gnd_net_),
            .in3(N__3317),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_9_6_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_10_LC_9_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_10_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_10_LC_9_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_10_LC_9_6_1  (
            .in0(_gnd_net_),
            .in1(N__3898),
            .in2(_gnd_net_),
            .in3(N__3314),
            .lcout(\U409_TICK.COUNTER50Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .clk(N__4170),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_9_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_9_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_11_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(N__3979),
            .in2(_gnd_net_),
            .in3(N__3311),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_12_LC_9_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_12_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_12_LC_9_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_12_LC_9_6_3  (
            .in0(_gnd_net_),
            .in1(N__3913),
            .in2(_gnd_net_),
            .in3(N__3308),
            .lcout(\U409_TICK.COUNTER50Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .clk(N__4170),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_9_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_9_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_13_LC_9_6_4  (
            .in0(_gnd_net_),
            .in1(N__4000),
            .in2(_gnd_net_),
            .in3(N__3305),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_9_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_9_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_14_LC_9_6_5  (
            .in0(_gnd_net_),
            .in1(N__3961),
            .in2(_gnd_net_),
            .in3(N__3302),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_9_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_9_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_15_LC_9_6_6  (
            .in0(_gnd_net_),
            .in1(N__3940),
            .in2(_gnd_net_),
            .in3(N__3299),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_16_LC_9_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_16_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_16_LC_9_6_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER50_16_LC_9_6_7  (
            .in0(_gnd_net_),
            .in1(N__3770),
            .in2(_gnd_net_),
            .in3(N__3296),
            .lcout(\U409_TICK.COUNTER50Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4170),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK60_LC_9_7_4 .C_ON=1'b0;
    defparam \U409_TICK.TICK60_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK60_LC_9_7_4 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \U409_TICK.TICK60_LC_9_7_4  (
            .in0(N__3430),
            .in1(N__3571),
            .in2(N__3380),
            .in3(N__3406),
            .lcout(TICK60_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4171),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_9_LC_9_8_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_9_LC_9_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_9_LC_9_8_1 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_9_LC_9_8_1  (
            .in0(N__3410),
            .in1(N__3443),
            .in2(N__3560),
            .in3(N__3374),
            .lcout(\U409_TICK.COUNTER60Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4173),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_9_8_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_9_8_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER60_RNICDC71_14_LC_9_8_2  (
            .in0(N__3551),
            .in1(N__3539),
            .in2(N__3509),
            .in3(N__3332),
            .lcout(\U409_TICK.TICK603_9 ),
            .ltout(\U409_TICK.TICK603_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_15_LC_9_8_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_15_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_15_LC_9_8_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_15_LC_9_8_3  (
            .in0(N__3408),
            .in1(N__3441),
            .in2(N__3527),
            .in3(N__3524),
            .lcout(\U409_TICK.COUNTER60Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4173),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_8_LC_9_8_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_8_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_8_LC_9_8_5 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_8_LC_9_8_5  (
            .in0(N__3409),
            .in1(N__3442),
            .in2(N__3518),
            .in3(N__3373),
            .lcout(\U409_TICK.COUNTER60Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4173),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_9_8_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_9_8_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_TICK.COUNTER60_RNI2USG_10_LC_9_8_6  (
            .in0(N__3494),
            .in1(N__3482),
            .in2(N__3470),
            .in3(N__3455),
            .lcout(\U409_TICK.TICK603_10 ),
            .ltout(\U409_TICK.TICK603_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_14_LC_9_8_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_14_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_14_LC_9_8_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_14_LC_9_8_7  (
            .in0(N__3407),
            .in1(N__3372),
            .in2(N__3341),
            .in3(N__3338),
            .lcout(\U409_TICK.COUNTER60Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4173),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_RNO_0_LC_9_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_RNO_0_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_RNO_0_LC_9_9_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_RNO_0_LC_9_9_0  (
            .in0(N__5562),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.RESETn_c_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_9_9_1 .C_ON=1'b0;
    defparam \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_9_9_1 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_9_9_1  (
            .in0(N__3707),
            .in1(N__4492),
            .in2(N__3683),
            .in3(N__3721),
            .lcout(CIA_ENABLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_HOLD_LC_9_9_5 .C_ON=1'b0;
    defparam \U409_CIA.CIA_HOLD_LC_9_9_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_HOLD_LC_9_9_5 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U409_CIA.CIA_HOLD_LC_9_9_5  (
            .in0(N__3706),
            .in1(N__4491),
            .in2(N__3682),
            .in3(N__3720),
            .lcout(\U409_CIA.CIA_HOLDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4623),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_9_10_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_9_10_4 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_9_10_4  (
            .in0(N__3725),
            .in1(N__3697),
            .in2(N__4496),
            .in3(N__3670),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .ce(),
            .sr(N__3647));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_9_12_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_9_12_0 .LUT_INIT=16'b1100110000010011;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_9_12_0  (
            .in0(N__3596),
            .in1(N__3630),
            .in2(N__4969),
            .in3(N__3610),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_9_12_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_9_12_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_9_12_1 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_LC_9_12_1  (
            .in0(N__3612),
            .in1(N__5592),
            .in2(N__3638),
            .in3(N__4421),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_9_12_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_9_12_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_9_12_2  (
            .in0(N__3595),
            .in1(N__3629),
            .in2(N__4968),
            .in3(N__3611),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_9_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_9_12_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_9_12_3 .LUT_INIT=16'b0100000011001000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_9_12_3  (
            .in0(N__3613),
            .in1(N__5590),
            .in2(N__3635),
            .in3(N__3631),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_9_12_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_9_12_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_9_12_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_9_12_7  (
            .in0(N__3614),
            .in1(N__5591),
            .in2(_gnd_net_),
            .in3(N__3632),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa_0_LC_9_13_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa_0_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa_0_LC_9_13_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxa_0_LC_9_13_0  (
            .in0(N__5349),
            .in1(N__5266),
            .in2(N__5604),
            .in3(N__5004),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_EN_0_sqmuxaZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_10_5_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_10_5_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_TICK.COUNTER50_RNID6CP_3_LC_10_5_0  (
            .in0(N__3827),
            .in1(N__3926),
            .in2(_gnd_net_),
            .in3(N__3881),
            .lcout(),
            .ltout(\U409_TICK.TICK503_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_10_5_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_10_5_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_10_5_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER50_RNITU182_10_LC_10_5_1  (
            .in0(N__3758),
            .in1(N__3914),
            .in2(N__3902),
            .in3(N__3899),
            .lcout(\U409_TICK.TICK503_14 ),
            .ltout(\U409_TICK.TICK503_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_0_LC_10_5_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_0_LC_10_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_0_LC_10_5_2 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \U409_TICK.COUNTER50_0_LC_10_5_2  (
            .in0(N__4306),
            .in1(N__4233),
            .in2(N__3887),
            .in3(N__3882),
            .lcout(\U409_TICK.COUNTER50Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4166),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_1_LC_10_5_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_1_LC_10_5_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_1_LC_10_5_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER50_1_LC_10_5_3  (
            .in0(N__3883),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3790),
            .lcout(\U409_TICK.COUNTER50Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4166),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_10_5_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_10_5_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_10_5_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNII24V_14_LC_10_5_4  (
            .in0(N__3863),
            .in1(N__3962),
            .in2(N__3851),
            .in3(N__3941),
            .lcout(\U409_TICK.TICK503_10 ),
            .ltout(\U409_TICK.TICK503_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_5_LC_10_5_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_5_LC_10_5_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_5_LC_10_5_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_5_LC_10_5_5  (
            .in0(N__4231),
            .in1(N__4270),
            .in2(N__3836),
            .in3(N__3833),
            .lcout(\U409_TICK.COUNTER50Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4166),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_10_5_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_10_5_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_10_5_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER50_RNIUHF01_16_LC_10_5_6  (
            .in0(N__3815),
            .in1(N__3803),
            .in2(N__3791),
            .in3(N__3769),
            .lcout(\U409_TICK.TICK503_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_6_LC_10_5_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_6_LC_10_5_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_6_LC_10_5_7 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_6_LC_10_5_7  (
            .in0(N__4232),
            .in1(N__4271),
            .in2(N__3752),
            .in3(N__4307),
            .lcout(\U409_TICK.COUNTER50Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4166),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_13_LC_10_6_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_13_LC_10_6_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_13_LC_10_6_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_13_LC_10_6_0  (
            .in0(N__4273),
            .in1(N__4229),
            .in2(N__4318),
            .in3(N__3743),
            .lcout(\U409_TICK.COUNTER50Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4169),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_10_6_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_10_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_10_6_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNIH14V_11_LC_10_6_4  (
            .in0(N__3980),
            .in1(N__4189),
            .in2(N__4016),
            .in3(N__4001),
            .lcout(\U409_TICK.TICK503_9 ),
            .ltout(\U409_TICK.TICK503_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_11_LC_10_6_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_11_LC_10_6_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_11_LC_10_6_5 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \U409_TICK.COUNTER50_11_LC_10_6_5  (
            .in0(N__3989),
            .in1(N__4272),
            .in2(N__3983),
            .in3(N__4308),
            .lcout(\U409_TICK.COUNTER50Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4169),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_14_LC_10_6_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_14_LC_10_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_14_LC_10_6_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_14_LC_10_6_6  (
            .in0(N__4274),
            .in1(N__4230),
            .in2(N__4319),
            .in3(N__3968),
            .lcout(\U409_TICK.COUNTER50Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4169),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_15_LC_10_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_15_LC_10_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_15_LC_10_6_7 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_15_LC_10_6_7  (
            .in0(N__4228),
            .in1(N__4275),
            .in2(N__3950),
            .in3(N__4315),
            .lcout(\U409_TICK.COUNTER50Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4169),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_10_7_5 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_10_7_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_10_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_0_LC_10_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4720),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4625),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_10_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_10_9_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_10_9_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_0_LC_10_9_5  (
            .in0(N__5535),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4642),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_10_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_10_10_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_10_10_0 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_1_LC_10_10_0  (
            .in0(N__4127),
            .in1(_gnd_net_),
            .in2(N__5576),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_10_10_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_10_10_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_10_10_1  (
            .in0(N__4066),
            .in1(N__4136),
            .in2(N__4965),
            .in3(N__4126),
            .lcout(\U409_TRANSFER_ACK.N_97 ),
            .ltout(\U409_TRANSFER_ACK.N_97_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_10_10_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_10_10_2 .LUT_INIT=16'b0000010100100111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_10_10_2  (
            .in0(N__4040),
            .in1(N__4437),
            .in2(N__3929),
            .in3(N__4457),
            .lcout(\U409_TRANSFER_ACK.m9_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_10_10_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_10_10_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(N__4135),
            .in2(_gnd_net_),
            .in3(N__4125),
            .lcout(\U409_TRANSFER_ACK.N_4 ),
            .ltout(\U409_TRANSFER_ACK.N_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_10_10_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_10_10_4 .LUT_INIT=16'b0001000100001111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_10_10_4  (
            .in0(N__4442),
            .in1(N__4458),
            .in2(N__4115),
            .in3(N__4068),
            .lcout(\U409_TRANSFER_ACK.i6_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_10_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_10_10_5 .LUT_INIT=16'b0001101100001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_10_10_5  (
            .in0(N__4067),
            .in1(N__4112),
            .in2(N__4048),
            .in3(N__4097),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.CIA_TACK_EN_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_10_10_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_10_10_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_10_10_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_LC_10_10_6  (
            .in0(N__5537),
            .in1(_gnd_net_),
            .in2(N__4106),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_10_10_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_10_10_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_10_10_7 .LUT_INIT=16'b0000100011001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_1_LC_10_10_7  (
            .in0(N__4069),
            .in1(N__5536),
            .in2(N__4049),
            .in3(N__4103),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIHST5_LC_10_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIHST5_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIHST5_LC_10_11_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNIHST5_LC_10_11_2  (
            .in0(_gnd_net_),
            .in1(N__4882),
            .in2(_gnd_net_),
            .in3(N__4096),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_10_11_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_10_11_3 .LUT_INIT=16'b1111011100000111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_10_11_3  (
            .in0(N__4438),
            .in1(N__4459),
            .in2(N__4047),
            .in3(N__4085),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.m9_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_10_11_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_10_11_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_10_11_4 .LUT_INIT=16'b0010001000001010;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_0_LC_10_11_4  (
            .in0(N__5542),
            .in1(N__4079),
            .in2(N__4073),
            .in3(N__4070),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_10_11_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_10_11_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_10_11_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_10_11_5  (
            .in0(_gnd_net_),
            .in1(N__5541),
            .in2(_gnd_net_),
            .in3(N__4460),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNIURL11_LC_10_12_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNIURL11_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNIURL11_LC_10_12_0 .LUT_INIT=16'b0000010000000101;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNIURL11_LC_10_12_0  (
            .in0(N__4356),
            .in1(N__4420),
            .in2(N__4373),
            .in3(N__4409),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_10_12_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_10_12_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_10_12_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4403),
            .in3(N__5579),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_10_12_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_10_12_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_10_12_5 .LUT_INIT=16'b0000101011101010;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_LC_10_12_5  (
            .in0(N__4384),
            .in1(N__4372),
            .in2(N__5600),
            .in3(N__4778),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_10_12_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_10_12_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_10_12_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_10_12_6  (
            .in0(N__4358),
            .in1(_gnd_net_),
            .in2(N__5599),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_10_12_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_10_12_7 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_10_12_7  (
            .in0(N__5583),
            .in1(N__4371),
            .in2(_gnd_net_),
            .in3(N__4357),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK50_LC_11_5_5 .C_ON=1'b0;
    defparam \U409_TICK.TICK50_LC_11_5_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK50_LC_11_5_5 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \U409_TICK.TICK50_LC_11_5_5  (
            .in0(N__4316),
            .in1(N__4330),
            .in2(N__4241),
            .in3(N__4276),
            .lcout(TICK50_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4165),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_9_LC_11_6_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_9_LC_11_6_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_9_LC_11_6_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_9_LC_11_6_5  (
            .in0(N__4317),
            .in1(N__4277),
            .in2(N__4240),
            .in3(N__4199),
            .lcout(\U409_TICK.COUNTER50Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4167),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_11_7_0 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_11_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__4677),
            .in2(N__4721),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_11_7_1 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_11_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_2_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(N__4559),
            .in2(_gnd_net_),
            .in3(N__4532),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .clk(N__4624),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_11_7_2 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_11_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__4751),
            .in2(_gnd_net_),
            .in3(N__4529),
            .lcout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_11_7_3 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_11_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_4_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(N__4581),
            .in2(_gnd_net_),
            .in3(N__4526),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .clk(N__4624),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_11_7_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_11_7_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(N__4602),
            .in2(_gnd_net_),
            .in3(N__4523),
            .lcout(),
            .ltout(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_11_7_5 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_11_7_5 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_5_LC_11_7_5  (
            .in0(N__4753),
            .in1(N__4507),
            .in2(N__4520),
            .in3(N__4714),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4624),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_11_7_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_11_7_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_11_7_6 .LUT_INIT=16'b0011001101001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_3_LC_11_7_6  (
            .in0(N__4715),
            .in1(N__4517),
            .in2(N__4511),
            .in3(N__4752),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4624),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_11_7_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_11_7_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_11_7_7  (
            .in0(N__4678),
            .in1(N__4582),
            .in2(N__4607),
            .in3(N__4560),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_0_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_0_LC_11_8_0 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_0_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_0_LC_11_8_0 .LUT_INIT=16'b0100010000100010;
    LogicCell40 \U409_CIA.VMA_RNO_0_LC_11_8_0  (
            .in0(N__4755),
            .in1(N__4717),
            .in2(_gnd_net_),
            .in3(N__4680),
            .lcout(),
            .ltout(\U409_CIA.N_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_LC_11_8_1 .C_ON=1'b0;
    defparam \U409_CIA.VMA_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.VMA_LC_11_8_1 .LUT_INIT=16'b0011101010101010;
    LogicCell40 \U409_CIA.VMA_LC_11_8_1  (
            .in0(N__4479),
            .in1(N__4757),
            .in2(N__4499),
            .in3(N__4544),
            .lcout(\U409_CIA.VMAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4622),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_11_8_2 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_11_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_1_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(N__4719),
            .in2(_gnd_net_),
            .in3(N__4681),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4622),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_RNO_1_LC_11_8_3 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_RNO_1_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLKCIA_RNO_1_LC_11_8_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_CIA.CLKCIA_RNO_1_LC_11_8_3  (
            .in0(N__4583),
            .in1(N__4756),
            .in2(N__4606),
            .in3(N__4562),
            .lcout(\U409_CIA.CLKCIA6_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_RNO_2_LC_11_8_4 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_RNO_2_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLKCIA_RNO_2_LC_11_8_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_CIA.CLKCIA_RNO_2_LC_11_8_4  (
            .in0(N__4754),
            .in1(N__4716),
            .in2(_gnd_net_),
            .in3(N__4679),
            .lcout(),
            .ltout(\U409_CIA.N_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_RNO_0_LC_11_8_5 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_RNO_0_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLKCIA_RNO_0_LC_11_8_5 .LUT_INIT=16'b1111110011001100;
    LogicCell40 \U409_CIA.CLKCIA_RNO_0_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(N__4641),
            .in2(N__4730),
            .in3(N__4543),
            .lcout(),
            .ltout(\U409_CIA.CLKCIAZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_LC_11_8_6 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_LC_11_8_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CLKCIA_LC_11_8_6 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \U409_CIA.CLKCIA_LC_11_8_6  (
            .in0(N__4727),
            .in1(N__4718),
            .in2(N__4685),
            .in3(N__4682),
            .lcout(CLKCIA_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4622),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_11_8_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_11_8_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_11_8_7  (
            .in0(N__4598),
            .in1(N__4580),
            .in2(_gnd_net_),
            .in3(N__4561),
            .lcout(\U409_CIA.CLKCIA8_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_9_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_9_0 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_9_0  (
            .in0(N__5149),
            .in1(N__5207),
            .in2(N__5195),
            .in3(N__5101),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__5420));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_9_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_9_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_9_1  (
            .in0(N__5205),
            .in1(N__5100),
            .in2(_gnd_net_),
            .in3(N__5148),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_9_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_9_2 .LUT_INIT=16'b0000001100110000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__5188),
            .in2(N__4535),
            .in3(N__5062),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__5420));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_9_3 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_9_3 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_9_3  (
            .in0(N__5061),
            .in1(N__5078),
            .in2(N__5024),
            .in3(N__5193),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__5420));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_9_5 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_9_5 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_9_5  (
            .in0(N__5618),
            .in1(N__5125),
            .in2(_gnd_net_),
            .in3(N__5192),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__5420));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_11_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_11_9_6 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_11_9_6  (
            .in0(N__4967),
            .in1(N__5008),
            .in2(N__5165),
            .in3(N__5037),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_9_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_9_7 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_9_7  (
            .in0(N__5206),
            .in1(_gnd_net_),
            .in2(N__5015),
            .in3(N__5150),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__5420));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_11_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_11_10_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_11_10_0 .LUT_INIT=16'b0000000001110101;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_11_10_0  (
            .in0(N__5039),
            .in1(N__5012),
            .in2(N__4966),
            .in3(N__5672),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5418));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_10_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_10_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_10_1 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_10_1  (
            .in0(N__4883),
            .in1(N__5038),
            .in2(_gnd_net_),
            .in3(N__5164),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5418));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_11_10_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_11_10_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_11_10_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_11_10_7  (
            .in0(N__5671),
            .in1(N__5641),
            .in2(_gnd_net_),
            .in3(N__5696),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5418));
    defparam \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_11_11_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_11_11_4 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_11_11_4  (
            .in0(N__4860),
            .in1(N__4829),
            .in2(_gnd_net_),
            .in3(N__5351),
            .lcout(U409_ADDRESS_DECODE_un1_nRAMSPACE_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_11_12_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_11_12_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_11_12_5 .LUT_INIT=16'b0111011101110111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_i_LC_11_12_5  (
            .in0(N__5577),
            .in1(N__4777),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(TACK_EN_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_EN_iC_net ),
            .ce(N__4766),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMENm_i_LC_11_13_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMENm_i_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMENm_i_LC_11_13_4 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \U409_ADDRESS_DECODE.ROMENm_i_LC_11_13_4  (
            .in0(N__5350),
            .in1(N__5267),
            .in2(_gnd_net_),
            .in3(N__5578),
            .lcout(ROMENm_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_1_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_1_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_1_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_1_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_12_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_12_9_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_12_9_0  (
            .in0(N__5667),
            .in1(N__5640),
            .in2(N__5126),
            .in3(N__5694),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_12_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_12_9_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_12_9_2 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_12_9_2  (
            .in0(N__5669),
            .in1(N__5695),
            .in2(_gnd_net_),
            .in3(N__5194),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__5419));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_12_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_12_9_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_12_9_3  (
            .in0(N__5124),
            .in1(N__5666),
            .in2(N__5063),
            .in3(N__5076),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_12_9_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_12_9_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_12_9_4  (
            .in0(N__5147),
            .in1(N__5099),
            .in2(N__5168),
            .in3(N__5707),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_12_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_12_9_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_12_9_5  (
            .in0(N__5146),
            .in1(N__5120),
            .in2(N__5102),
            .in3(N__5077),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_12_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_12_9_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_12_9_6  (
            .in0(N__5668),
            .in1(N__5060),
            .in2(N__5042),
            .in3(N__5708),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_12_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_12_10_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(N__5692),
            .in2(_gnd_net_),
            .in3(N__5636),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_12_10_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_12_10_1 .LUT_INIT=16'b1000000010000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_12_10_1  (
            .in0(N__5693),
            .in1(N__5670),
            .in2(N__5642),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_13_10_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_13_10_3 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_13_10_3  (
            .in0(N__5523),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5441),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TACKn_iobuf_RNO_LC_15_15_3.C_ON=1'b0;
    defparam TACKn_iobuf_RNO_LC_15_15_3.SEQ_MODE=4'b0000;
    defparam TACKn_iobuf_RNO_LC_15_15_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 TACKn_iobuf_RNO_LC_15_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5384),
            .lcout(N_347_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U409_TOP

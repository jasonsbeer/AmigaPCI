-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 29 2025 20:48:25

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    CMA : out std_logic_vector(10 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    A : in std_logic_vector(20 downto 0);
    RAMENn : out std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    DBRn : in std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__11587\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10434\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7827\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7434\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7260\ : std_logic;
signal \N__7257\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3959\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3900\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_16\ : std_logic;
signal \N_848_i\ : std_logic;
signal \N_336\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER18_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_371_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0\ : std_logic;
signal \U712_CHIP_RAM.N_321\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.N_371\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \U712_CHIP_RAM.N_285_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_309_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_311\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_55_i_a2_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_212\ : std_logic;
signal \U712_CHIP_RAM.N_326_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0_cascade_\ : std_logic;
signal \A_c_12\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \U712_REG_SM.N_294_cascade_\ : std_logic;
signal \TSn_c\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \U712_CHIP_RAM.LATCH_CLK_8_i_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_368_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_323_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_359_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER15\ : std_logic;
signal \U712_CHIP_RAM.N_330_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_331\ : std_logic;
signal \U712_CHIP_RAM.BANK0_9_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_16\ : std_logic;
signal \U712_CHIP_RAM.N_49_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_55_i_a2_0_a2_0_0\ : std_logic;
signal \A_c_15\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.N_217\ : std_logic;
signal \U712_CHIP_RAM.N_361\ : std_logic;
signal \U712_CHIP_RAM.N_217_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_222\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.N_262\ : std_logic;
signal \U712_CHIP_RAM.N_354_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_408\ : std_logic;
signal \U712_CHIP_RAM.N_408_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_359\ : std_logic;
signal \U712_CHIP_RAM.N_305\ : std_logic;
signal \U712_CYCLE_TERM.N_236_i_0_en_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.N_236_i_0_en_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTc_1_0\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_255\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_srsts_i_0_a2_0_0_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.N_264\ : std_logic;
signal \U712_REG_SM.N_24\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_323\ : std_logic;
signal \U712_CHIP_RAM.N_63\ : std_logic;
signal \LATCH_CLK_c\ : std_logic;
signal \U712_CHIP_RAM.N_363\ : std_logic;
signal \U712_CHIP_RAM.N_363_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_369\ : std_logic;
signal \U712_CHIP_RAM.N_397\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0\ : std_logic;
signal \U712_CHIP_RAM.N_306\ : std_logic;
signal \bfn_10_6_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.N_49\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.N_352_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_328_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un3_DMA_CYCLE_START\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_207\ : std_logic;
signal \U712_CHIP_RAM.CLK_EN_5_0_a2_1_a2_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_370\ : std_logic;
signal \U712_CHIP_RAM.N_307\ : std_logic;
signal \U712_CHIP_RAM.N_411\ : std_logic;
signal \U712_CHIP_RAM.N_403\ : std_logic;
signal \U712_CHIP_RAM.N_411_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_308\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.N_352\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_232\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_REG_SM.N_289\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_254\ : std_logic;
signal \U712_REG_SM.N_254_cascade_\ : std_logic;
signal \U712_REG_SM.N_26\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.N_216\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.N_239\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.N_239_0_0\ : std_logic;
signal \RnW_c\ : std_logic;
signal \WRITE_CYCLEm\ : std_logic;
signal \N_259\ : std_logic;
signal \U712_CHIP_RAM.N_360\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0_0\ : std_logic;
signal \U712_CHIP_RAM.CLK_EN_5_0\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.N_404\ : std_logic;
signal \U712_CHIP_RAM.N_313_2\ : std_logic;
signal \U712_CHIP_RAM.N_312_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_314\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_37\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_396\ : std_logic;
signal \U712_CHIP_RAM.N_400\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lt7\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.N_231_cascade_\ : std_logic;
signal \A_c_14\ : std_logic;
signal \CLK40_PLL_i\ : std_logic;
signal \CLK40_PLL_i_i\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\ : std_logic;
signal \A_c_3\ : std_logic;
signal \A_c_10\ : std_logic;
signal \N_180_i\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1_cascade_\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_9\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \U712_BYTE_ENABLE.N_342\ : std_logic;
signal \U712_BYTE_ENABLE.N_341_cascade_\ : std_logic;
signal \N_55_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_320\ : std_logic;
signal \U712_BYTE_ENABLE.N_318_cascade_\ : std_logic;
signal \N_105_i\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \N_57_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_339\ : std_logic;
signal \U712_BYTE_ENABLE.N_206_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_316\ : std_logic;
signal \N_277_i\ : std_logic;
signal \LLBE_i_o2_i\ : std_logic;
signal \WEn_c\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \A_c_19\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\ : std_logic;
signal \A_c_13\ : std_logic;
signal \A_c_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z20\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A20C_net\ : std_logic;
signal \UMBEn_c\ : std_logic;
signal \A_c_1\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \N_276_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \RASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \CASn_c\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNIHMEAZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_0\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \un1_LDSn_i_0\ : std_logic;
signal \DS_ENm\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \N_87\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL_i\,
            REFERENCECLK => \N__3921\,
            RESETB => \N__7143\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11587\,
            DIN => \N__11586\,
            DOUT => \N__11585\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11587\,
            PADOUT => \N__11586\,
            PADIN => \N__11585\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7737\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11578\,
            DIN => \N__11577\,
            DOUT => \N__11576\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11578\,
            PADOUT => \N__11577\,
            PADIN => \N__11576\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11569\,
            DIN => \N__11568\,
            DOUT => \N__11567\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11569\,
            PADOUT => \N__11568\,
            PADIN => \N__11567\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9540\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11560\,
            DIN => \N__11559\,
            DOUT => \N__11558\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11560\,
            PADOUT => \N__11559\,
            PADIN => \N__11558\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6183\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11551\,
            DIN => \N__11550\,
            DOUT => \N__11549\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11551\,
            PADOUT => \N__11550\,
            PADIN => \N__11549\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11542\,
            DIN => \N__11541\,
            DOUT => \N__11540\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11542\,
            PADOUT => \N__11541\,
            PADIN => \N__11540\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11533\,
            DIN => \N__11532\,
            DOUT => \N__11531\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11533\,
            PADOUT => \N__11532\,
            PADIN => \N__11531\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11524\,
            DIN => \N__11523\,
            DOUT => \N__11522\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11524\,
            PADOUT => \N__11523\,
            PADIN => \N__11522\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11515\,
            DIN => \N__11514\,
            DOUT => \N__11513\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11515\,
            PADOUT => \N__11514\,
            PADIN => \N__11513\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11506\,
            DIN => \N__11505\,
            DOUT => \N__11504\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11506\,
            PADOUT => \N__11505\,
            PADIN => \N__11504\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11497\,
            DIN => \N__11496\,
            DOUT => \N__11495\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11497\,
            PADOUT => \N__11496\,
            PADIN => \N__11495\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9114\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11488\,
            DIN => \N__11487\,
            DOUT => \N__11486\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11488\,
            PADOUT => \N__11487\,
            PADIN => \N__11486\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8253\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11479\,
            DIN => \N__11478\,
            DOUT => \N__11477\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11479\,
            PADOUT => \N__11478\,
            PADIN => \N__11477\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11470\,
            DIN => \N__11469\,
            DOUT => \N__11468\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11470\,
            PADOUT => \N__11469\,
            PADIN => \N__11468\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4379\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11461\,
            DIN => \N__11460\,
            DOUT => \N__11459\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11461\,
            PADOUT => \N__11460\,
            PADIN => \N__11459\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11452\,
            DIN => \N__11451\,
            DOUT => \N__11450\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11452\,
            PADOUT => \N__11451\,
            PADIN => \N__11450\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11443\,
            DIN => \N__11442\,
            DOUT => \N__11441\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11443\,
            PADOUT => \N__11442\,
            PADIN => \N__11441\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4014\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11434\,
            DIN => \N__11433\,
            DOUT => \N__11432\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11434\,
            PADOUT => \N__11433\,
            PADIN => \N__11432\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11425\,
            DIN => \N__11424\,
            DOUT => \N__11423\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11425\,
            PADOUT => \N__11424\,
            PADIN => \N__11423\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11416\,
            DIN => \N__11415\,
            DOUT => \N__11414\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11416\,
            PADOUT => \N__11415\,
            PADIN => \N__11414\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8727\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11407\,
            DIN => \N__11406\,
            DOUT => \N__11405\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11407\,
            PADOUT => \N__11406\,
            PADIN => \N__11405\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11398\,
            DIN => \N__11397\,
            DOUT => \N__11396\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11398\,
            PADOUT => \N__11397\,
            PADIN => \N__11396\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8319\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11389\,
            DIN => \N__11388\,
            DOUT => \N__11387\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11389\,
            PADOUT => \N__11388\,
            PADIN => \N__11387\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11380\,
            DIN => \N__11379\,
            DOUT => \N__11378\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11380\,
            PADOUT => \N__11379\,
            PADIN => \N__11378\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8241\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11371\,
            DIN => \N__11370\,
            DOUT => \N__11369\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11371\,
            PADOUT => \N__11370\,
            PADIN => \N__11369\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11362\,
            DIN => \N__11361\,
            DOUT => \N__11360\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11362\,
            PADOUT => \N__11361\,
            PADIN => \N__11360\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11353\,
            DIN => \N__11352\,
            DOUT => \N__11351\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11353\,
            PADOUT => \N__11352\,
            PADIN => \N__11351\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11344\,
            DIN => \N__11343\,
            DOUT => \N__11342\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11344\,
            PADOUT => \N__11343\,
            PADIN => \N__11342\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11335\,
            DIN => \N__11334\,
            DOUT => \N__11333\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11335\,
            PADOUT => \N__11334\,
            PADIN => \N__11333\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11326\,
            DIN => \N__11325\,
            DOUT => \N__11324\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11326\,
            PADOUT => \N__11325\,
            PADIN => \N__11324\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4026\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11317\,
            DIN => \N__11316\,
            DOUT => \N__11315\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11317\,
            PADOUT => \N__11316\,
            PADIN => \N__11315\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11308\,
            DIN => \N__11307\,
            DOUT => \N__11306\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11308\,
            PADOUT => \N__11307\,
            PADIN => \N__11306\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11299\,
            DIN => \N__11298\,
            DOUT => \N__11297\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11299\,
            PADOUT => \N__11298\,
            PADIN => \N__11297\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11290\,
            DIN => \N__11289\,
            DOUT => \N__11288\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11290\,
            PADOUT => \N__11289\,
            PADIN => \N__11288\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11281\,
            DIN => \N__11280\,
            DOUT => \N__11279\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11281\,
            PADOUT => \N__11280\,
            PADIN => \N__11279\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11272\,
            DIN => \N__11271\,
            DOUT => \N__11270\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11272\,
            PADOUT => \N__11271\,
            PADIN => \N__11270\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5088\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11263\,
            DIN => \N__11262\,
            DOUT => \N__11261\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11263\,
            PADOUT => \N__11262\,
            PADIN => \N__11261\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9900\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11254\,
            DIN => \N__11253\,
            DOUT => \N__11252\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11254\,
            PADOUT => \N__11253\,
            PADIN => \N__11252\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7029\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11245\,
            DIN => \N__11244\,
            DOUT => \N__11243\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11245\,
            PADOUT => \N__11244\,
            PADIN => \N__11243\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11236\,
            DIN => \N__11235\,
            DOUT => \N__11234\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11236\,
            PADOUT => \N__11235\,
            PADIN => \N__11234\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8379\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11227\,
            DIN => \N__11226\,
            DOUT => \N__11225\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11227\,
            PADOUT => \N__11226\,
            PADIN => \N__11225\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11218\,
            DIN => \N__11217\,
            DOUT => \N__11216\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11218\,
            PADOUT => \N__11217\,
            PADIN => \N__11216\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4461\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11209\,
            DIN => \N__11208\,
            DOUT => \N__11207\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11209\,
            PADOUT => \N__11208\,
            PADIN => \N__11207\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7025\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11200\,
            DIN => \N__11199\,
            DOUT => \N__11198\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11200\,
            PADOUT => \N__11199\,
            PADIN => \N__11198\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3999\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11191\,
            DIN => \N__11190\,
            DOUT => \N__11189\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11191\,
            PADOUT => \N__11190\,
            PADIN => \N__11189\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11182\,
            DIN => \N__11181\,
            DOUT => \N__11180\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11182\,
            PADOUT => \N__11181\,
            PADIN => \N__11180\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6342\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11173\,
            DIN => \N__11172\,
            DOUT => \N__11171\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11173\,
            PADOUT => \N__11172\,
            PADIN => \N__11171\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7236\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11164\,
            DIN => \N__11163\,
            DOUT => \N__11162\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11164\,
            PADOUT => \N__11163\,
            PADIN => \N__11162\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11155\,
            DIN => \N__11154\,
            DOUT => \N__11153\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11155\,
            PADOUT => \N__11154\,
            PADIN => \N__11153\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11146\,
            DIN => \N__11145\,
            DOUT => \N__11144\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11146\,
            PADOUT => \N__11145\,
            PADIN => \N__11144\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11137\,
            DIN => \N__11136\,
            DOUT => \N__11135\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11137\,
            PADOUT => \N__11136\,
            PADIN => \N__11135\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11128\,
            DIN => \N__11127\,
            DOUT => \N__11126\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11128\,
            PADOUT => \N__11127\,
            PADIN => \N__11126\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8031\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11119\,
            DIN => \N__11118\,
            DOUT => \N__11117\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11119\,
            PADOUT => \N__11118\,
            PADIN => \N__11117\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11110\,
            DIN => \N__11109\,
            DOUT => \N__11108\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11110\,
            PADOUT => \N__11109\,
            PADIN => \N__11108\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7018\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11101\,
            DIN => \N__11100\,
            DOUT => \N__11099\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11101\,
            PADOUT => \N__11100\,
            PADIN => \N__11099\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9135\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11092\,
            DIN => \N__11091\,
            DOUT => \N__11090\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11092\,
            PADOUT => \N__11091\,
            PADIN => \N__11090\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4380\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11083\,
            DIN => \N__11082\,
            DOUT => \N__11081\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11083\,
            PADOUT => \N__11082\,
            PADIN => \N__11081\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7467\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11074\,
            DIN => \N__11073\,
            DOUT => \N__11072\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11074\,
            PADOUT => \N__11073\,
            PADIN => \N__11072\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8124\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11065\,
            DIN => \N__11064\,
            DOUT => \N__11063\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11065\,
            PADOUT => \N__11064\,
            PADIN => \N__11063\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6338\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11056\,
            DIN => \N__11055\,
            DOUT => \N__11054\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11056\,
            PADOUT => \N__11055\,
            PADIN => \N__11054\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11047\,
            DIN => \N__11046\,
            DOUT => \N__11045\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11047\,
            PADOUT => \N__11046\,
            PADIN => \N__11045\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11038\,
            DIN => \N__11037\,
            DOUT => \N__11036\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11038\,
            PADOUT => \N__11037\,
            PADIN => \N__11036\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7680\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11029\,
            DIN => \N__11028\,
            DOUT => \N__11027\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11029\,
            PADOUT => \N__11028\,
            PADIN => \N__11027\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8226\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11020\,
            DIN => \N__11019\,
            DOUT => \N__11018\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11020\,
            PADOUT => \N__11019\,
            PADIN => \N__11018\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4182\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11011\,
            DIN => \N__11010\,
            DOUT => \N__11009\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11011\,
            PADOUT => \N__11010\,
            PADIN => \N__11009\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8001\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11002\,
            DIN => \N__11001\,
            DOUT => \N__11000\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11002\,
            PADOUT => \N__11001\,
            PADIN => \N__11000\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10993\,
            DIN => \N__10992\,
            DOUT => \N__10991\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10993\,
            PADOUT => \N__10992\,
            PADIN => \N__10991\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10984\,
            DIN => \N__10983\,
            DOUT => \N__10982\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10984\,
            PADOUT => \N__10983\,
            PADIN => \N__10982\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10975\,
            DIN => \N__10974\,
            DOUT => \N__10973\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10975\,
            PADOUT => \N__10974\,
            PADIN => \N__10973\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10966\,
            DIN => \N__10965\,
            DOUT => \N__10964\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10966\,
            PADOUT => \N__10965\,
            PADIN => \N__10964\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7212\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10957\,
            DIN => \N__10956\,
            DOUT => \N__10955\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10957\,
            PADOUT => \N__10956\,
            PADIN => \N__10955\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8457\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10948\,
            DIN => \N__10947\,
            DOUT => \N__10946\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10948\,
            PADOUT => \N__10947\,
            PADIN => \N__10946\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10939\,
            DIN => \N__10938\,
            DOUT => \N__10937\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10939\,
            PADOUT => \N__10938\,
            PADIN => \N__10937\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7398\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10930\,
            DIN => \N__10929\,
            DOUT => \N__10928\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__10930\,
            PADOUT => \N__10929\,
            PADIN => \N__10928\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4044\,
            DIN0 => OPEN,
            DOUT0 => \N__6567\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10921\,
            DIN => \N__10920\,
            DOUT => \N__10919\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10921\,
            PADOUT => \N__10920\,
            PADIN => \N__10919\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7977\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10912\,
            DIN => \N__10911\,
            DOUT => \N__10910\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10912\,
            PADOUT => \N__10911\,
            PADIN => \N__10910\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10903\,
            DIN => \N__10902\,
            DOUT => \N__10901\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10903\,
            PADOUT => \N__10902\,
            PADIN => \N__10901\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10894\,
            DIN => \N__10893\,
            DOUT => \N__10892\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10894\,
            PADOUT => \N__10893\,
            PADIN => \N__10892\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8187\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10885\,
            DIN => \N__10884\,
            DOUT => \N__10883\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10885\,
            PADOUT => \N__10884\,
            PADIN => \N__10883\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10876\,
            DIN => \N__10875\,
            DOUT => \N__10874\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10876\,
            PADOUT => \N__10875\,
            PADIN => \N__10874\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10867\,
            DIN => \N__10866\,
            DOUT => \N__10865\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10867\,
            PADOUT => \N__10866\,
            PADIN => \N__10865\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10858\,
            DIN => \N__10857\,
            DOUT => \N__10856\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10858\,
            PADOUT => \N__10857\,
            PADIN => \N__10856\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10849\,
            DIN => \N__10848\,
            DOUT => \N__10847\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10849\,
            PADOUT => \N__10848\,
            PADIN => \N__10847\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7632\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10840\,
            DIN => \N__10839\,
            DOUT => \N__10838\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10840\,
            PADOUT => \N__10839\,
            PADIN => \N__10838\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9660\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10831\,
            DIN => \N__10830\,
            DOUT => \N__10829\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10831\,
            PADOUT => \N__10830\,
            PADIN => \N__10829\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8610\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10822\,
            DIN => \N__10821\,
            DOUT => \N__10820\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10822\,
            PADOUT => \N__10821\,
            PADIN => \N__10820\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6093\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10813\,
            DIN => \N__10812\,
            DOUT => \N__10811\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10813\,
            PADOUT => \N__10812\,
            PADIN => \N__10811\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10804\,
            DIN => \N__10803\,
            DOUT => \N__10802\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10804\,
            PADOUT => \N__10803\,
            PADIN => \N__10802\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10795\,
            DIN => \N__10794\,
            DOUT => \N__10793\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10795\,
            PADOUT => \N__10794\,
            PADIN => \N__10793\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8988\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10786\,
            DIN => \N__10785\,
            DOUT => \N__10784\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10786\,
            PADOUT => \N__10785\,
            PADIN => \N__10784\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2625\ : InMux
    port map (
            O => \N__10767\,
            I => \N__10763\
        );

    \I__2624\ : CascadeMux
    port map (
            O => \N__10766\,
            I => \N__10760\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__10763\,
            I => \N__10757\
        );

    \I__2622\ : InMux
    port map (
            O => \N__10760\,
            I => \N__10754\
        );

    \I__2621\ : Span4Mux_h
    port map (
            O => \N__10757\,
            I => \N__10748\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__10754\,
            I => \N__10748\
        );

    \I__2619\ : InMux
    port map (
            O => \N__10753\,
            I => \N__10745\
        );

    \I__2618\ : Span4Mux_v
    port map (
            O => \N__10748\,
            I => \N__10741\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__10745\,
            I => \N__10738\
        );

    \I__2616\ : InMux
    port map (
            O => \N__10744\,
            I => \N__10735\
        );

    \I__2615\ : Sp12to4
    port map (
            O => \N__10741\,
            I => \N__10732\
        );

    \I__2614\ : Sp12to4
    port map (
            O => \N__10738\,
            I => \N__10727\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__10735\,
            I => \N__10727\
        );

    \I__2612\ : Span12Mux_h
    port map (
            O => \N__10732\,
            I => \N__10724\
        );

    \I__2611\ : Span12Mux_v
    port map (
            O => \N__10727\,
            I => \N__10721\
        );

    \I__2610\ : Span12Mux_v
    port map (
            O => \N__10724\,
            I => \N__10718\
        );

    \I__2609\ : Span12Mux_v
    port map (
            O => \N__10721\,
            I => \N__10715\
        );

    \I__2608\ : Odrv12
    port map (
            O => \N__10718\,
            I => \DRA_c_9\
        );

    \I__2607\ : Odrv12
    port map (
            O => \N__10715\,
            I => \DRA_c_9\
        );

    \I__2606\ : InMux
    port map (
            O => \N__10710\,
            I => \N__10704\
        );

    \I__2605\ : CascadeMux
    port map (
            O => \N__10709\,
            I => \N__10699\
        );

    \I__2604\ : CascadeMux
    port map (
            O => \N__10708\,
            I => \N__10689\
        );

    \I__2603\ : CascadeMux
    port map (
            O => \N__10707\,
            I => \N__10685\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__10704\,
            I => \N__10681\
        );

    \I__2601\ : InMux
    port map (
            O => \N__10703\,
            I => \N__10676\
        );

    \I__2600\ : InMux
    port map (
            O => \N__10702\,
            I => \N__10665\
        );

    \I__2599\ : InMux
    port map (
            O => \N__10699\,
            I => \N__10665\
        );

    \I__2598\ : InMux
    port map (
            O => \N__10698\,
            I => \N__10665\
        );

    \I__2597\ : InMux
    port map (
            O => \N__10697\,
            I => \N__10665\
        );

    \I__2596\ : InMux
    port map (
            O => \N__10696\,
            I => \N__10665\
        );

    \I__2595\ : CascadeMux
    port map (
            O => \N__10695\,
            I => \N__10662\
        );

    \I__2594\ : CascadeMux
    port map (
            O => \N__10694\,
            I => \N__10657\
        );

    \I__2593\ : CascadeMux
    port map (
            O => \N__10693\,
            I => \N__10654\
        );

    \I__2592\ : InMux
    port map (
            O => \N__10692\,
            I => \N__10646\
        );

    \I__2591\ : InMux
    port map (
            O => \N__10689\,
            I => \N__10646\
        );

    \I__2590\ : InMux
    port map (
            O => \N__10688\,
            I => \N__10646\
        );

    \I__2589\ : InMux
    port map (
            O => \N__10685\,
            I => \N__10641\
        );

    \I__2588\ : InMux
    port map (
            O => \N__10684\,
            I => \N__10641\
        );

    \I__2587\ : Span4Mux_v
    port map (
            O => \N__10681\,
            I => \N__10638\
        );

    \I__2586\ : InMux
    port map (
            O => \N__10680\,
            I => \N__10635\
        );

    \I__2585\ : InMux
    port map (
            O => \N__10679\,
            I => \N__10632\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__10676\,
            I => \N__10627\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__10665\,
            I => \N__10627\
        );

    \I__2582\ : InMux
    port map (
            O => \N__10662\,
            I => \N__10622\
        );

    \I__2581\ : InMux
    port map (
            O => \N__10661\,
            I => \N__10622\
        );

    \I__2580\ : InMux
    port map (
            O => \N__10660\,
            I => \N__10612\
        );

    \I__2579\ : InMux
    port map (
            O => \N__10657\,
            I => \N__10612\
        );

    \I__2578\ : InMux
    port map (
            O => \N__10654\,
            I => \N__10612\
        );

    \I__2577\ : InMux
    port map (
            O => \N__10653\,
            I => \N__10612\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__10646\,
            I => \N__10607\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__10641\,
            I => \N__10607\
        );

    \I__2574\ : Span4Mux_h
    port map (
            O => \N__10638\,
            I => \N__10596\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__10635\,
            I => \N__10596\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__10632\,
            I => \N__10596\
        );

    \I__2571\ : Span4Mux_v
    port map (
            O => \N__10627\,
            I => \N__10596\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__10622\,
            I => \N__10596\
        );

    \I__2569\ : InMux
    port map (
            O => \N__10621\,
            I => \N__10593\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__10612\,
            I => \N__10590\
        );

    \I__2567\ : Span4Mux_v
    port map (
            O => \N__10607\,
            I => \N__10583\
        );

    \I__2566\ : Span4Mux_h
    port map (
            O => \N__10596\,
            I => \N__10583\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__10593\,
            I => \N__10583\
        );

    \I__2564\ : Span4Mux_v
    port map (
            O => \N__10590\,
            I => \N__10580\
        );

    \I__2563\ : Span4Mux_h
    port map (
            O => \N__10583\,
            I => \N__10577\
        );

    \I__2562\ : Span4Mux_v
    port map (
            O => \N__10580\,
            I => \N__10574\
        );

    \I__2561\ : Span4Mux_h
    port map (
            O => \N__10577\,
            I => \N__10571\
        );

    \I__2560\ : Sp12to4
    port map (
            O => \N__10574\,
            I => \N__10568\
        );

    \I__2559\ : Sp12to4
    port map (
            O => \N__10571\,
            I => \N__10565\
        );

    \I__2558\ : Span12Mux_h
    port map (
            O => \N__10568\,
            I => \N__10562\
        );

    \I__2557\ : Span12Mux_v
    port map (
            O => \N__10565\,
            I => \N__10559\
        );

    \I__2556\ : Odrv12
    port map (
            O => \N__10562\,
            I => \AGNUS_REV_c\
        );

    \I__2555\ : Odrv12
    port map (
            O => \N__10559\,
            I => \AGNUS_REV_c\
        );

    \I__2554\ : InMux
    port map (
            O => \N__10554\,
            I => \N__10550\
        );

    \I__2553\ : InMux
    port map (
            O => \N__10553\,
            I => \N__10547\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__10550\,
            I => \N__10541\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__10547\,
            I => \N__10541\
        );

    \I__2550\ : InMux
    port map (
            O => \N__10546\,
            I => \N__10538\
        );

    \I__2549\ : Span4Mux_v
    port map (
            O => \N__10541\,
            I => \N__10532\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__10538\,
            I => \N__10532\
        );

    \I__2547\ : InMux
    port map (
            O => \N__10537\,
            I => \N__10529\
        );

    \I__2546\ : Sp12to4
    port map (
            O => \N__10532\,
            I => \N__10524\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__10529\,
            I => \N__10524\
        );

    \I__2544\ : Odrv12
    port map (
            O => \N__10524\,
            I => \DRA_c_8\
        );

    \I__2543\ : InMux
    port map (
            O => \N__10521\,
            I => \N__10518\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__10518\,
            I => \N__10515\
        );

    \I__2541\ : Span4Mux_h
    port map (
            O => \N__10515\,
            I => \N__10512\
        );

    \I__2540\ : Odrv4
    port map (
            O => \N__10512\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__2539\ : CEMux
    port map (
            O => \N__10509\,
            I => \N__10485\
        );

    \I__2538\ : CEMux
    port map (
            O => \N__10508\,
            I => \N__10485\
        );

    \I__2537\ : CEMux
    port map (
            O => \N__10507\,
            I => \N__10485\
        );

    \I__2536\ : CEMux
    port map (
            O => \N__10506\,
            I => \N__10485\
        );

    \I__2535\ : CEMux
    port map (
            O => \N__10505\,
            I => \N__10485\
        );

    \I__2534\ : CEMux
    port map (
            O => \N__10504\,
            I => \N__10485\
        );

    \I__2533\ : CEMux
    port map (
            O => \N__10503\,
            I => \N__10485\
        );

    \I__2532\ : CEMux
    port map (
            O => \N__10502\,
            I => \N__10485\
        );

    \I__2531\ : GlobalMux
    port map (
            O => \N__10485\,
            I => \N__10482\
        );

    \I__2530\ : gio2CtrlBuf
    port map (
            O => \N__10482\,
            I => \DBRn_c_i_0_g\
        );

    \I__2529\ : InMux
    port map (
            O => \N__10479\,
            I => \N__10470\
        );

    \I__2528\ : InMux
    port map (
            O => \N__10478\,
            I => \N__10465\
        );

    \I__2527\ : InMux
    port map (
            O => \N__10477\,
            I => \N__10465\
        );

    \I__2526\ : InMux
    port map (
            O => \N__10476\,
            I => \N__10462\
        );

    \I__2525\ : InMux
    port map (
            O => \N__10475\,
            I => \N__10459\
        );

    \I__2524\ : InMux
    port map (
            O => \N__10474\,
            I => \N__10456\
        );

    \I__2523\ : InMux
    port map (
            O => \N__10473\,
            I => \N__10453\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__10470\,
            I => \N__10448\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__10465\,
            I => \N__10439\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__10462\,
            I => \N__10431\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__10459\,
            I => \N__10417\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__10456\,
            I => \N__10406\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__10453\,
            I => \N__10395\
        );

    \I__2516\ : SRMux
    port map (
            O => \N__10452\,
            I => \N__10299\
        );

    \I__2515\ : SRMux
    port map (
            O => \N__10451\,
            I => \N__10299\
        );

    \I__2514\ : Glb2LocalMux
    port map (
            O => \N__10448\,
            I => \N__10299\
        );

    \I__2513\ : SRMux
    port map (
            O => \N__10447\,
            I => \N__10299\
        );

    \I__2512\ : SRMux
    port map (
            O => \N__10446\,
            I => \N__10299\
        );

    \I__2511\ : SRMux
    port map (
            O => \N__10445\,
            I => \N__10299\
        );

    \I__2510\ : SRMux
    port map (
            O => \N__10444\,
            I => \N__10299\
        );

    \I__2509\ : SRMux
    port map (
            O => \N__10443\,
            I => \N__10299\
        );

    \I__2508\ : SRMux
    port map (
            O => \N__10442\,
            I => \N__10299\
        );

    \I__2507\ : Glb2LocalMux
    port map (
            O => \N__10439\,
            I => \N__10299\
        );

    \I__2506\ : SRMux
    port map (
            O => \N__10438\,
            I => \N__10299\
        );

    \I__2505\ : SRMux
    port map (
            O => \N__10437\,
            I => \N__10299\
        );

    \I__2504\ : SRMux
    port map (
            O => \N__10436\,
            I => \N__10299\
        );

    \I__2503\ : SRMux
    port map (
            O => \N__10435\,
            I => \N__10299\
        );

    \I__2502\ : SRMux
    port map (
            O => \N__10434\,
            I => \N__10299\
        );

    \I__2501\ : Glb2LocalMux
    port map (
            O => \N__10431\,
            I => \N__10299\
        );

    \I__2500\ : SRMux
    port map (
            O => \N__10430\,
            I => \N__10299\
        );

    \I__2499\ : SRMux
    port map (
            O => \N__10429\,
            I => \N__10299\
        );

    \I__2498\ : SRMux
    port map (
            O => \N__10428\,
            I => \N__10299\
        );

    \I__2497\ : SRMux
    port map (
            O => \N__10427\,
            I => \N__10299\
        );

    \I__2496\ : SRMux
    port map (
            O => \N__10426\,
            I => \N__10299\
        );

    \I__2495\ : SRMux
    port map (
            O => \N__10425\,
            I => \N__10299\
        );

    \I__2494\ : SRMux
    port map (
            O => \N__10424\,
            I => \N__10299\
        );

    \I__2493\ : SRMux
    port map (
            O => \N__10423\,
            I => \N__10299\
        );

    \I__2492\ : SRMux
    port map (
            O => \N__10422\,
            I => \N__10299\
        );

    \I__2491\ : SRMux
    port map (
            O => \N__10421\,
            I => \N__10299\
        );

    \I__2490\ : SRMux
    port map (
            O => \N__10420\,
            I => \N__10299\
        );

    \I__2489\ : Glb2LocalMux
    port map (
            O => \N__10417\,
            I => \N__10299\
        );

    \I__2488\ : SRMux
    port map (
            O => \N__10416\,
            I => \N__10299\
        );

    \I__2487\ : SRMux
    port map (
            O => \N__10415\,
            I => \N__10299\
        );

    \I__2486\ : SRMux
    port map (
            O => \N__10414\,
            I => \N__10299\
        );

    \I__2485\ : SRMux
    port map (
            O => \N__10413\,
            I => \N__10299\
        );

    \I__2484\ : SRMux
    port map (
            O => \N__10412\,
            I => \N__10299\
        );

    \I__2483\ : SRMux
    port map (
            O => \N__10411\,
            I => \N__10299\
        );

    \I__2482\ : SRMux
    port map (
            O => \N__10410\,
            I => \N__10299\
        );

    \I__2481\ : SRMux
    port map (
            O => \N__10409\,
            I => \N__10299\
        );

    \I__2480\ : Glb2LocalMux
    port map (
            O => \N__10406\,
            I => \N__10299\
        );

    \I__2479\ : SRMux
    port map (
            O => \N__10405\,
            I => \N__10299\
        );

    \I__2478\ : SRMux
    port map (
            O => \N__10404\,
            I => \N__10299\
        );

    \I__2477\ : SRMux
    port map (
            O => \N__10403\,
            I => \N__10299\
        );

    \I__2476\ : SRMux
    port map (
            O => \N__10402\,
            I => \N__10299\
        );

    \I__2475\ : SRMux
    port map (
            O => \N__10401\,
            I => \N__10299\
        );

    \I__2474\ : SRMux
    port map (
            O => \N__10400\,
            I => \N__10299\
        );

    \I__2473\ : SRMux
    port map (
            O => \N__10399\,
            I => \N__10299\
        );

    \I__2472\ : SRMux
    port map (
            O => \N__10398\,
            I => \N__10299\
        );

    \I__2471\ : Glb2LocalMux
    port map (
            O => \N__10395\,
            I => \N__10299\
        );

    \I__2470\ : SRMux
    port map (
            O => \N__10394\,
            I => \N__10299\
        );

    \I__2469\ : GlobalMux
    port map (
            O => \N__10299\,
            I => \N__10296\
        );

    \I__2468\ : gio2CtrlBuf
    port map (
            O => \N__10296\,
            I => \RESETn_c_i_g\
        );

    \I__2467\ : InMux
    port map (
            O => \N__10293\,
            I => \N__10290\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__10290\,
            I => \N__10287\
        );

    \I__2465\ : Odrv12
    port map (
            O => \N__10287\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__2464\ : InMux
    port map (
            O => \N__10284\,
            I => \N__10278\
        );

    \I__2463\ : InMux
    port map (
            O => \N__10283\,
            I => \N__10278\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__10278\,
            I => \N__10273\
        );

    \I__2461\ : InMux
    port map (
            O => \N__10277\,
            I => \N__10268\
        );

    \I__2460\ : InMux
    port map (
            O => \N__10276\,
            I => \N__10268\
        );

    \I__2459\ : Span4Mux_h
    port map (
            O => \N__10273\,
            I => \N__10263\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__10268\,
            I => \N__10263\
        );

    \I__2457\ : Sp12to4
    port map (
            O => \N__10263\,
            I => \N__10260\
        );

    \I__2456\ : Span12Mux_v
    port map (
            O => \N__10260\,
            I => \N__10257\
        );

    \I__2455\ : Odrv12
    port map (
            O => \N__10257\,
            I => \DRA_c_3\
        );

    \I__2454\ : InMux
    port map (
            O => \N__10254\,
            I => \N__10251\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__10251\,
            I => \N__10248\
        );

    \I__2452\ : Odrv4
    port map (
            O => \N__10248\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__2451\ : InMux
    port map (
            O => \N__10245\,
            I => \N__10239\
        );

    \I__2450\ : InMux
    port map (
            O => \N__10244\,
            I => \N__10239\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__10239\,
            I => \N__10236\
        );

    \I__2448\ : Span4Mux_v
    port map (
            O => \N__10236\,
            I => \N__10231\
        );

    \I__2447\ : InMux
    port map (
            O => \N__10235\,
            I => \N__10228\
        );

    \I__2446\ : InMux
    port map (
            O => \N__10234\,
            I => \N__10225\
        );

    \I__2445\ : Sp12to4
    port map (
            O => \N__10231\,
            I => \N__10220\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__10228\,
            I => \N__10220\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__10225\,
            I => \N__10217\
        );

    \I__2442\ : Span12Mux_h
    port map (
            O => \N__10220\,
            I => \N__10214\
        );

    \I__2441\ : Sp12to4
    port map (
            O => \N__10217\,
            I => \N__10211\
        );

    \I__2440\ : Span12Mux_v
    port map (
            O => \N__10214\,
            I => \N__10208\
        );

    \I__2439\ : Span12Mux_v
    port map (
            O => \N__10211\,
            I => \N__10205\
        );

    \I__2438\ : Odrv12
    port map (
            O => \N__10208\,
            I => \DRA_c_1\
        );

    \I__2437\ : Odrv12
    port map (
            O => \N__10205\,
            I => \DRA_c_1\
        );

    \I__2436\ : InMux
    port map (
            O => \N__10200\,
            I => \N__10196\
        );

    \I__2435\ : InMux
    port map (
            O => \N__10199\,
            I => \N__10193\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__10196\,
            I => \N__10188\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__10193\,
            I => \N__10188\
        );

    \I__2432\ : Span4Mux_h
    port map (
            O => \N__10188\,
            I => \N__10185\
        );

    \I__2431\ : Sp12to4
    port map (
            O => \N__10185\,
            I => \N__10182\
        );

    \I__2430\ : Span12Mux_v
    port map (
            O => \N__10182\,
            I => \N__10179\
        );

    \I__2429\ : Odrv12
    port map (
            O => \N__10179\,
            I => \DRA_c_0\
        );

    \I__2428\ : InMux
    port map (
            O => \N__10176\,
            I => \N__10173\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__10173\,
            I => \N__10170\
        );

    \I__2426\ : Span4Mux_v
    port map (
            O => \N__10170\,
            I => \N__10167\
        );

    \I__2425\ : Sp12to4
    port map (
            O => \N__10167\,
            I => \N__10164\
        );

    \I__2424\ : Odrv12
    port map (
            O => \N__10164\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__2423\ : InMux
    port map (
            O => \N__10161\,
            I => \N__10158\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__10158\,
            I => \N__10155\
        );

    \I__2421\ : Span4Mux_h
    port map (
            O => \N__10155\,
            I => \N__10152\
        );

    \I__2420\ : Span4Mux_h
    port map (
            O => \N__10152\,
            I => \N__10149\
        );

    \I__2419\ : Odrv4
    port map (
            O => \N__10149\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__2418\ : InMux
    port map (
            O => \N__10146\,
            I => \N__10143\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__10143\,
            I => \N__10140\
        );

    \I__2416\ : Span4Mux_v
    port map (
            O => \N__10140\,
            I => \N__10137\
        );

    \I__2415\ : Odrv4
    port map (
            O => \N__10137\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__2414\ : InMux
    port map (
            O => \N__10134\,
            I => \N__10128\
        );

    \I__2413\ : InMux
    port map (
            O => \N__10133\,
            I => \N__10125\
        );

    \I__2412\ : InMux
    port map (
            O => \N__10132\,
            I => \N__10122\
        );

    \I__2411\ : InMux
    port map (
            O => \N__10131\,
            I => \N__10119\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__10128\,
            I => \N__10110\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__10125\,
            I => \N__10110\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__10122\,
            I => \N__10110\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__10119\,
            I => \N__10110\
        );

    \I__2406\ : Span4Mux_v
    port map (
            O => \N__10110\,
            I => \N__10107\
        );

    \I__2405\ : Sp12to4
    port map (
            O => \N__10107\,
            I => \N__10104\
        );

    \I__2404\ : Span12Mux_h
    port map (
            O => \N__10104\,
            I => \N__10101\
        );

    \I__2403\ : Odrv12
    port map (
            O => \N__10101\,
            I => \DRA_c_7\
        );

    \I__2402\ : InMux
    port map (
            O => \N__10098\,
            I => \N__10095\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__10095\,
            I => \N__10092\
        );

    \I__2400\ : Span4Mux_h
    port map (
            O => \N__10092\,
            I => \N__10089\
        );

    \I__2399\ : Odrv4
    port map (
            O => \N__10089\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__2398\ : InMux
    port map (
            O => \N__10086\,
            I => \N__10079\
        );

    \I__2397\ : InMux
    port map (
            O => \N__10085\,
            I => \N__10079\
        );

    \I__2396\ : InMux
    port map (
            O => \N__10084\,
            I => \N__10076\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__10079\,
            I => \N__10072\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__10076\,
            I => \N__10069\
        );

    \I__2393\ : InMux
    port map (
            O => \N__10075\,
            I => \N__10066\
        );

    \I__2392\ : Span4Mux_v
    port map (
            O => \N__10072\,
            I => \N__10063\
        );

    \I__2391\ : Span4Mux_h
    port map (
            O => \N__10069\,
            I => \N__10058\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__10066\,
            I => \N__10058\
        );

    \I__2389\ : Span4Mux_v
    port map (
            O => \N__10063\,
            I => \N__10055\
        );

    \I__2388\ : Span4Mux_v
    port map (
            O => \N__10058\,
            I => \N__10052\
        );

    \I__2387\ : Span4Mux_h
    port map (
            O => \N__10055\,
            I => \N__10049\
        );

    \I__2386\ : Span4Mux_v
    port map (
            O => \N__10052\,
            I => \N__10046\
        );

    \I__2385\ : Sp12to4
    port map (
            O => \N__10049\,
            I => \N__10041\
        );

    \I__2384\ : Sp12to4
    port map (
            O => \N__10046\,
            I => \N__10041\
        );

    \I__2383\ : Odrv12
    port map (
            O => \N__10041\,
            I => \DRA_c_4\
        );

    \I__2382\ : InMux
    port map (
            O => \N__10038\,
            I => \N__10035\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__10035\,
            I => \N__10032\
        );

    \I__2380\ : Span4Mux_v
    port map (
            O => \N__10032\,
            I => \N__10029\
        );

    \I__2379\ : Odrv4
    port map (
            O => \N__10029\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2378\ : InMux
    port map (
            O => \N__10026\,
            I => \N__10023\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__10023\,
            I => \N__10017\
        );

    \I__2376\ : InMux
    port map (
            O => \N__10022\,
            I => \N__10014\
        );

    \I__2375\ : InMux
    port map (
            O => \N__10021\,
            I => \N__10011\
        );

    \I__2374\ : InMux
    port map (
            O => \N__10020\,
            I => \N__10008\
        );

    \I__2373\ : Span4Mux_v
    port map (
            O => \N__10017\,
            I => \N__10005\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__10014\,
            I => \N__9998\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__10011\,
            I => \N__9998\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__10008\,
            I => \N__9998\
        );

    \I__2369\ : Span4Mux_v
    port map (
            O => \N__10005\,
            I => \N__9995\
        );

    \I__2368\ : Sp12to4
    port map (
            O => \N__9998\,
            I => \N__9992\
        );

    \I__2367\ : Sp12to4
    port map (
            O => \N__9995\,
            I => \N__9987\
        );

    \I__2366\ : Span12Mux_v
    port map (
            O => \N__9992\,
            I => \N__9987\
        );

    \I__2365\ : Odrv12
    port map (
            O => \N__9987\,
            I => \DRA_c_6\
        );

    \I__2364\ : InMux
    port map (
            O => \N__9984\,
            I => \N__9981\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__9981\,
            I => \N__9975\
        );

    \I__2362\ : InMux
    port map (
            O => \N__9980\,
            I => \N__9972\
        );

    \I__2361\ : InMux
    port map (
            O => \N__9979\,
            I => \N__9967\
        );

    \I__2360\ : InMux
    port map (
            O => \N__9978\,
            I => \N__9967\
        );

    \I__2359\ : Span4Mux_h
    port map (
            O => \N__9975\,
            I => \N__9962\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__9972\,
            I => \N__9962\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__9967\,
            I => \N__9957\
        );

    \I__2356\ : Sp12to4
    port map (
            O => \N__9962\,
            I => \N__9957\
        );

    \I__2355\ : Span12Mux_v
    port map (
            O => \N__9957\,
            I => \N__9954\
        );

    \I__2354\ : Odrv12
    port map (
            O => \N__9954\,
            I => \DRA_c_5\
        );

    \I__2353\ : InMux
    port map (
            O => \N__9951\,
            I => \N__9945\
        );

    \I__2352\ : InMux
    port map (
            O => \N__9950\,
            I => \N__9945\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__9945\,
            I => \N__9942\
        );

    \I__2350\ : Span12Mux_v
    port map (
            O => \N__9942\,
            I => \N__9939\
        );

    \I__2349\ : Odrv12
    port map (
            O => \N__9939\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__2348\ : ClkMux
    port map (
            O => \N__9936\,
            I => \N__9924\
        );

    \I__2347\ : ClkMux
    port map (
            O => \N__9935\,
            I => \N__9924\
        );

    \I__2346\ : ClkMux
    port map (
            O => \N__9934\,
            I => \N__9924\
        );

    \I__2345\ : ClkMux
    port map (
            O => \N__9933\,
            I => \N__9924\
        );

    \I__2344\ : GlobalMux
    port map (
            O => \N__9924\,
            I => \N__9921\
        );

    \I__2343\ : gio2CtrlBuf
    port map (
            O => \N__9921\,
            I => \C3_c_g\
        );

    \I__2342\ : InMux
    port map (
            O => \N__9918\,
            I => \N__9915\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__9915\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2340\ : InMux
    port map (
            O => \N__9912\,
            I => \N__9909\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__9909\,
            I => \N__9906\
        );

    \I__2338\ : Span4Mux_h
    port map (
            O => \N__9906\,
            I => \N__9903\
        );

    \I__2337\ : Odrv4
    port map (
            O => \N__9903\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__2336\ : IoInMux
    port map (
            O => \N__9900\,
            I => \N__9897\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__9897\,
            I => \N__9894\
        );

    \I__2334\ : Span4Mux_s3_v
    port map (
            O => \N__9894\,
            I => \N__9891\
        );

    \I__2333\ : Span4Mux_h
    port map (
            O => \N__9891\,
            I => \N__9888\
        );

    \I__2332\ : Span4Mux_v
    port map (
            O => \N__9888\,
            I => \N__9885\
        );

    \I__2331\ : Odrv4
    port map (
            O => \N__9885\,
            I => \un1_LDSn_i_0\
        );

    \I__2330\ : InMux
    port map (
            O => \N__9882\,
            I => \N__9878\
        );

    \I__2329\ : InMux
    port map (
            O => \N__9881\,
            I => \N__9875\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__9878\,
            I => \N__9870\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__9875\,
            I => \N__9870\
        );

    \I__2326\ : Span4Mux_v
    port map (
            O => \N__9870\,
            I => \N__9867\
        );

    \I__2325\ : Span4Mux_h
    port map (
            O => \N__9867\,
            I => \N__9864\
        );

    \I__2324\ : Span4Mux_v
    port map (
            O => \N__9864\,
            I => \N__9860\
        );

    \I__2323\ : InMux
    port map (
            O => \N__9863\,
            I => \N__9857\
        );

    \I__2322\ : Odrv4
    port map (
            O => \N__9860\,
            I => \DS_ENm\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__9857\,
            I => \DS_ENm\
        );

    \I__2320\ : InMux
    port map (
            O => \N__9852\,
            I => \N__9843\
        );

    \I__2319\ : InMux
    port map (
            O => \N__9851\,
            I => \N__9843\
        );

    \I__2318\ : InMux
    port map (
            O => \N__9850\,
            I => \N__9838\
        );

    \I__2317\ : InMux
    port map (
            O => \N__9849\,
            I => \N__9838\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__9848\,
            I => \N__9835\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__9843\,
            I => \N__9827\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__9838\,
            I => \N__9824\
        );

    \I__2313\ : InMux
    port map (
            O => \N__9835\,
            I => \N__9821\
        );

    \I__2312\ : InMux
    port map (
            O => \N__9834\,
            I => \N__9818\
        );

    \I__2311\ : InMux
    port map (
            O => \N__9833\,
            I => \N__9813\
        );

    \I__2310\ : InMux
    port map (
            O => \N__9832\,
            I => \N__9813\
        );

    \I__2309\ : InMux
    port map (
            O => \N__9831\,
            I => \N__9810\
        );

    \I__2308\ : InMux
    port map (
            O => \N__9830\,
            I => \N__9807\
        );

    \I__2307\ : Span4Mux_v
    port map (
            O => \N__9827\,
            I => \N__9804\
        );

    \I__2306\ : Span4Mux_v
    port map (
            O => \N__9824\,
            I => \N__9801\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__9821\,
            I => \N__9794\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__9818\,
            I => \N__9794\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__9813\,
            I => \N__9794\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__9810\,
            I => \N__9789\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__9807\,
            I => \N__9789\
        );

    \I__2300\ : Span4Mux_v
    port map (
            O => \N__9804\,
            I => \N__9786\
        );

    \I__2299\ : Span4Mux_v
    port map (
            O => \N__9801\,
            I => \N__9781\
        );

    \I__2298\ : Span4Mux_v
    port map (
            O => \N__9794\,
            I => \N__9781\
        );

    \I__2297\ : Span12Mux_s10_v
    port map (
            O => \N__9789\,
            I => \N__9778\
        );

    \I__2296\ : Span4Mux_h
    port map (
            O => \N__9786\,
            I => \N__9775\
        );

    \I__2295\ : Sp12to4
    port map (
            O => \N__9781\,
            I => \N__9772\
        );

    \I__2294\ : Span12Mux_h
    port map (
            O => \N__9778\,
            I => \N__9769\
        );

    \I__2293\ : Sp12to4
    port map (
            O => \N__9775\,
            I => \N__9764\
        );

    \I__2292\ : Span12Mux_h
    port map (
            O => \N__9772\,
            I => \N__9764\
        );

    \I__2291\ : Odrv12
    port map (
            O => \N__9769\,
            I => \A_c_0\
        );

    \I__2290\ : Odrv12
    port map (
            O => \N__9764\,
            I => \A_c_0\
        );

    \I__2289\ : CascadeMux
    port map (
            O => \N__9759\,
            I => \N__9755\
        );

    \I__2288\ : InMux
    port map (
            O => \N__9758\,
            I => \N__9750\
        );

    \I__2287\ : InMux
    port map (
            O => \N__9755\,
            I => \N__9750\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__9750\,
            I => \N__9744\
        );

    \I__2285\ : InMux
    port map (
            O => \N__9749\,
            I => \N__9740\
        );

    \I__2284\ : InMux
    port map (
            O => \N__9748\,
            I => \N__9737\
        );

    \I__2283\ : InMux
    port map (
            O => \N__9747\,
            I => \N__9734\
        );

    \I__2282\ : Span4Mux_v
    port map (
            O => \N__9744\,
            I => \N__9729\
        );

    \I__2281\ : InMux
    port map (
            O => \N__9743\,
            I => \N__9726\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__9740\,
            I => \N__9723\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__9737\,
            I => \N__9718\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__9734\,
            I => \N__9718\
        );

    \I__2277\ : InMux
    port map (
            O => \N__9733\,
            I => \N__9713\
        );

    \I__2276\ : InMux
    port map (
            O => \N__9732\,
            I => \N__9713\
        );

    \I__2275\ : Span4Mux_v
    port map (
            O => \N__9729\,
            I => \N__9707\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__9726\,
            I => \N__9707\
        );

    \I__2273\ : Span4Mux_v
    port map (
            O => \N__9723\,
            I => \N__9700\
        );

    \I__2272\ : Span4Mux_h
    port map (
            O => \N__9718\,
            I => \N__9700\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__9713\,
            I => \N__9700\
        );

    \I__2270\ : InMux
    port map (
            O => \N__9712\,
            I => \N__9697\
        );

    \I__2269\ : Span4Mux_v
    port map (
            O => \N__9707\,
            I => \N__9694\
        );

    \I__2268\ : Span4Mux_h
    port map (
            O => \N__9700\,
            I => \N__9691\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__9697\,
            I => \N__9688\
        );

    \I__2266\ : Span4Mux_v
    port map (
            O => \N__9694\,
            I => \N__9685\
        );

    \I__2265\ : Span4Mux_v
    port map (
            O => \N__9691\,
            I => \N__9682\
        );

    \I__2264\ : Span12Mux_v
    port map (
            O => \N__9688\,
            I => \N__9679\
        );

    \I__2263\ : Span4Mux_h
    port map (
            O => \N__9685\,
            I => \N__9676\
        );

    \I__2262\ : Span4Mux_h
    port map (
            O => \N__9682\,
            I => \N__9673\
        );

    \I__2261\ : Span12Mux_h
    port map (
            O => \N__9679\,
            I => \N__9670\
        );

    \I__2260\ : Sp12to4
    port map (
            O => \N__9676\,
            I => \N__9665\
        );

    \I__2259\ : Sp12to4
    port map (
            O => \N__9673\,
            I => \N__9665\
        );

    \I__2258\ : Odrv12
    port map (
            O => \N__9670\,
            I => \SIZ_c_0\
        );

    \I__2257\ : Odrv12
    port map (
            O => \N__9665\,
            I => \SIZ_c_0\
        );

    \I__2256\ : IoInMux
    port map (
            O => \N__9660\,
            I => \N__9657\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__9657\,
            I => \N__9654\
        );

    \I__2254\ : Span4Mux_s2_v
    port map (
            O => \N__9654\,
            I => \N__9651\
        );

    \I__2253\ : Span4Mux_h
    port map (
            O => \N__9651\,
            I => \N__9648\
        );

    \I__2252\ : Span4Mux_v
    port map (
            O => \N__9648\,
            I => \N__9645\
        );

    \I__2251\ : Odrv4
    port map (
            O => \N__9645\,
            I => \N_87\
        );

    \I__2250\ : InMux
    port map (
            O => \N__9642\,
            I => \N__9639\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__9639\,
            I => \N__9636\
        );

    \I__2248\ : Odrv4
    port map (
            O => \N__9636\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__2247\ : InMux
    port map (
            O => \N__9633\,
            I => \N__9630\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__9630\,
            I => \N__9627\
        );

    \I__2245\ : Span4Mux_h
    port map (
            O => \N__9627\,
            I => \N__9624\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__9624\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__2243\ : InMux
    port map (
            O => \N__9621\,
            I => \N__9618\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__9618\,
            I => \N__9615\
        );

    \I__2241\ : Span4Mux_h
    port map (
            O => \N__9615\,
            I => \N__9612\
        );

    \I__2240\ : Odrv4
    port map (
            O => \N__9612\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__2239\ : InMux
    port map (
            O => \N__9609\,
            I => \N__9606\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__9606\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2237\ : InMux
    port map (
            O => \N__9603\,
            I => \N__9600\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__9600\,
            I => \N__9594\
        );

    \I__2235\ : InMux
    port map (
            O => \N__9599\,
            I => \N__9591\
        );

    \I__2234\ : InMux
    port map (
            O => \N__9598\,
            I => \N__9588\
        );

    \I__2233\ : InMux
    port map (
            O => \N__9597\,
            I => \N__9585\
        );

    \I__2232\ : Span4Mux_v
    port map (
            O => \N__9594\,
            I => \N__9582\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__9591\,
            I => \N__9577\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__9588\,
            I => \N__9577\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__9585\,
            I => \N__9574\
        );

    \I__2228\ : Sp12to4
    port map (
            O => \N__9582\,
            I => \N__9571\
        );

    \I__2227\ : Span4Mux_v
    port map (
            O => \N__9577\,
            I => \N__9566\
        );

    \I__2226\ : Span4Mux_h
    port map (
            O => \N__9574\,
            I => \N__9566\
        );

    \I__2225\ : Span12Mux_h
    port map (
            O => \N__9571\,
            I => \N__9563\
        );

    \I__2224\ : Sp12to4
    port map (
            O => \N__9566\,
            I => \N__9560\
        );

    \I__2223\ : Span12Mux_v
    port map (
            O => \N__9563\,
            I => \N__9557\
        );

    \I__2222\ : Span12Mux_v
    port map (
            O => \N__9560\,
            I => \N__9554\
        );

    \I__2221\ : Odrv12
    port map (
            O => \N__9557\,
            I => \DRA_c_2\
        );

    \I__2220\ : Odrv12
    port map (
            O => \N__9554\,
            I => \DRA_c_2\
        );

    \I__2219\ : InMux
    port map (
            O => \N__9549\,
            I => \N__9546\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__9546\,
            I => \N__9543\
        );

    \I__2217\ : Odrv12
    port map (
            O => \N__9543\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__2216\ : IoInMux
    port map (
            O => \N__9540\,
            I => \N__9537\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__9537\,
            I => \N__9534\
        );

    \I__2214\ : Span4Mux_s2_v
    port map (
            O => \N__9534\,
            I => \N__9531\
        );

    \I__2213\ : Span4Mux_v
    port map (
            O => \N__9531\,
            I => \N__9528\
        );

    \I__2212\ : Span4Mux_v
    port map (
            O => \N__9528\,
            I => \N__9525\
        );

    \I__2211\ : Span4Mux_h
    port map (
            O => \N__9525\,
            I => \N__9522\
        );

    \I__2210\ : Odrv4
    port map (
            O => \N__9522\,
            I => \CASn_c\
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__9519\,
            I => \N__9508\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__9518\,
            I => \N__9505\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__9517\,
            I => \N__9498\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__9516\,
            I => \N__9495\
        );

    \I__2205\ : CascadeMux
    port map (
            O => \N__9515\,
            I => \N__9491\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__9514\,
            I => \N__9488\
        );

    \I__2203\ : CascadeMux
    port map (
            O => \N__9513\,
            I => \N__9484\
        );

    \I__2202\ : CascadeMux
    port map (
            O => \N__9512\,
            I => \N__9480\
        );

    \I__2201\ : CascadeMux
    port map (
            O => \N__9511\,
            I => \N__9477\
        );

    \I__2200\ : InMux
    port map (
            O => \N__9508\,
            I => \N__9467\
        );

    \I__2199\ : InMux
    port map (
            O => \N__9505\,
            I => \N__9467\
        );

    \I__2198\ : InMux
    port map (
            O => \N__9504\,
            I => \N__9458\
        );

    \I__2197\ : InMux
    port map (
            O => \N__9503\,
            I => \N__9458\
        );

    \I__2196\ : InMux
    port map (
            O => \N__9502\,
            I => \N__9458\
        );

    \I__2195\ : InMux
    port map (
            O => \N__9501\,
            I => \N__9458\
        );

    \I__2194\ : InMux
    port map (
            O => \N__9498\,
            I => \N__9455\
        );

    \I__2193\ : InMux
    port map (
            O => \N__9495\,
            I => \N__9450\
        );

    \I__2192\ : InMux
    port map (
            O => \N__9494\,
            I => \N__9450\
        );

    \I__2191\ : InMux
    port map (
            O => \N__9491\,
            I => \N__9447\
        );

    \I__2190\ : InMux
    port map (
            O => \N__9488\,
            I => \N__9444\
        );

    \I__2189\ : InMux
    port map (
            O => \N__9487\,
            I => \N__9439\
        );

    \I__2188\ : InMux
    port map (
            O => \N__9484\,
            I => \N__9439\
        );

    \I__2187\ : InMux
    port map (
            O => \N__9483\,
            I => \N__9434\
        );

    \I__2186\ : InMux
    port map (
            O => \N__9480\,
            I => \N__9434\
        );

    \I__2185\ : InMux
    port map (
            O => \N__9477\,
            I => \N__9431\
        );

    \I__2184\ : InMux
    port map (
            O => \N__9476\,
            I => \N__9428\
        );

    \I__2183\ : InMux
    port map (
            O => \N__9475\,
            I => \N__9425\
        );

    \I__2182\ : InMux
    port map (
            O => \N__9474\,
            I => \N__9417\
        );

    \I__2181\ : InMux
    port map (
            O => \N__9473\,
            I => \N__9417\
        );

    \I__2180\ : InMux
    port map (
            O => \N__9472\,
            I => \N__9414\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__9467\,
            I => \N__9405\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__9458\,
            I => \N__9405\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__9455\,
            I => \N__9405\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__9450\,
            I => \N__9405\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__9447\,
            I => \N__9400\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__9444\,
            I => \N__9400\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__9439\,
            I => \N__9397\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__9434\,
            I => \N__9393\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__9431\,
            I => \N__9388\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__9428\,
            I => \N__9388\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__9425\,
            I => \N__9385\
        );

    \I__2168\ : InMux
    port map (
            O => \N__9424\,
            I => \N__9382\
        );

    \I__2167\ : InMux
    port map (
            O => \N__9423\,
            I => \N__9379\
        );

    \I__2166\ : InMux
    port map (
            O => \N__9422\,
            I => \N__9375\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__9417\,
            I => \N__9372\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__9414\,
            I => \N__9369\
        );

    \I__2163\ : Span4Mux_v
    port map (
            O => \N__9405\,
            I => \N__9366\
        );

    \I__2162\ : Span4Mux_h
    port map (
            O => \N__9400\,
            I => \N__9361\
        );

    \I__2161\ : Span4Mux_v
    port map (
            O => \N__9397\,
            I => \N__9361\
        );

    \I__2160\ : InMux
    port map (
            O => \N__9396\,
            I => \N__9358\
        );

    \I__2159\ : Span4Mux_v
    port map (
            O => \N__9393\,
            I => \N__9351\
        );

    \I__2158\ : Span4Mux_h
    port map (
            O => \N__9388\,
            I => \N__9351\
        );

    \I__2157\ : Span4Mux_h
    port map (
            O => \N__9385\,
            I => \N__9351\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__9382\,
            I => \N__9348\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__9379\,
            I => \N__9345\
        );

    \I__2154\ : InMux
    port map (
            O => \N__9378\,
            I => \N__9342\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__9375\,
            I => \N__9329\
        );

    \I__2152\ : Span12Mux_v
    port map (
            O => \N__9372\,
            I => \N__9329\
        );

    \I__2151\ : Span12Mux_h
    port map (
            O => \N__9369\,
            I => \N__9329\
        );

    \I__2150\ : Sp12to4
    port map (
            O => \N__9366\,
            I => \N__9329\
        );

    \I__2149\ : Sp12to4
    port map (
            O => \N__9361\,
            I => \N__9329\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__9358\,
            I => \N__9329\
        );

    \I__2147\ : Span4Mux_h
    port map (
            O => \N__9351\,
            I => \N__9326\
        );

    \I__2146\ : Span4Mux_v
    port map (
            O => \N__9348\,
            I => \N__9323\
        );

    \I__2145\ : Odrv4
    port map (
            O => \N__9345\,
            I => \CPU_CYCLEm\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__9342\,
            I => \CPU_CYCLEm\
        );

    \I__2143\ : Odrv12
    port map (
            O => \N__9329\,
            I => \CPU_CYCLEm\
        );

    \I__2142\ : Odrv4
    port map (
            O => \N__9326\,
            I => \CPU_CYCLEm\
        );

    \I__2141\ : Odrv4
    port map (
            O => \N__9323\,
            I => \CPU_CYCLEm\
        );

    \I__2140\ : InMux
    port map (
            O => \N__9312\,
            I => \N__9309\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__9309\,
            I => \N__9306\
        );

    \I__2138\ : Span12Mux_h
    port map (
            O => \N__9306\,
            I => \N__9303\
        );

    \I__2137\ : Odrv12
    port map (
            O => \N__9303\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__2136\ : CascadeMux
    port map (
            O => \N__9300\,
            I => \N__9296\
        );

    \I__2135\ : InMux
    port map (
            O => \N__9299\,
            I => \N__9291\
        );

    \I__2134\ : InMux
    port map (
            O => \N__9296\,
            I => \N__9288\
        );

    \I__2133\ : CascadeMux
    port map (
            O => \N__9295\,
            I => \N__9285\
        );

    \I__2132\ : InMux
    port map (
            O => \N__9294\,
            I => \N__9275\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__9291\,
            I => \N__9267\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__9288\,
            I => \N__9267\
        );

    \I__2129\ : InMux
    port map (
            O => \N__9285\,
            I => \N__9264\
        );

    \I__2128\ : InMux
    port map (
            O => \N__9284\,
            I => \N__9259\
        );

    \I__2127\ : InMux
    port map (
            O => \N__9283\,
            I => \N__9259\
        );

    \I__2126\ : InMux
    port map (
            O => \N__9282\,
            I => \N__9252\
        );

    \I__2125\ : InMux
    port map (
            O => \N__9281\,
            I => \N__9252\
        );

    \I__2124\ : InMux
    port map (
            O => \N__9280\,
            I => \N__9252\
        );

    \I__2123\ : InMux
    port map (
            O => \N__9279\,
            I => \N__9245\
        );

    \I__2122\ : InMux
    port map (
            O => \N__9278\,
            I => \N__9245\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__9275\,
            I => \N__9241\
        );

    \I__2120\ : InMux
    port map (
            O => \N__9274\,
            I => \N__9236\
        );

    \I__2119\ : InMux
    port map (
            O => \N__9273\,
            I => \N__9236\
        );

    \I__2118\ : CascadeMux
    port map (
            O => \N__9272\,
            I => \N__9232\
        );

    \I__2117\ : Span4Mux_v
    port map (
            O => \N__9267\,
            I => \N__9223\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__9264\,
            I => \N__9223\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__9259\,
            I => \N__9223\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__9252\,
            I => \N__9223\
        );

    \I__2113\ : InMux
    port map (
            O => \N__9251\,
            I => \N__9218\
        );

    \I__2112\ : InMux
    port map (
            O => \N__9250\,
            I => \N__9218\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__9245\,
            I => \N__9215\
        );

    \I__2110\ : CascadeMux
    port map (
            O => \N__9244\,
            I => \N__9210\
        );

    \I__2109\ : Span4Mux_v
    port map (
            O => \N__9241\,
            I => \N__9206\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__9236\,
            I => \N__9203\
        );

    \I__2107\ : InMux
    port map (
            O => \N__9235\,
            I => \N__9200\
        );

    \I__2106\ : InMux
    port map (
            O => \N__9232\,
            I => \N__9194\
        );

    \I__2105\ : Span4Mux_h
    port map (
            O => \N__9223\,
            I => \N__9187\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__9218\,
            I => \N__9187\
        );

    \I__2103\ : Span4Mux_v
    port map (
            O => \N__9215\,
            I => \N__9187\
        );

    \I__2102\ : InMux
    port map (
            O => \N__9214\,
            I => \N__9180\
        );

    \I__2101\ : InMux
    port map (
            O => \N__9213\,
            I => \N__9180\
        );

    \I__2100\ : InMux
    port map (
            O => \N__9210\,
            I => \N__9180\
        );

    \I__2099\ : InMux
    port map (
            O => \N__9209\,
            I => \N__9177\
        );

    \I__2098\ : Span4Mux_h
    port map (
            O => \N__9206\,
            I => \N__9170\
        );

    \I__2097\ : Span4Mux_v
    port map (
            O => \N__9203\,
            I => \N__9170\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__9200\,
            I => \N__9170\
        );

    \I__2095\ : InMux
    port map (
            O => \N__9199\,
            I => \N__9167\
        );

    \I__2094\ : InMux
    port map (
            O => \N__9198\,
            I => \N__9162\
        );

    \I__2093\ : InMux
    port map (
            O => \N__9197\,
            I => \N__9162\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__9194\,
            I => \N__9155\
        );

    \I__2091\ : Sp12to4
    port map (
            O => \N__9187\,
            I => \N__9155\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__9180\,
            I => \N__9155\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__9177\,
            I => \N__9150\
        );

    \I__2088\ : Span4Mux_h
    port map (
            O => \N__9170\,
            I => \N__9150\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__9167\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__9162\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2085\ : Odrv12
    port map (
            O => \N__9155\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2084\ : Odrv4
    port map (
            O => \N__9150\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2083\ : InMux
    port map (
            O => \N__9141\,
            I => \N__9138\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__9138\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__2081\ : IoInMux
    port map (
            O => \N__9135\,
            I => \N__9132\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__9132\,
            I => \N__9129\
        );

    \I__2079\ : Sp12to4
    port map (
            O => \N__9129\,
            I => \N__9126\
        );

    \I__2078\ : Span12Mux_h
    port map (
            O => \N__9126\,
            I => \N__9123\
        );

    \I__2077\ : Odrv12
    port map (
            O => \N__9123\,
            I => \CMA_c_4\
        );

    \I__2076\ : InMux
    port map (
            O => \N__9120\,
            I => \N__9117\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__9117\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__2074\ : IoInMux
    port map (
            O => \N__9114\,
            I => \N__9111\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__9111\,
            I => \N__9108\
        );

    \I__2072\ : Span4Mux_s2_h
    port map (
            O => \N__9108\,
            I => \N__9105\
        );

    \I__2071\ : Sp12to4
    port map (
            O => \N__9105\,
            I => \N__9102\
        );

    \I__2070\ : Span12Mux_v
    port map (
            O => \N__9102\,
            I => \N__9099\
        );

    \I__2069\ : Odrv12
    port map (
            O => \N__9099\,
            I => \CMA_c_7\
        );

    \I__2068\ : InMux
    port map (
            O => \N__9096\,
            I => \N__9091\
        );

    \I__2067\ : InMux
    port map (
            O => \N__9095\,
            I => \N__9086\
        );

    \I__2066\ : InMux
    port map (
            O => \N__9094\,
            I => \N__9086\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__9091\,
            I => \N__9079\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__9086\,
            I => \N__9079\
        );

    \I__2063\ : InMux
    port map (
            O => \N__9085\,
            I => \N__9076\
        );

    \I__2062\ : InMux
    port map (
            O => \N__9084\,
            I => \N__9070\
        );

    \I__2061\ : Span4Mux_h
    port map (
            O => \N__9079\,
            I => \N__9065\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__9076\,
            I => \N__9065\
        );

    \I__2059\ : InMux
    port map (
            O => \N__9075\,
            I => \N__9062\
        );

    \I__2058\ : InMux
    port map (
            O => \N__9074\,
            I => \N__9059\
        );

    \I__2057\ : InMux
    port map (
            O => \N__9073\,
            I => \N__9056\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__9070\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2055\ : Odrv4
    port map (
            O => \N__9065\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__9062\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__9059\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__9056\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2051\ : CascadeMux
    port map (
            O => \N__9045\,
            I => \N__9038\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__9044\,
            I => \N__9035\
        );

    \I__2049\ : CascadeMux
    port map (
            O => \N__9043\,
            I => \N__9032\
        );

    \I__2048\ : CascadeMux
    port map (
            O => \N__9042\,
            I => \N__9028\
        );

    \I__2047\ : InMux
    port map (
            O => \N__9041\,
            I => \N__9021\
        );

    \I__2046\ : InMux
    port map (
            O => \N__9038\,
            I => \N__9021\
        );

    \I__2045\ : InMux
    port map (
            O => \N__9035\,
            I => \N__9021\
        );

    \I__2044\ : InMux
    port map (
            O => \N__9032\,
            I => \N__9018\
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__9031\,
            I => \N__9015\
        );

    \I__2042\ : InMux
    port map (
            O => \N__9028\,
            I => \N__9012\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__9021\,
            I => \N__9007\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__9018\,
            I => \N__9007\
        );

    \I__2039\ : InMux
    port map (
            O => \N__9015\,
            I => \N__9004\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__9012\,
            I => \N__8999\
        );

    \I__2037\ : Span4Mux_v
    port map (
            O => \N__9007\,
            I => \N__8999\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__9004\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNIHMEAZ0Z_1\
        );

    \I__2035\ : Odrv4
    port map (
            O => \N__8999\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNIHMEAZ0Z_1\
        );

    \I__2034\ : InMux
    port map (
            O => \N__8994\,
            I => \N__8991\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__8991\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__2032\ : IoInMux
    port map (
            O => \N__8988\,
            I => \N__8985\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__8985\,
            I => \N__8982\
        );

    \I__2030\ : Span4Mux_s3_h
    port map (
            O => \N__8982\,
            I => \N__8979\
        );

    \I__2029\ : Sp12to4
    port map (
            O => \N__8979\,
            I => \N__8976\
        );

    \I__2028\ : Span12Mux_v
    port map (
            O => \N__8976\,
            I => \N__8973\
        );

    \I__2027\ : Odrv12
    port map (
            O => \N__8973\,
            I => \CMA_c_6\
        );

    \I__2026\ : InMux
    port map (
            O => \N__8970\,
            I => \N__8967\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__8967\,
            I => \N__8940\
        );

    \I__2024\ : ClkMux
    port map (
            O => \N__8966\,
            I => \N__8844\
        );

    \I__2023\ : ClkMux
    port map (
            O => \N__8965\,
            I => \N__8844\
        );

    \I__2022\ : ClkMux
    port map (
            O => \N__8964\,
            I => \N__8844\
        );

    \I__2021\ : ClkMux
    port map (
            O => \N__8963\,
            I => \N__8844\
        );

    \I__2020\ : ClkMux
    port map (
            O => \N__8962\,
            I => \N__8844\
        );

    \I__2019\ : ClkMux
    port map (
            O => \N__8961\,
            I => \N__8844\
        );

    \I__2018\ : ClkMux
    port map (
            O => \N__8960\,
            I => \N__8844\
        );

    \I__2017\ : ClkMux
    port map (
            O => \N__8959\,
            I => \N__8844\
        );

    \I__2016\ : ClkMux
    port map (
            O => \N__8958\,
            I => \N__8844\
        );

    \I__2015\ : ClkMux
    port map (
            O => \N__8957\,
            I => \N__8844\
        );

    \I__2014\ : ClkMux
    port map (
            O => \N__8956\,
            I => \N__8844\
        );

    \I__2013\ : ClkMux
    port map (
            O => \N__8955\,
            I => \N__8844\
        );

    \I__2012\ : ClkMux
    port map (
            O => \N__8954\,
            I => \N__8844\
        );

    \I__2011\ : ClkMux
    port map (
            O => \N__8953\,
            I => \N__8844\
        );

    \I__2010\ : ClkMux
    port map (
            O => \N__8952\,
            I => \N__8844\
        );

    \I__2009\ : ClkMux
    port map (
            O => \N__8951\,
            I => \N__8844\
        );

    \I__2008\ : ClkMux
    port map (
            O => \N__8950\,
            I => \N__8844\
        );

    \I__2007\ : ClkMux
    port map (
            O => \N__8949\,
            I => \N__8844\
        );

    \I__2006\ : ClkMux
    port map (
            O => \N__8948\,
            I => \N__8844\
        );

    \I__2005\ : ClkMux
    port map (
            O => \N__8947\,
            I => \N__8844\
        );

    \I__2004\ : ClkMux
    port map (
            O => \N__8946\,
            I => \N__8844\
        );

    \I__2003\ : ClkMux
    port map (
            O => \N__8945\,
            I => \N__8844\
        );

    \I__2002\ : ClkMux
    port map (
            O => \N__8944\,
            I => \N__8844\
        );

    \I__2001\ : ClkMux
    port map (
            O => \N__8943\,
            I => \N__8844\
        );

    \I__2000\ : Glb2LocalMux
    port map (
            O => \N__8940\,
            I => \N__8844\
        );

    \I__1999\ : ClkMux
    port map (
            O => \N__8939\,
            I => \N__8844\
        );

    \I__1998\ : ClkMux
    port map (
            O => \N__8938\,
            I => \N__8844\
        );

    \I__1997\ : ClkMux
    port map (
            O => \N__8937\,
            I => \N__8844\
        );

    \I__1996\ : ClkMux
    port map (
            O => \N__8936\,
            I => \N__8844\
        );

    \I__1995\ : ClkMux
    port map (
            O => \N__8935\,
            I => \N__8844\
        );

    \I__1994\ : ClkMux
    port map (
            O => \N__8934\,
            I => \N__8844\
        );

    \I__1993\ : ClkMux
    port map (
            O => \N__8933\,
            I => \N__8844\
        );

    \I__1992\ : ClkMux
    port map (
            O => \N__8932\,
            I => \N__8844\
        );

    \I__1991\ : ClkMux
    port map (
            O => \N__8931\,
            I => \N__8844\
        );

    \I__1990\ : ClkMux
    port map (
            O => \N__8930\,
            I => \N__8844\
        );

    \I__1989\ : ClkMux
    port map (
            O => \N__8929\,
            I => \N__8844\
        );

    \I__1988\ : ClkMux
    port map (
            O => \N__8928\,
            I => \N__8844\
        );

    \I__1987\ : ClkMux
    port map (
            O => \N__8927\,
            I => \N__8844\
        );

    \I__1986\ : ClkMux
    port map (
            O => \N__8926\,
            I => \N__8844\
        );

    \I__1985\ : ClkMux
    port map (
            O => \N__8925\,
            I => \N__8844\
        );

    \I__1984\ : GlobalMux
    port map (
            O => \N__8844\,
            I => \CLK80_PLL\
        );

    \I__1983\ : CEMux
    port map (
            O => \N__8841\,
            I => \N__8838\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__8838\,
            I => \N__8832\
        );

    \I__1981\ : CEMux
    port map (
            O => \N__8837\,
            I => \N__8828\
        );

    \I__1980\ : CEMux
    port map (
            O => \N__8836\,
            I => \N__8825\
        );

    \I__1979\ : CEMux
    port map (
            O => \N__8835\,
            I => \N__8822\
        );

    \I__1978\ : Span4Mux_h
    port map (
            O => \N__8832\,
            I => \N__8819\
        );

    \I__1977\ : CEMux
    port map (
            O => \N__8831\,
            I => \N__8816\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__8828\,
            I => \N__8812\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__8825\,
            I => \N__8807\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__8822\,
            I => \N__8807\
        );

    \I__1973\ : Span4Mux_h
    port map (
            O => \N__8819\,
            I => \N__8802\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__8816\,
            I => \N__8802\
        );

    \I__1971\ : CEMux
    port map (
            O => \N__8815\,
            I => \N__8799\
        );

    \I__1970\ : Span4Mux_v
    port map (
            O => \N__8812\,
            I => \N__8796\
        );

    \I__1969\ : Sp12to4
    port map (
            O => \N__8807\,
            I => \N__8793\
        );

    \I__1968\ : Sp12to4
    port map (
            O => \N__8802\,
            I => \N__8788\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__8799\,
            I => \N__8788\
        );

    \I__1966\ : Odrv4
    port map (
            O => \N__8796\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1965\ : Odrv12
    port map (
            O => \N__8793\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1964\ : Odrv12
    port map (
            O => \N__8788\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1963\ : InMux
    port map (
            O => \N__8781\,
            I => \N__8778\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__8778\,
            I => \N__8775\
        );

    \I__1961\ : Span12Mux_h
    port map (
            O => \N__8775\,
            I => \N__8772\
        );

    \I__1960\ : Odrv12
    port map (
            O => \N__8772\,
            I => \RAS0n_c\
        );

    \I__1959\ : InMux
    port map (
            O => \N__8769\,
            I => \N__8766\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__8766\,
            I => \N__8763\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__8763\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__1956\ : InMux
    port map (
            O => \N__8760\,
            I => \N__8754\
        );

    \I__1955\ : InMux
    port map (
            O => \N__8759\,
            I => \N__8754\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__8754\,
            I => \N__8751\
        );

    \I__1953\ : Span4Mux_v
    port map (
            O => \N__8751\,
            I => \N__8748\
        );

    \I__1952\ : Span4Mux_h
    port map (
            O => \N__8748\,
            I => \N__8745\
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__8745\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__1950\ : CascadeMux
    port map (
            O => \N__8742\,
            I => \N__8739\
        );

    \I__1949\ : InMux
    port map (
            O => \N__8739\,
            I => \N__8736\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__8736\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__1947\ : InMux
    port map (
            O => \N__8733\,
            I => \N__8730\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__8730\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__1945\ : IoInMux
    port map (
            O => \N__8727\,
            I => \N__8724\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__8724\,
            I => \N__8721\
        );

    \I__1943\ : Span4Mux_s0_v
    port map (
            O => \N__8721\,
            I => \N__8718\
        );

    \I__1942\ : Span4Mux_v
    port map (
            O => \N__8718\,
            I => \N__8715\
        );

    \I__1941\ : Span4Mux_v
    port map (
            O => \N__8715\,
            I => \N__8712\
        );

    \I__1940\ : Span4Mux_v
    port map (
            O => \N__8712\,
            I => \N__8709\
        );

    \I__1939\ : Odrv4
    port map (
            O => \N__8709\,
            I => \CMA_c_0\
        );

    \I__1938\ : InMux
    port map (
            O => \N__8706\,
            I => \N__8703\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__8703\,
            I => \N__8700\
        );

    \I__1936\ : Span4Mux_h
    port map (
            O => \N__8700\,
            I => \N__8697\
        );

    \I__1935\ : Odrv4
    port map (
            O => \N__8697\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\
        );

    \I__1934\ : InMux
    port map (
            O => \N__8694\,
            I => \N__8691\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__8691\,
            I => \N__8688\
        );

    \I__1932\ : Span4Mux_v
    port map (
            O => \N__8688\,
            I => \N__8685\
        );

    \I__1931\ : Sp12to4
    port map (
            O => \N__8685\,
            I => \N__8682\
        );

    \I__1930\ : Span12Mux_h
    port map (
            O => \N__8682\,
            I => \N__8679\
        );

    \I__1929\ : Odrv12
    port map (
            O => \N__8679\,
            I => \A_c_13\
        );

    \I__1928\ : InMux
    port map (
            O => \N__8676\,
            I => \N__8673\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__8673\,
            I => \N__8670\
        );

    \I__1926\ : Span4Mux_h
    port map (
            O => \N__8670\,
            I => \N__8667\
        );

    \I__1925\ : Span4Mux_v
    port map (
            O => \N__8667\,
            I => \N__8664\
        );

    \I__1924\ : Sp12to4
    port map (
            O => \N__8664\,
            I => \N__8661\
        );

    \I__1923\ : Span12Mux_h
    port map (
            O => \N__8661\,
            I => \N__8658\
        );

    \I__1922\ : Odrv12
    port map (
            O => \N__8658\,
            I => \A_c_6\
        );

    \I__1921\ : CascadeMux
    port map (
            O => \N__8655\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\
        );

    \I__1920\ : InMux
    port map (
            O => \N__8652\,
            I => \N__8649\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__8649\,
            I => \N__8645\
        );

    \I__1918\ : InMux
    port map (
            O => \N__8648\,
            I => \N__8642\
        );

    \I__1917\ : Span4Mux_h
    port map (
            O => \N__8645\,
            I => \N__8639\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__8642\,
            I => \N__8636\
        );

    \I__1915\ : Span4Mux_h
    port map (
            O => \N__8639\,
            I => \N__8631\
        );

    \I__1914\ : Span4Mux_v
    port map (
            O => \N__8636\,
            I => \N__8631\
        );

    \I__1913\ : Odrv4
    port map (
            O => \N__8631\,
            I => \DBRn_c_i\
        );

    \I__1912\ : InMux
    port map (
            O => \N__8628\,
            I => \N__8625\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__8625\,
            I => \N__8621\
        );

    \I__1910\ : InMux
    port map (
            O => \N__8624\,
            I => \N__8618\
        );

    \I__1909\ : Span12Mux_h
    port map (
            O => \N__8621\,
            I => \N__8615\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__8618\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__1907\ : Odrv12
    port map (
            O => \N__8615\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__1906\ : IoInMux
    port map (
            O => \N__8610\,
            I => \N__8607\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__8607\,
            I => \N__8604\
        );

    \I__1904\ : Span12Mux_s7_v
    port map (
            O => \N__8604\,
            I => \N__8601\
        );

    \I__1903\ : Odrv12
    port map (
            O => \N__8601\,
            I => \UMBEn_c\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__8598\,
            I => \N__8595\
        );

    \I__1901\ : InMux
    port map (
            O => \N__8595\,
            I => \N__8587\
        );

    \I__1900\ : InMux
    port map (
            O => \N__8594\,
            I => \N__8587\
        );

    \I__1899\ : InMux
    port map (
            O => \N__8593\,
            I => \N__8582\
        );

    \I__1898\ : InMux
    port map (
            O => \N__8592\,
            I => \N__8582\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__8587\,
            I => \N__8578\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__8582\,
            I => \N__8575\
        );

    \I__1895\ : CascadeMux
    port map (
            O => \N__8581\,
            I => \N__8571\
        );

    \I__1894\ : Span4Mux_v
    port map (
            O => \N__8578\,
            I => \N__8567\
        );

    \I__1893\ : Span4Mux_v
    port map (
            O => \N__8575\,
            I => \N__8564\
        );

    \I__1892\ : InMux
    port map (
            O => \N__8574\,
            I => \N__8561\
        );

    \I__1891\ : InMux
    port map (
            O => \N__8571\,
            I => \N__8556\
        );

    \I__1890\ : InMux
    port map (
            O => \N__8570\,
            I => \N__8556\
        );

    \I__1889\ : Span4Mux_v
    port map (
            O => \N__8567\,
            I => \N__8553\
        );

    \I__1888\ : Span4Mux_v
    port map (
            O => \N__8564\,
            I => \N__8550\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__8561\,
            I => \N__8545\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__8556\,
            I => \N__8545\
        );

    \I__1885\ : Span4Mux_v
    port map (
            O => \N__8553\,
            I => \N__8541\
        );

    \I__1884\ : Span4Mux_v
    port map (
            O => \N__8550\,
            I => \N__8536\
        );

    \I__1883\ : Span4Mux_v
    port map (
            O => \N__8545\,
            I => \N__8536\
        );

    \I__1882\ : InMux
    port map (
            O => \N__8544\,
            I => \N__8533\
        );

    \I__1881\ : Sp12to4
    port map (
            O => \N__8541\,
            I => \N__8526\
        );

    \I__1880\ : Sp12to4
    port map (
            O => \N__8536\,
            I => \N__8526\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__8533\,
            I => \N__8526\
        );

    \I__1878\ : Span12Mux_h
    port map (
            O => \N__8526\,
            I => \N__8523\
        );

    \I__1877\ : Odrv12
    port map (
            O => \N__8523\,
            I => \A_c_1\
        );

    \I__1876\ : CascadeMux
    port map (
            O => \N__8520\,
            I => \N__8517\
        );

    \I__1875\ : InMux
    port map (
            O => \N__8517\,
            I => \N__8512\
        );

    \I__1874\ : InMux
    port map (
            O => \N__8516\,
            I => \N__8509\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8515\,
            I => \N__8506\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__8512\,
            I => \N__8502\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__8509\,
            I => \N__8499\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__8506\,
            I => \N__8496\
        );

    \I__1869\ : CascadeMux
    port map (
            O => \N__8505\,
            I => \N__8492\
        );

    \I__1868\ : Span4Mux_v
    port map (
            O => \N__8502\,
            I => \N__8489\
        );

    \I__1867\ : Span4Mux_v
    port map (
            O => \N__8499\,
            I => \N__8484\
        );

    \I__1866\ : Span4Mux_h
    port map (
            O => \N__8496\,
            I => \N__8484\
        );

    \I__1865\ : InMux
    port map (
            O => \N__8495\,
            I => \N__8479\
        );

    \I__1864\ : InMux
    port map (
            O => \N__8492\,
            I => \N__8479\
        );

    \I__1863\ : Span4Mux_v
    port map (
            O => \N__8489\,
            I => \N__8476\
        );

    \I__1862\ : Span4Mux_v
    port map (
            O => \N__8484\,
            I => \N__8473\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__8479\,
            I => \N__8470\
        );

    \I__1860\ : Sp12to4
    port map (
            O => \N__8476\,
            I => \N__8463\
        );

    \I__1859\ : Sp12to4
    port map (
            O => \N__8473\,
            I => \N__8463\
        );

    \I__1858\ : Span12Mux_v
    port map (
            O => \N__8470\,
            I => \N__8463\
        );

    \I__1857\ : Span12Mux_h
    port map (
            O => \N__8463\,
            I => \N__8460\
        );

    \I__1856\ : Odrv12
    port map (
            O => \N__8460\,
            I => \SIZ_c_1\
        );

    \I__1855\ : IoInMux
    port map (
            O => \N__8457\,
            I => \N__8454\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__8454\,
            I => \N__8451\
        );

    \I__1853\ : Span4Mux_s3_v
    port map (
            O => \N__8451\,
            I => \N__8448\
        );

    \I__1852\ : Odrv4
    port map (
            O => \N__8448\,
            I => \N_276_i\
        );

    \I__1851\ : InMux
    port map (
            O => \N__8445\,
            I => \N__8441\
        );

    \I__1850\ : InMux
    port map (
            O => \N__8444\,
            I => \N__8438\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__8441\,
            I => \N__8434\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__8438\,
            I => \N__8430\
        );

    \I__1847\ : InMux
    port map (
            O => \N__8437\,
            I => \N__8427\
        );

    \I__1846\ : Span4Mux_h
    port map (
            O => \N__8434\,
            I => \N__8424\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__8433\,
            I => \N__8419\
        );

    \I__1844\ : Span4Mux_h
    port map (
            O => \N__8430\,
            I => \N__8414\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__8427\,
            I => \N__8414\
        );

    \I__1842\ : Span4Mux_v
    port map (
            O => \N__8424\,
            I => \N__8411\
        );

    \I__1841\ : InMux
    port map (
            O => \N__8423\,
            I => \N__8408\
        );

    \I__1840\ : InMux
    port map (
            O => \N__8422\,
            I => \N__8405\
        );

    \I__1839\ : InMux
    port map (
            O => \N__8419\,
            I => \N__8401\
        );

    \I__1838\ : Span4Mux_h
    port map (
            O => \N__8414\,
            I => \N__8398\
        );

    \I__1837\ : Sp12to4
    port map (
            O => \N__8411\,
            I => \N__8391\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__8408\,
            I => \N__8391\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__8405\,
            I => \N__8391\
        );

    \I__1834\ : InMux
    port map (
            O => \N__8404\,
            I => \N__8388\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__8401\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__8398\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1831\ : Odrv12
    port map (
            O => \N__8391\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8388\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1829\ : IoInMux
    port map (
            O => \N__8379\,
            I => \N__8376\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__8376\,
            I => \N__8373\
        );

    \I__1827\ : Span4Mux_s2_v
    port map (
            O => \N__8373\,
            I => \N__8370\
        );

    \I__1826\ : Span4Mux_v
    port map (
            O => \N__8370\,
            I => \N__8367\
        );

    \I__1825\ : Span4Mux_h
    port map (
            O => \N__8367\,
            I => \N__8364\
        );

    \I__1824\ : Odrv4
    port map (
            O => \N__8364\,
            I => \RASn_c\
        );

    \I__1823\ : CascadeMux
    port map (
            O => \N__8361\,
            I => \N__8358\
        );

    \I__1822\ : InMux
    port map (
            O => \N__8358\,
            I => \N__8354\
        );

    \I__1821\ : InMux
    port map (
            O => \N__8357\,
            I => \N__8351\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__8354\,
            I => \N__8348\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__8351\,
            I => \N__8341\
        );

    \I__1818\ : Sp12to4
    port map (
            O => \N__8348\,
            I => \N__8341\
        );

    \I__1817\ : InMux
    port map (
            O => \N__8347\,
            I => \N__8338\
        );

    \I__1816\ : InMux
    port map (
            O => \N__8346\,
            I => \N__8334\
        );

    \I__1815\ : Span12Mux_v
    port map (
            O => \N__8341\,
            I => \N__8329\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__8338\,
            I => \N__8329\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8337\,
            I => \N__8326\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__8334\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1811\ : Odrv12
    port map (
            O => \N__8329\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__8326\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1809\ : IoInMux
    port map (
            O => \N__8319\,
            I => \N__8316\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__8316\,
            I => \N__8313\
        );

    \I__1807\ : Span4Mux_s2_v
    port map (
            O => \N__8313\,
            I => \N__8310\
        );

    \I__1806\ : Span4Mux_v
    port map (
            O => \N__8310\,
            I => \N__8307\
        );

    \I__1805\ : Span4Mux_h
    port map (
            O => \N__8307\,
            I => \N__8304\
        );

    \I__1804\ : Odrv4
    port map (
            O => \N__8304\,
            I => \CRCSn_c\
        );

    \I__1803\ : InMux
    port map (
            O => \N__8301\,
            I => \N__8298\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__8298\,
            I => \U712_BYTE_ENABLE.N_339\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8295\,
            I => \N__8289\
        );

    \I__1800\ : InMux
    port map (
            O => \N__8294\,
            I => \N__8289\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__8289\,
            I => \N__8286\
        );

    \I__1798\ : Span4Mux_v
    port map (
            O => \N__8286\,
            I => \N__8281\
        );

    \I__1797\ : InMux
    port map (
            O => \N__8285\,
            I => \N__8276\
        );

    \I__1796\ : InMux
    port map (
            O => \N__8284\,
            I => \N__8276\
        );

    \I__1795\ : Span4Mux_v
    port map (
            O => \N__8281\,
            I => \N__8273\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__8276\,
            I => \N__8270\
        );

    \I__1793\ : Odrv4
    port map (
            O => \N__8273\,
            I => \U712_BYTE_ENABLE.N_206_i\
        );

    \I__1792\ : Odrv12
    port map (
            O => \N__8270\,
            I => \U712_BYTE_ENABLE.N_206_i\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8265\,
            I => \N__8262\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__8262\,
            I => \N__8259\
        );

    \I__1789\ : Span4Mux_h
    port map (
            O => \N__8259\,
            I => \N__8256\
        );

    \I__1788\ : Odrv4
    port map (
            O => \N__8256\,
            I => \U712_BYTE_ENABLE.N_316\
        );

    \I__1787\ : IoInMux
    port map (
            O => \N__8253\,
            I => \N__8250\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__8250\,
            I => \N__8247\
        );

    \I__1785\ : Span4Mux_s3_v
    port map (
            O => \N__8247\,
            I => \N__8244\
        );

    \I__1784\ : Odrv4
    port map (
            O => \N__8244\,
            I => \N_277_i\
        );

    \I__1783\ : IoInMux
    port map (
            O => \N__8241\,
            I => \N__8238\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__8238\,
            I => \N__8235\
        );

    \I__1781\ : Span4Mux_s2_v
    port map (
            O => \N__8235\,
            I => \N__8232\
        );

    \I__1780\ : Span4Mux_v
    port map (
            O => \N__8232\,
            I => \N__8229\
        );

    \I__1779\ : Odrv4
    port map (
            O => \N__8229\,
            I => \LLBE_i_o2_i\
        );

    \I__1778\ : IoInMux
    port map (
            O => \N__8226\,
            I => \N__8223\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__8223\,
            I => \N__8220\
        );

    \I__1776\ : IoSpan4Mux
    port map (
            O => \N__8220\,
            I => \N__8217\
        );

    \I__1775\ : Sp12to4
    port map (
            O => \N__8217\,
            I => \N__8214\
        );

    \I__1774\ : Span12Mux_s7_v
    port map (
            O => \N__8214\,
            I => \N__8211\
        );

    \I__1773\ : Span12Mux_h
    port map (
            O => \N__8211\,
            I => \N__8208\
        );

    \I__1772\ : Odrv12
    port map (
            O => \N__8208\,
            I => \WEn_c\
        );

    \I__1771\ : InMux
    port map (
            O => \N__8205\,
            I => \N__8202\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__8202\,
            I => \N__8199\
        );

    \I__1769\ : Sp12to4
    port map (
            O => \N__8199\,
            I => \N__8196\
        );

    \I__1768\ : Span12Mux_v
    port map (
            O => \N__8196\,
            I => \N__8193\
        );

    \I__1767\ : Span12Mux_h
    port map (
            O => \N__8193\,
            I => \N__8190\
        );

    \I__1766\ : Odrv12
    port map (
            O => \N__8190\,
            I => \A_c_17\
        );

    \I__1765\ : IoInMux
    port map (
            O => \N__8187\,
            I => \N__8184\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8184\,
            I => \N__8181\
        );

    \I__1763\ : IoSpan4Mux
    port map (
            O => \N__8181\,
            I => \N__8178\
        );

    \I__1762\ : IoSpan4Mux
    port map (
            O => \N__8178\,
            I => \N__8175\
        );

    \I__1761\ : Span4Mux_s2_h
    port map (
            O => \N__8175\,
            I => \N__8172\
        );

    \I__1760\ : Sp12to4
    port map (
            O => \N__8172\,
            I => \N__8169\
        );

    \I__1759\ : Odrv12
    port map (
            O => \N__8169\,
            I => \CMA_c_8\
        );

    \I__1758\ : InMux
    port map (
            O => \N__8166\,
            I => \N__8163\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__8163\,
            I => \N__8160\
        );

    \I__1756\ : Sp12to4
    port map (
            O => \N__8160\,
            I => \N__8157\
        );

    \I__1755\ : Span12Mux_v
    port map (
            O => \N__8157\,
            I => \N__8154\
        );

    \I__1754\ : Span12Mux_h
    port map (
            O => \N__8154\,
            I => \N__8151\
        );

    \I__1753\ : Odrv12
    port map (
            O => \N__8151\,
            I => \A_c_19\
        );

    \I__1752\ : InMux
    port map (
            O => \N__8148\,
            I => \N__8142\
        );

    \I__1751\ : InMux
    port map (
            O => \N__8147\,
            I => \N__8142\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__8142\,
            I => \N__8139\
        );

    \I__1749\ : Span4Mux_h
    port map (
            O => \N__8139\,
            I => \N__8134\
        );

    \I__1748\ : InMux
    port map (
            O => \N__8138\,
            I => \N__8129\
        );

    \I__1747\ : InMux
    port map (
            O => \N__8137\,
            I => \N__8129\
        );

    \I__1746\ : Odrv4
    port map (
            O => \N__8134\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__8129\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1744\ : IoInMux
    port map (
            O => \N__8124\,
            I => \N__8121\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__8121\,
            I => \N__8118\
        );

    \I__1742\ : IoSpan4Mux
    port map (
            O => \N__8118\,
            I => \N__8115\
        );

    \I__1741\ : Span4Mux_s3_h
    port map (
            O => \N__8115\,
            I => \N__8112\
        );

    \I__1740\ : Sp12to4
    port map (
            O => \N__8112\,
            I => \N__8109\
        );

    \I__1739\ : Span12Mux_h
    port map (
            O => \N__8109\,
            I => \N__8106\
        );

    \I__1738\ : Odrv12
    port map (
            O => \N__8106\,
            I => \CMA_c_9\
        );

    \I__1737\ : InMux
    port map (
            O => \N__8103\,
            I => \N__8098\
        );

    \I__1736\ : InMux
    port map (
            O => \N__8102\,
            I => \N__8094\
        );

    \I__1735\ : CascadeMux
    port map (
            O => \N__8101\,
            I => \N__8090\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__8098\,
            I => \N__8086\
        );

    \I__1733\ : InMux
    port map (
            O => \N__8097\,
            I => \N__8083\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__8094\,
            I => \N__8080\
        );

    \I__1731\ : InMux
    port map (
            O => \N__8093\,
            I => \N__8077\
        );

    \I__1730\ : InMux
    port map (
            O => \N__8090\,
            I => \N__8073\
        );

    \I__1729\ : InMux
    port map (
            O => \N__8089\,
            I => \N__8070\
        );

    \I__1728\ : Span4Mux_h
    port map (
            O => \N__8086\,
            I => \N__8065\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__8083\,
            I => \N__8065\
        );

    \I__1726\ : Span4Mux_v
    port map (
            O => \N__8080\,
            I => \N__8062\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__8077\,
            I => \N__8059\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__8076\,
            I => \N__8056\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__8073\,
            I => \N__8053\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__8070\,
            I => \N__8048\
        );

    \I__1721\ : Span4Mux_v
    port map (
            O => \N__8065\,
            I => \N__8048\
        );

    \I__1720\ : Span4Mux_h
    port map (
            O => \N__8062\,
            I => \N__8043\
        );

    \I__1719\ : Span4Mux_h
    port map (
            O => \N__8059\,
            I => \N__8043\
        );

    \I__1718\ : InMux
    port map (
            O => \N__8056\,
            I => \N__8040\
        );

    \I__1717\ : Odrv4
    port map (
            O => \N__8053\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1716\ : Odrv4
    port map (
            O => \N__8048\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1715\ : Odrv4
    port map (
            O => \N__8043\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__8040\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1713\ : IoInMux
    port map (
            O => \N__8031\,
            I => \N__8028\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__8028\,
            I => \N__8025\
        );

    \I__1711\ : Span4Mux_s3_v
    port map (
            O => \N__8025\,
            I => \N__8022\
        );

    \I__1710\ : Span4Mux_v
    port map (
            O => \N__8022\,
            I => \N__8019\
        );

    \I__1709\ : Span4Mux_v
    port map (
            O => \N__8019\,
            I => \N__8016\
        );

    \I__1708\ : Span4Mux_h
    port map (
            O => \N__8016\,
            I => \N__8013\
        );

    \I__1707\ : Odrv4
    port map (
            O => \N__8013\,
            I => \CMA_c_10\
        );

    \I__1706\ : InMux
    port map (
            O => \N__8010\,
            I => \N__8007\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__8007\,
            I => \U712_BYTE_ENABLE.N_320\
        );

    \I__1704\ : CascadeMux
    port map (
            O => \N__8004\,
            I => \U712_BYTE_ENABLE.N_318_cascade_\
        );

    \I__1703\ : IoInMux
    port map (
            O => \N__8001\,
            I => \N__7998\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__7998\,
            I => \N__7995\
        );

    \I__1701\ : IoSpan4Mux
    port map (
            O => \N__7995\,
            I => \N__7992\
        );

    \I__1700\ : Span4Mux_s3_h
    port map (
            O => \N__7992\,
            I => \N__7989\
        );

    \I__1699\ : Sp12to4
    port map (
            O => \N__7989\,
            I => \N__7986\
        );

    \I__1698\ : Span12Mux_s10_v
    port map (
            O => \N__7986\,
            I => \N__7983\
        );

    \I__1697\ : Span12Mux_h
    port map (
            O => \N__7983\,
            I => \N__7980\
        );

    \I__1696\ : Odrv12
    port map (
            O => \N__7980\,
            I => \N_105_i\
        );

    \I__1695\ : IoInMux
    port map (
            O => \N__7977\,
            I => \N__7974\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__7974\,
            I => \N__7971\
        );

    \I__1693\ : Span4Mux_s3_v
    port map (
            O => \N__7971\,
            I => \N__7968\
        );

    \I__1692\ : Span4Mux_v
    port map (
            O => \N__7968\,
            I => \N__7965\
        );

    \I__1691\ : Span4Mux_v
    port map (
            O => \N__7965\,
            I => \N__7962\
        );

    \I__1690\ : Odrv4
    port map (
            O => \N__7962\,
            I => \CMA_c_2\
        );

    \I__1689\ : InMux
    port map (
            O => \N__7959\,
            I => \N__7956\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__7956\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i\
        );

    \I__1687\ : InMux
    port map (
            O => \N__7953\,
            I => \N__7950\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__7950\,
            I => \N__7947\
        );

    \I__1685\ : Span12Mux_v
    port map (
            O => \N__7947\,
            I => \N__7944\
        );

    \I__1684\ : Span12Mux_h
    port map (
            O => \N__7944\,
            I => \N__7941\
        );

    \I__1683\ : Odrv12
    port map (
            O => \N__7941\,
            I => \A_c_4\
        );

    \I__1682\ : InMux
    port map (
            O => \N__7938\,
            I => \N__7935\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__7935\,
            I => \N__7932\
        );

    \I__1680\ : Span4Mux_v
    port map (
            O => \N__7932\,
            I => \N__7929\
        );

    \I__1679\ : Sp12to4
    port map (
            O => \N__7929\,
            I => \N__7926\
        );

    \I__1678\ : Span12Mux_h
    port map (
            O => \N__7926\,
            I => \N__7923\
        );

    \I__1677\ : Odrv12
    port map (
            O => \N__7923\,
            I => \A_c_11\
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__7920\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\
        );

    \I__1675\ : InMux
    port map (
            O => \N__7917\,
            I => \N__7914\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__7914\,
            I => \N__7911\
        );

    \I__1673\ : Odrv4
    port map (
            O => \N__7911\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__1672\ : InMux
    port map (
            O => \N__7908\,
            I => \N__7905\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__7905\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\
        );

    \I__1670\ : InMux
    port map (
            O => \N__7902\,
            I => \N__7894\
        );

    \I__1669\ : InMux
    port map (
            O => \N__7901\,
            I => \N__7889\
        );

    \I__1668\ : InMux
    port map (
            O => \N__7900\,
            I => \N__7889\
        );

    \I__1667\ : InMux
    port map (
            O => \N__7899\,
            I => \N__7886\
        );

    \I__1666\ : InMux
    port map (
            O => \N__7898\,
            I => \N__7883\
        );

    \I__1665\ : InMux
    port map (
            O => \N__7897\,
            I => \N__7880\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__7894\,
            I => \N__7877\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__7889\,
            I => \N__7871\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__7886\,
            I => \N__7871\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__7883\,
            I => \N__7868\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__7880\,
            I => \N__7865\
        );

    \I__1659\ : Span4Mux_v
    port map (
            O => \N__7877\,
            I => \N__7861\
        );

    \I__1658\ : InMux
    port map (
            O => \N__7876\,
            I => \N__7858\
        );

    \I__1657\ : Span4Mux_v
    port map (
            O => \N__7871\,
            I => \N__7853\
        );

    \I__1656\ : Span4Mux_v
    port map (
            O => \N__7868\,
            I => \N__7853\
        );

    \I__1655\ : Span4Mux_h
    port map (
            O => \N__7865\,
            I => \N__7850\
        );

    \I__1654\ : InMux
    port map (
            O => \N__7864\,
            I => \N__7847\
        );

    \I__1653\ : Odrv4
    port map (
            O => \N__7861\,
            I => \DMA_CYCLEm\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__7858\,
            I => \DMA_CYCLEm\
        );

    \I__1651\ : Odrv4
    port map (
            O => \N__7853\,
            I => \DMA_CYCLEm\
        );

    \I__1650\ : Odrv4
    port map (
            O => \N__7850\,
            I => \DMA_CYCLEm\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__7847\,
            I => \DMA_CYCLEm\
        );

    \I__1648\ : InMux
    port map (
            O => \N__7836\,
            I => \N__7833\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__7833\,
            I => \N__7828\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__7832\,
            I => \N__7824\
        );

    \I__1645\ : CascadeMux
    port map (
            O => \N__7831\,
            I => \N__7820\
        );

    \I__1644\ : Span4Mux_v
    port map (
            O => \N__7828\,
            I => \N__7817\
        );

    \I__1643\ : InMux
    port map (
            O => \N__7827\,
            I => \N__7814\
        );

    \I__1642\ : InMux
    port map (
            O => \N__7824\,
            I => \N__7811\
        );

    \I__1641\ : InMux
    port map (
            O => \N__7823\,
            I => \N__7808\
        );

    \I__1640\ : InMux
    port map (
            O => \N__7820\,
            I => \N__7805\
        );

    \I__1639\ : Span4Mux_v
    port map (
            O => \N__7817\,
            I => \N__7800\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__7814\,
            I => \N__7800\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__7811\,
            I => \N__7797\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__7808\,
            I => \N__7794\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__7805\,
            I => \N__7790\
        );

    \I__1634\ : Span4Mux_v
    port map (
            O => \N__7800\,
            I => \N__7787\
        );

    \I__1633\ : Span4Mux_v
    port map (
            O => \N__7797\,
            I => \N__7782\
        );

    \I__1632\ : Span4Mux_v
    port map (
            O => \N__7794\,
            I => \N__7782\
        );

    \I__1631\ : InMux
    port map (
            O => \N__7793\,
            I => \N__7779\
        );

    \I__1630\ : Span12Mux_v
    port map (
            O => \N__7790\,
            I => \N__7776\
        );

    \I__1629\ : Span4Mux_v
    port map (
            O => \N__7787\,
            I => \N__7773\
        );

    \I__1628\ : Sp12to4
    port map (
            O => \N__7782\,
            I => \N__7770\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__7779\,
            I => \N__7767\
        );

    \I__1626\ : Span12Mux_h
    port map (
            O => \N__7776\,
            I => \N__7764\
        );

    \I__1625\ : Sp12to4
    port map (
            O => \N__7773\,
            I => \N__7761\
        );

    \I__1624\ : Span12Mux_h
    port map (
            O => \N__7770\,
            I => \N__7758\
        );

    \I__1623\ : Span12Mux_v
    port map (
            O => \N__7767\,
            I => \N__7755\
        );

    \I__1622\ : Span12Mux_v
    port map (
            O => \N__7764\,
            I => \N__7752\
        );

    \I__1621\ : Span12Mux_h
    port map (
            O => \N__7761\,
            I => \N__7749\
        );

    \I__1620\ : Span12Mux_v
    port map (
            O => \N__7758\,
            I => \N__7744\
        );

    \I__1619\ : Span12Mux_h
    port map (
            O => \N__7755\,
            I => \N__7744\
        );

    \I__1618\ : Odrv12
    port map (
            O => \N__7752\,
            I => \CASUn_c\
        );

    \I__1617\ : Odrv12
    port map (
            O => \N__7749\,
            I => \CASUn_c\
        );

    \I__1616\ : Odrv12
    port map (
            O => \N__7744\,
            I => \CASUn_c\
        );

    \I__1615\ : IoInMux
    port map (
            O => \N__7737\,
            I => \N__7734\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__7734\,
            I => \N__7730\
        );

    \I__1613\ : InMux
    port map (
            O => \N__7733\,
            I => \N__7727\
        );

    \I__1612\ : IoSpan4Mux
    port map (
            O => \N__7730\,
            I => \N__7721\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__7727\,
            I => \N__7718\
        );

    \I__1610\ : InMux
    port map (
            O => \N__7726\,
            I => \N__7713\
        );

    \I__1609\ : InMux
    port map (
            O => \N__7725\,
            I => \N__7713\
        );

    \I__1608\ : InMux
    port map (
            O => \N__7724\,
            I => \N__7710\
        );

    \I__1607\ : Span4Mux_s2_v
    port map (
            O => \N__7721\,
            I => \N__7707\
        );

    \I__1606\ : Span4Mux_v
    port map (
            O => \N__7718\,
            I => \N__7700\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__7713\,
            I => \N__7700\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__7710\,
            I => \N__7700\
        );

    \I__1603\ : Span4Mux_v
    port map (
            O => \N__7707\,
            I => \N__7697\
        );

    \I__1602\ : Span4Mux_h
    port map (
            O => \N__7700\,
            I => \N__7694\
        );

    \I__1601\ : Span4Mux_v
    port map (
            O => \N__7697\,
            I => \N__7688\
        );

    \I__1600\ : Span4Mux_v
    port map (
            O => \N__7694\,
            I => \N__7688\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7693\,
            I => \N__7685\
        );

    \I__1598\ : Odrv4
    port map (
            O => \N__7688\,
            I => \DBENn_c\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__7685\,
            I => \DBENn_c\
        );

    \I__1596\ : IoInMux
    port map (
            O => \N__7680\,
            I => \N__7677\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__7677\,
            I => \N__7674\
        );

    \I__1594\ : IoSpan4Mux
    port map (
            O => \N__7674\,
            I => \N__7671\
        );

    \I__1593\ : Span4Mux_s3_h
    port map (
            O => \N__7671\,
            I => \N__7668\
        );

    \I__1592\ : Sp12to4
    port map (
            O => \N__7668\,
            I => \N__7665\
        );

    \I__1591\ : Span12Mux_h
    port map (
            O => \N__7665\,
            I => \N__7662\
        );

    \I__1590\ : Odrv12
    port map (
            O => \N__7662\,
            I => \N_57_i\
        );

    \I__1589\ : CascadeMux
    port map (
            O => \N__7659\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_\
        );

    \I__1588\ : InMux
    port map (
            O => \N__7656\,
            I => \N__7653\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__7653\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__1586\ : InMux
    port map (
            O => \N__7650\,
            I => \N__7647\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__7647\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\
        );

    \I__1584\ : InMux
    port map (
            O => \N__7644\,
            I => \N__7641\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__7641\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\
        );

    \I__1582\ : InMux
    port map (
            O => \N__7638\,
            I => \N__7635\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__7635\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\
        );

    \I__1580\ : IoInMux
    port map (
            O => \N__7632\,
            I => \N__7629\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__7629\,
            I => \N__7626\
        );

    \I__1578\ : Span4Mux_s3_h
    port map (
            O => \N__7626\,
            I => \N__7623\
        );

    \I__1577\ : Span4Mux_v
    port map (
            O => \N__7623\,
            I => \N__7620\
        );

    \I__1576\ : Sp12to4
    port map (
            O => \N__7620\,
            I => \N__7617\
        );

    \I__1575\ : Span12Mux_h
    port map (
            O => \N__7617\,
            I => \N__7614\
        );

    \I__1574\ : Odrv12
    port map (
            O => \N__7614\,
            I => \CMA_c_5\
        );

    \I__1573\ : InMux
    port map (
            O => \N__7611\,
            I => \N__7608\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__7608\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\
        );

    \I__1571\ : InMux
    port map (
            O => \N__7605\,
            I => \N__7602\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__7602\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\
        );

    \I__1569\ : InMux
    port map (
            O => \N__7599\,
            I => \N__7596\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__7596\,
            I => \N__7593\
        );

    \I__1567\ : Span4Mux_v
    port map (
            O => \N__7593\,
            I => \N__7590\
        );

    \I__1566\ : Sp12to4
    port map (
            O => \N__7590\,
            I => \N__7587\
        );

    \I__1565\ : Span12Mux_h
    port map (
            O => \N__7587\,
            I => \N__7584\
        );

    \I__1564\ : Span12Mux_v
    port map (
            O => \N__7584\,
            I => \N__7581\
        );

    \I__1563\ : Odrv12
    port map (
            O => \N__7581\,
            I => \A_c_2\
        );

    \I__1562\ : InMux
    port map (
            O => \N__7578\,
            I => \N__7575\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__7575\,
            I => \N__7572\
        );

    \I__1560\ : Span4Mux_v
    port map (
            O => \N__7572\,
            I => \N__7569\
        );

    \I__1559\ : Sp12to4
    port map (
            O => \N__7569\,
            I => \N__7566\
        );

    \I__1558\ : Span12Mux_h
    port map (
            O => \N__7566\,
            I => \N__7563\
        );

    \I__1557\ : Odrv12
    port map (
            O => \N__7563\,
            I => \A_c_9\
        );

    \I__1556\ : InMux
    port map (
            O => \N__7560\,
            I => \N__7557\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__7557\,
            I => \N__7554\
        );

    \I__1554\ : Span4Mux_v
    port map (
            O => \N__7554\,
            I => \N__7547\
        );

    \I__1553\ : InMux
    port map (
            O => \N__7553\,
            I => \N__7544\
        );

    \I__1552\ : CascadeMux
    port map (
            O => \N__7552\,
            I => \N__7541\
        );

    \I__1551\ : InMux
    port map (
            O => \N__7551\,
            I => \N__7536\
        );

    \I__1550\ : InMux
    port map (
            O => \N__7550\,
            I => \N__7536\
        );

    \I__1549\ : Span4Mux_v
    port map (
            O => \N__7547\,
            I => \N__7531\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__7544\,
            I => \N__7531\
        );

    \I__1547\ : InMux
    port map (
            O => \N__7541\,
            I => \N__7528\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__7536\,
            I => \N__7524\
        );

    \I__1545\ : Span4Mux_v
    port map (
            O => \N__7531\,
            I => \N__7521\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__7528\,
            I => \N__7518\
        );

    \I__1543\ : InMux
    port map (
            O => \N__7527\,
            I => \N__7515\
        );

    \I__1542\ : Span4Mux_v
    port map (
            O => \N__7524\,
            I => \N__7512\
        );

    \I__1541\ : Span4Mux_h
    port map (
            O => \N__7521\,
            I => \N__7507\
        );

    \I__1540\ : Span4Mux_v
    port map (
            O => \N__7518\,
            I => \N__7507\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__7515\,
            I => \N__7504\
        );

    \I__1538\ : Sp12to4
    port map (
            O => \N__7512\,
            I => \N__7501\
        );

    \I__1537\ : Span4Mux_v
    port map (
            O => \N__7507\,
            I => \N__7498\
        );

    \I__1536\ : Span12Mux_v
    port map (
            O => \N__7504\,
            I => \N__7495\
        );

    \I__1535\ : Span12Mux_h
    port map (
            O => \N__7501\,
            I => \N__7492\
        );

    \I__1534\ : Sp12to4
    port map (
            O => \N__7498\,
            I => \N__7489\
        );

    \I__1533\ : Span12Mux_h
    port map (
            O => \N__7495\,
            I => \N__7486\
        );

    \I__1532\ : Span12Mux_v
    port map (
            O => \N__7492\,
            I => \N__7481\
        );

    \I__1531\ : Span12Mux_h
    port map (
            O => \N__7489\,
            I => \N__7481\
        );

    \I__1530\ : Odrv12
    port map (
            O => \N__7486\,
            I => \CASLn_c\
        );

    \I__1529\ : Odrv12
    port map (
            O => \N__7481\,
            I => \CASLn_c\
        );

    \I__1528\ : InMux
    port map (
            O => \N__7476\,
            I => \N__7473\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7473\,
            I => \U712_BYTE_ENABLE.N_342\
        );

    \I__1526\ : CascadeMux
    port map (
            O => \N__7470\,
            I => \U712_BYTE_ENABLE.N_341_cascade_\
        );

    \I__1525\ : IoInMux
    port map (
            O => \N__7467\,
            I => \N__7464\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__7464\,
            I => \N__7461\
        );

    \I__1523\ : Span4Mux_s2_v
    port map (
            O => \N__7461\,
            I => \N__7458\
        );

    \I__1522\ : Span4Mux_h
    port map (
            O => \N__7458\,
            I => \N__7455\
        );

    \I__1521\ : Sp12to4
    port map (
            O => \N__7455\,
            I => \N__7452\
        );

    \I__1520\ : Span12Mux_v
    port map (
            O => \N__7452\,
            I => \N__7449\
        );

    \I__1519\ : Odrv12
    port map (
            O => \N__7449\,
            I => \N_55_i\
        );

    \I__1518\ : InMux
    port map (
            O => \N__7446\,
            I => \N__7443\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__7443\,
            I => \N__7440\
        );

    \I__1516\ : Odrv12
    port map (
            O => \N__7440\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\
        );

    \I__1515\ : InMux
    port map (
            O => \N__7437\,
            I => \N__7434\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__7434\,
            I => \N__7431\
        );

    \I__1513\ : Span4Mux_v
    port map (
            O => \N__7431\,
            I => \N__7428\
        );

    \I__1512\ : Sp12to4
    port map (
            O => \N__7428\,
            I => \N__7425\
        );

    \I__1511\ : Span12Mux_h
    port map (
            O => \N__7425\,
            I => \N__7422\
        );

    \I__1510\ : Span12Mux_v
    port map (
            O => \N__7422\,
            I => \N__7419\
        );

    \I__1509\ : Odrv12
    port map (
            O => \N__7419\,
            I => \A_c_3\
        );

    \I__1508\ : InMux
    port map (
            O => \N__7416\,
            I => \N__7413\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__7413\,
            I => \N__7410\
        );

    \I__1506\ : Span4Mux_v
    port map (
            O => \N__7410\,
            I => \N__7407\
        );

    \I__1505\ : Sp12to4
    port map (
            O => \N__7407\,
            I => \N__7404\
        );

    \I__1504\ : Span12Mux_h
    port map (
            O => \N__7404\,
            I => \N__7401\
        );

    \I__1503\ : Odrv12
    port map (
            O => \N__7401\,
            I => \A_c_10\
        );

    \I__1502\ : IoInMux
    port map (
            O => \N__7398\,
            I => \N__7395\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__7395\,
            I => \N__7392\
        );

    \I__1500\ : IoSpan4Mux
    port map (
            O => \N__7392\,
            I => \N__7389\
        );

    \I__1499\ : IoSpan4Mux
    port map (
            O => \N__7389\,
            I => \N__7386\
        );

    \I__1498\ : Span4Mux_s3_h
    port map (
            O => \N__7386\,
            I => \N__7383\
        );

    \I__1497\ : Sp12to4
    port map (
            O => \N__7383\,
            I => \N__7380\
        );

    \I__1496\ : Odrv12
    port map (
            O => \N__7380\,
            I => \N_180_i\
        );

    \I__1495\ : InMux
    port map (
            O => \N__7377\,
            I => \N__7367\
        );

    \I__1494\ : InMux
    port map (
            O => \N__7376\,
            I => \N__7367\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7375\,
            I => \N__7362\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7374\,
            I => \N__7362\
        );

    \I__1491\ : InMux
    port map (
            O => \N__7373\,
            I => \N__7357\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7372\,
            I => \N__7357\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__7367\,
            I => \N__7346\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__7362\,
            I => \N__7346\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__7357\,
            I => \N__7346\
        );

    \I__1486\ : InMux
    port map (
            O => \N__7356\,
            I => \N__7343\
        );

    \I__1485\ : InMux
    port map (
            O => \N__7355\,
            I => \N__7339\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7354\,
            I => \N__7336\
        );

    \I__1483\ : InMux
    port map (
            O => \N__7353\,
            I => \N__7333\
        );

    \I__1482\ : Span4Mux_h
    port map (
            O => \N__7346\,
            I => \N__7324\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__7343\,
            I => \N__7324\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7342\,
            I => \N__7321\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__7339\,
            I => \N__7318\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__7336\,
            I => \N__7315\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__7333\,
            I => \N__7312\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7332\,
            I => \N__7307\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7331\,
            I => \N__7307\
        );

    \I__1474\ : InMux
    port map (
            O => \N__7330\,
            I => \N__7304\
        );

    \I__1473\ : InMux
    port map (
            O => \N__7329\,
            I => \N__7301\
        );

    \I__1472\ : Span4Mux_h
    port map (
            O => \N__7324\,
            I => \N__7296\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__7321\,
            I => \N__7296\
        );

    \I__1470\ : Span4Mux_v
    port map (
            O => \N__7318\,
            I => \N__7293\
        );

    \I__1469\ : Span4Mux_v
    port map (
            O => \N__7315\,
            I => \N__7282\
        );

    \I__1468\ : Span4Mux_v
    port map (
            O => \N__7312\,
            I => \N__7282\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__7307\,
            I => \N__7282\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7304\,
            I => \N__7282\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__7301\,
            I => \N__7282\
        );

    \I__1464\ : Span4Mux_v
    port map (
            O => \N__7296\,
            I => \N__7278\
        );

    \I__1463\ : Span4Mux_v
    port map (
            O => \N__7293\,
            I => \N__7273\
        );

    \I__1462\ : Span4Mux_v
    port map (
            O => \N__7282\,
            I => \N__7273\
        );

    \I__1461\ : InMux
    port map (
            O => \N__7281\,
            I => \N__7270\
        );

    \I__1460\ : Sp12to4
    port map (
            O => \N__7278\,
            I => \N__7263\
        );

    \I__1459\ : Sp12to4
    port map (
            O => \N__7273\,
            I => \N__7263\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__7270\,
            I => \N__7263\
        );

    \I__1457\ : Span12Mux_h
    port map (
            O => \N__7263\,
            I => \N__7260\
        );

    \I__1456\ : Odrv12
    port map (
            O => \N__7260\,
            I => \RESETn_c\
        );

    \I__1455\ : IoInMux
    port map (
            O => \N__7257\,
            I => \N__7254\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__7254\,
            I => \N__7251\
        );

    \I__1453\ : Sp12to4
    port map (
            O => \N__7251\,
            I => \N__7248\
        );

    \I__1452\ : Odrv12
    port map (
            O => \N__7248\,
            I => \RESETn_c_i\
        );

    \I__1451\ : InMux
    port map (
            O => \N__7245\,
            I => \N__7242\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__7242\,
            I => \N__7239\
        );

    \I__1449\ : Odrv4
    port map (
            O => \N__7239\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__1448\ : IoInMux
    port map (
            O => \N__7236\,
            I => \N__7233\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__7233\,
            I => \N__7230\
        );

    \I__1446\ : IoSpan4Mux
    port map (
            O => \N__7230\,
            I => \N__7227\
        );

    \I__1445\ : Span4Mux_s1_h
    port map (
            O => \N__7227\,
            I => \N__7224\
        );

    \I__1444\ : Sp12to4
    port map (
            O => \N__7224\,
            I => \N__7221\
        );

    \I__1443\ : Span12Mux_h
    port map (
            O => \N__7221\,
            I => \N__7218\
        );

    \I__1442\ : Odrv12
    port map (
            O => \N__7218\,
            I => \CMA_c_3\
        );

    \I__1441\ : CascadeMux
    port map (
            O => \N__7215\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1_cascade_\
        );

    \I__1440\ : IoInMux
    port map (
            O => \N__7212\,
            I => \N__7209\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__7209\,
            I => \N__7206\
        );

    \I__1438\ : Span4Mux_s2_v
    port map (
            O => \N__7206\,
            I => \N__7203\
        );

    \I__1437\ : Sp12to4
    port map (
            O => \N__7203\,
            I => \N__7200\
        );

    \I__1436\ : Span12Mux_h
    port map (
            O => \N__7200\,
            I => \N__7197\
        );

    \I__1435\ : Odrv12
    port map (
            O => \N__7197\,
            I => \CMA_c_1\
        );

    \I__1434\ : SRMux
    port map (
            O => \N__7194\,
            I => \N__7191\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__7191\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__1432\ : InMux
    port map (
            O => \N__7188\,
            I => \N__7184\
        );

    \I__1431\ : InMux
    port map (
            O => \N__7187\,
            I => \N__7181\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__7184\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__7181\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1428\ : InMux
    port map (
            O => \N__7176\,
            I => \N__7172\
        );

    \I__1427\ : InMux
    port map (
            O => \N__7175\,
            I => \N__7169\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__7172\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__7169\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1424\ : InMux
    port map (
            O => \N__7164\,
            I => \N__7160\
        );

    \I__1423\ : InMux
    port map (
            O => \N__7163\,
            I => \N__7157\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__7160\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__7157\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__1420\ : InMux
    port map (
            O => \N__7152\,
            I => \N__7149\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__7149\,
            I => \N__7146\
        );

    \I__1418\ : Odrv4
    port map (
            O => \N__7146\,
            I => \U712_CHIP_RAM.REFRESH5lt7\
        );

    \I__1417\ : IoInMux
    port map (
            O => \N__7143\,
            I => \N__7140\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__7140\,
            I => \N__7137\
        );

    \I__1415\ : Span4Mux_s2_v
    port map (
            O => \N__7137\,
            I => \N__7133\
        );

    \I__1414\ : InMux
    port map (
            O => \N__7136\,
            I => \N__7130\
        );

    \I__1413\ : Span4Mux_v
    port map (
            O => \N__7133\,
            I => \N__7127\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__7130\,
            I => \N__7124\
        );

    \I__1411\ : Span4Mux_v
    port map (
            O => \N__7127\,
            I => \N__7121\
        );

    \I__1410\ : Span4Mux_v
    port map (
            O => \N__7124\,
            I => \N__7118\
        );

    \I__1409\ : Odrv4
    port map (
            O => \N__7121\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1408\ : Odrv4
    port map (
            O => \N__7118\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1407\ : InMux
    port map (
            O => \N__7113\,
            I => \N__7110\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__7110\,
            I => \N__7107\
        );

    \I__1405\ : Span12Mux_v
    port map (
            O => \N__7107\,
            I => \N__7104\
        );

    \I__1404\ : Span12Mux_h
    port map (
            O => \N__7104\,
            I => \N__7101\
        );

    \I__1403\ : Odrv12
    port map (
            O => \N__7101\,
            I => \A_c_7\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__7098\,
            I => \U712_CHIP_RAM.N_231_cascade_\
        );

    \I__1401\ : CascadeMux
    port map (
            O => \N__7095\,
            I => \N__7092\
        );

    \I__1400\ : InMux
    port map (
            O => \N__7092\,
            I => \N__7086\
        );

    \I__1399\ : InMux
    port map (
            O => \N__7091\,
            I => \N__7086\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__7086\,
            I => \N__7083\
        );

    \I__1397\ : Span4Mux_v
    port map (
            O => \N__7083\,
            I => \N__7080\
        );

    \I__1396\ : Span4Mux_v
    port map (
            O => \N__7080\,
            I => \N__7077\
        );

    \I__1395\ : Sp12to4
    port map (
            O => \N__7077\,
            I => \N__7074\
        );

    \I__1394\ : Span12Mux_h
    port map (
            O => \N__7074\,
            I => \N__7071\
        );

    \I__1393\ : Odrv12
    port map (
            O => \N__7071\,
            I => \A_c_14\
        );

    \I__1392\ : CascadeMux
    port map (
            O => \N__7068\,
            I => \N__7064\
        );

    \I__1391\ : InMux
    port map (
            O => \N__7067\,
            I => \N__7059\
        );

    \I__1390\ : InMux
    port map (
            O => \N__7064\,
            I => \N__7056\
        );

    \I__1389\ : InMux
    port map (
            O => \N__7063\,
            I => \N__7051\
        );

    \I__1388\ : InMux
    port map (
            O => \N__7062\,
            I => \N__7051\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__7059\,
            I => \N__7044\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__7056\,
            I => \N__7044\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__7051\,
            I => \N__7044\
        );

    \I__1384\ : Span4Mux_v
    port map (
            O => \N__7044\,
            I => \N__7041\
        );

    \I__1383\ : Span4Mux_v
    port map (
            O => \N__7041\,
            I => \N__7038\
        );

    \I__1382\ : Span4Mux_v
    port map (
            O => \N__7038\,
            I => \N__7035\
        );

    \I__1381\ : IoSpan4Mux
    port map (
            O => \N__7035\,
            I => \N__7032\
        );

    \I__1380\ : Odrv4
    port map (
            O => \N__7032\,
            I => \CLK40_PLL_i\
        );

    \I__1379\ : IoInMux
    port map (
            O => \N__7029\,
            I => \N__7026\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__7026\,
            I => \N__7022\
        );

    \I__1377\ : IoInMux
    port map (
            O => \N__7025\,
            I => \N__7019\
        );

    \I__1376\ : IoSpan4Mux
    port map (
            O => \N__7022\,
            I => \N__7013\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__7019\,
            I => \N__7013\
        );

    \I__1374\ : IoInMux
    port map (
            O => \N__7018\,
            I => \N__7010\
        );

    \I__1373\ : IoSpan4Mux
    port map (
            O => \N__7013\,
            I => \N__7007\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__7010\,
            I => \N__7004\
        );

    \I__1371\ : IoSpan4Mux
    port map (
            O => \N__7007\,
            I => \N__7001\
        );

    \I__1370\ : Span4Mux_s3_h
    port map (
            O => \N__7004\,
            I => \N__6998\
        );

    \I__1369\ : Sp12to4
    port map (
            O => \N__7001\,
            I => \N__6995\
        );

    \I__1368\ : Span4Mux_h
    port map (
            O => \N__6998\,
            I => \N__6992\
        );

    \I__1367\ : Span12Mux_s6_v
    port map (
            O => \N__6995\,
            I => \N__6989\
        );

    \I__1366\ : Span4Mux_h
    port map (
            O => \N__6992\,
            I => \N__6986\
        );

    \I__1365\ : Span12Mux_v
    port map (
            O => \N__6989\,
            I => \N__6983\
        );

    \I__1364\ : Span4Mux_h
    port map (
            O => \N__6986\,
            I => \N__6980\
        );

    \I__1363\ : Odrv12
    port map (
            O => \N__6983\,
            I => \CLK40_PLL_i_i\
        );

    \I__1362\ : Odrv4
    port map (
            O => \N__6980\,
            I => \CLK40_PLL_i_i\
        );

    \I__1361\ : InMux
    port map (
            O => \N__6975\,
            I => \N__6968\
        );

    \I__1360\ : InMux
    port map (
            O => \N__6974\,
            I => \N__6968\
        );

    \I__1359\ : InMux
    port map (
            O => \N__6973\,
            I => \N__6965\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__6968\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__6965\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1356\ : InMux
    port map (
            O => \N__6960\,
            I => \N__6956\
        );

    \I__1355\ : InMux
    port map (
            O => \N__6959\,
            I => \N__6953\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__6956\,
            I => \N__6950\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__6953\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__1352\ : Odrv4
    port map (
            O => \N__6950\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__1351\ : InMux
    port map (
            O => \N__6945\,
            I => \N__6942\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__6942\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\
        );

    \I__1349\ : InMux
    port map (
            O => \N__6939\,
            I => \N__6936\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__6936\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__1347\ : InMux
    port map (
            O => \N__6933\,
            I => \bfn_11_10_0_\
        );

    \I__1346\ : InMux
    port map (
            O => \N__6930\,
            I => \N__6927\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__6927\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__1344\ : InMux
    port map (
            O => \N__6924\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__1343\ : InMux
    port map (
            O => \N__6921\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__1342\ : InMux
    port map (
            O => \N__6918\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__1341\ : InMux
    port map (
            O => \N__6915\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__1340\ : InMux
    port map (
            O => \N__6912\,
            I => \N__6908\
        );

    \I__1339\ : InMux
    port map (
            O => \N__6911\,
            I => \N__6905\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__6908\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__6905\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1336\ : InMux
    port map (
            O => \N__6900\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__1335\ : InMux
    port map (
            O => \N__6897\,
            I => \N__6893\
        );

    \I__1334\ : InMux
    port map (
            O => \N__6896\,
            I => \N__6890\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__6893\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__6890\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1331\ : InMux
    port map (
            O => \N__6885\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__1330\ : InMux
    port map (
            O => \N__6882\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__1329\ : CascadeMux
    port map (
            O => \N__6879\,
            I => \N__6876\
        );

    \I__1328\ : InMux
    port map (
            O => \N__6876\,
            I => \N__6872\
        );

    \I__1327\ : InMux
    port map (
            O => \N__6875\,
            I => \N__6869\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__6872\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__6869\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1324\ : ClkMux
    port map (
            O => \N__6864\,
            I => \N__6846\
        );

    \I__1323\ : ClkMux
    port map (
            O => \N__6863\,
            I => \N__6846\
        );

    \I__1322\ : ClkMux
    port map (
            O => \N__6862\,
            I => \N__6846\
        );

    \I__1321\ : ClkMux
    port map (
            O => \N__6861\,
            I => \N__6846\
        );

    \I__1320\ : ClkMux
    port map (
            O => \N__6860\,
            I => \N__6846\
        );

    \I__1319\ : ClkMux
    port map (
            O => \N__6859\,
            I => \N__6846\
        );

    \I__1318\ : GlobalMux
    port map (
            O => \N__6846\,
            I => \N__6843\
        );

    \I__1317\ : gio2CtrlBuf
    port map (
            O => \N__6843\,
            I => \C1_c_g\
        );

    \I__1316\ : CascadeMux
    port map (
            O => \N__6840\,
            I => \N__6836\
        );

    \I__1315\ : InMux
    port map (
            O => \N__6839\,
            I => \N__6833\
        );

    \I__1314\ : InMux
    port map (
            O => \N__6836\,
            I => \N__6830\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__6833\,
            I => \N__6827\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__6830\,
            I => \U712_CHIP_RAM.N_314\
        );

    \I__1311\ : Odrv4
    port map (
            O => \N__6827\,
            I => \U712_CHIP_RAM.N_314\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__6822\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_cascade_\
        );

    \I__1309\ : InMux
    port map (
            O => \N__6819\,
            I => \N__6816\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__6816\,
            I => \U712_CHIP_RAM.N_37\
        );

    \I__1307\ : InMux
    port map (
            O => \N__6813\,
            I => \N__6809\
        );

    \I__1306\ : InMux
    port map (
            O => \N__6812\,
            I => \N__6806\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__6809\,
            I => \N__6803\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__6806\,
            I => \CPU_TACKm\
        );

    \I__1303\ : Odrv4
    port map (
            O => \N__6803\,
            I => \CPU_TACKm\
        );

    \I__1302\ : InMux
    port map (
            O => \N__6798\,
            I => \N__6794\
        );

    \I__1301\ : InMux
    port map (
            O => \N__6797\,
            I => \N__6787\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__6794\,
            I => \N__6781\
        );

    \I__1299\ : InMux
    port map (
            O => \N__6793\,
            I => \N__6778\
        );

    \I__1298\ : InMux
    port map (
            O => \N__6792\,
            I => \N__6775\
        );

    \I__1297\ : InMux
    port map (
            O => \N__6791\,
            I => \N__6770\
        );

    \I__1296\ : InMux
    port map (
            O => \N__6790\,
            I => \N__6770\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__6787\,
            I => \N__6765\
        );

    \I__1294\ : InMux
    port map (
            O => \N__6786\,
            I => \N__6762\
        );

    \I__1293\ : InMux
    port map (
            O => \N__6785\,
            I => \N__6759\
        );

    \I__1292\ : InMux
    port map (
            O => \N__6784\,
            I => \N__6756\
        );

    \I__1291\ : Span4Mux_v
    port map (
            O => \N__6781\,
            I => \N__6747\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__6778\,
            I => \N__6747\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__6775\,
            I => \N__6747\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__6770\,
            I => \N__6743\
        );

    \I__1287\ : InMux
    port map (
            O => \N__6769\,
            I => \N__6737\
        );

    \I__1286\ : InMux
    port map (
            O => \N__6768\,
            I => \N__6734\
        );

    \I__1285\ : Span4Mux_h
    port map (
            O => \N__6765\,
            I => \N__6729\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__6762\,
            I => \N__6729\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__6759\,
            I => \N__6724\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__6756\,
            I => \N__6724\
        );

    \I__1281\ : InMux
    port map (
            O => \N__6755\,
            I => \N__6721\
        );

    \I__1280\ : InMux
    port map (
            O => \N__6754\,
            I => \N__6718\
        );

    \I__1279\ : Span4Mux_h
    port map (
            O => \N__6747\,
            I => \N__6715\
        );

    \I__1278\ : InMux
    port map (
            O => \N__6746\,
            I => \N__6712\
        );

    \I__1277\ : Span4Mux_h
    port map (
            O => \N__6743\,
            I => \N__6709\
        );

    \I__1276\ : InMux
    port map (
            O => \N__6742\,
            I => \N__6702\
        );

    \I__1275\ : InMux
    port map (
            O => \N__6741\,
            I => \N__6702\
        );

    \I__1274\ : InMux
    port map (
            O => \N__6740\,
            I => \N__6702\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__6737\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__6734\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1271\ : Odrv4
    port map (
            O => \N__6729\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1270\ : Odrv4
    port map (
            O => \N__6724\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__6721\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__6718\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1267\ : Odrv4
    port map (
            O => \N__6715\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__6712\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1265\ : Odrv4
    port map (
            O => \N__6709\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__6702\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1263\ : InMux
    port map (
            O => \N__6681\,
            I => \N__6675\
        );

    \I__1262\ : InMux
    port map (
            O => \N__6680\,
            I => \N__6675\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__6675\,
            I => \U712_CHIP_RAM.N_396\
        );

    \I__1260\ : InMux
    port map (
            O => \N__6672\,
            I => \N__6669\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__6669\,
            I => \N__6666\
        );

    \I__1258\ : Span4Mux_h
    port map (
            O => \N__6666\,
            I => \N__6661\
        );

    \I__1257\ : InMux
    port map (
            O => \N__6665\,
            I => \N__6658\
        );

    \I__1256\ : InMux
    port map (
            O => \N__6664\,
            I => \N__6655\
        );

    \I__1255\ : Odrv4
    port map (
            O => \N__6661\,
            I => \U712_CHIP_RAM.N_400\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__6658\,
            I => \U712_CHIP_RAM.N_400\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__6655\,
            I => \U712_CHIP_RAM.N_400\
        );

    \I__1252\ : InMux
    port map (
            O => \N__6648\,
            I => \N__6644\
        );

    \I__1251\ : CascadeMux
    port map (
            O => \N__6647\,
            I => \N__6640\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__6644\,
            I => \N__6637\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6643\,
            I => \N__6633\
        );

    \I__1248\ : InMux
    port map (
            O => \N__6640\,
            I => \N__6630\
        );

    \I__1247\ : Span4Mux_h
    port map (
            O => \N__6637\,
            I => \N__6627\
        );

    \I__1246\ : InMux
    port map (
            O => \N__6636\,
            I => \N__6624\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__6633\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__6630\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1243\ : Odrv4
    port map (
            O => \N__6627\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__6624\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1241\ : CascadeMux
    port map (
            O => \N__6615\,
            I => \N__6611\
        );

    \I__1240\ : InMux
    port map (
            O => \N__6614\,
            I => \N__6607\
        );

    \I__1239\ : InMux
    port map (
            O => \N__6611\,
            I => \N__6604\
        );

    \I__1238\ : CascadeMux
    port map (
            O => \N__6610\,
            I => \N__6601\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__6607\,
            I => \N__6596\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__6604\,
            I => \N__6596\
        );

    \I__1235\ : InMux
    port map (
            O => \N__6601\,
            I => \N__6593\
        );

    \I__1234\ : Span4Mux_h
    port map (
            O => \N__6596\,
            I => \N__6590\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__6593\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1232\ : Odrv4
    port map (
            O => \N__6590\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1231\ : InMux
    port map (
            O => \N__6585\,
            I => \N__6579\
        );

    \I__1230\ : InMux
    port map (
            O => \N__6584\,
            I => \N__6572\
        );

    \I__1229\ : InMux
    port map (
            O => \N__6583\,
            I => \N__6572\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6582\,
            I => \N__6572\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__6579\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__6572\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1225\ : IoInMux
    port map (
            O => \N__6567\,
            I => \N__6564\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__6564\,
            I => \N__6561\
        );

    \I__1223\ : Span12Mux_s8_h
    port map (
            O => \N__6561\,
            I => \N__6558\
        );

    \I__1222\ : Span12Mux_v
    port map (
            O => \N__6558\,
            I => \N__6554\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6557\,
            I => \N__6551\
        );

    \I__1220\ : Odrv12
    port map (
            O => \N__6554\,
            I => \TACK_OUTn\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__6551\,
            I => \TACK_OUTn\
        );

    \I__1218\ : CascadeMux
    port map (
            O => \N__6546\,
            I => \N__6543\
        );

    \I__1217\ : InMux
    port map (
            O => \N__6543\,
            I => \N__6539\
        );

    \I__1216\ : InMux
    port map (
            O => \N__6542\,
            I => \N__6536\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__6539\,
            I => \N__6531\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__6536\,
            I => \N__6531\
        );

    \I__1213\ : Span4Mux_v
    port map (
            O => \N__6531\,
            I => \N__6527\
        );

    \I__1212\ : InMux
    port map (
            O => \N__6530\,
            I => \N__6524\
        );

    \I__1211\ : Odrv4
    port map (
            O => \N__6527\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__6524\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1209\ : InMux
    port map (
            O => \N__6519\,
            I => \N__6516\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__6516\,
            I => \N__6512\
        );

    \I__1207\ : InMux
    port map (
            O => \N__6515\,
            I => \N__6509\
        );

    \I__1206\ : Span4Mux_v
    port map (
            O => \N__6512\,
            I => \N__6506\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__6509\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1204\ : Odrv4
    port map (
            O => \N__6506\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1203\ : InMux
    port map (
            O => \N__6501\,
            I => \N__6493\
        );

    \I__1202\ : InMux
    port map (
            O => \N__6500\,
            I => \N__6490\
        );

    \I__1201\ : InMux
    port map (
            O => \N__6499\,
            I => \N__6487\
        );

    \I__1200\ : InMux
    port map (
            O => \N__6498\,
            I => \N__6484\
        );

    \I__1199\ : InMux
    port map (
            O => \N__6497\,
            I => \N__6479\
        );

    \I__1198\ : InMux
    port map (
            O => \N__6496\,
            I => \N__6479\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__6493\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__6490\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__6487\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__6484\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__6479\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1192\ : InMux
    port map (
            O => \N__6468\,
            I => \N__6464\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6467\,
            I => \N__6461\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__6464\,
            I => \U712_REG_SM.N_216\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__6461\,
            I => \U712_REG_SM.N_216\
        );

    \I__1188\ : InMux
    port map (
            O => \N__6456\,
            I => \N__6448\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6455\,
            I => \N__6445\
        );

    \I__1186\ : InMux
    port map (
            O => \N__6454\,
            I => \N__6442\
        );

    \I__1185\ : InMux
    port map (
            O => \N__6453\,
            I => \N__6435\
        );

    \I__1184\ : InMux
    port map (
            O => \N__6452\,
            I => \N__6435\
        );

    \I__1183\ : InMux
    port map (
            O => \N__6451\,
            I => \N__6435\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__6448\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__6445\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6442\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__6435\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1178\ : InMux
    port map (
            O => \N__6426\,
            I => \N__6422\
        );

    \I__1177\ : InMux
    port map (
            O => \N__6425\,
            I => \N__6419\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__6422\,
            I => \U712_REG_SM.N_239\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6419\,
            I => \U712_REG_SM.N_239\
        );

    \I__1174\ : CascadeMux
    port map (
            O => \N__6414\,
            I => \N__6411\
        );

    \I__1173\ : InMux
    port map (
            O => \N__6411\,
            I => \N__6406\
        );

    \I__1172\ : InMux
    port map (
            O => \N__6410\,
            I => \N__6400\
        );

    \I__1171\ : InMux
    port map (
            O => \N__6409\,
            I => \N__6400\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__6406\,
            I => \N__6394\
        );

    \I__1169\ : InMux
    port map (
            O => \N__6405\,
            I => \N__6387\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__6400\,
            I => \N__6384\
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__6399\,
            I => \N__6381\
        );

    \I__1166\ : InMux
    port map (
            O => \N__6398\,
            I => \N__6376\
        );

    \I__1165\ : InMux
    port map (
            O => \N__6397\,
            I => \N__6376\
        );

    \I__1164\ : Span4Mux_h
    port map (
            O => \N__6394\,
            I => \N__6373\
        );

    \I__1163\ : InMux
    port map (
            O => \N__6393\,
            I => \N__6368\
        );

    \I__1162\ : InMux
    port map (
            O => \N__6392\,
            I => \N__6368\
        );

    \I__1161\ : InMux
    port map (
            O => \N__6391\,
            I => \N__6363\
        );

    \I__1160\ : InMux
    port map (
            O => \N__6390\,
            I => \N__6363\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__6387\,
            I => \N__6358\
        );

    \I__1158\ : Span4Mux_h
    port map (
            O => \N__6384\,
            I => \N__6358\
        );

    \I__1157\ : InMux
    port map (
            O => \N__6381\,
            I => \N__6355\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__6376\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1155\ : Odrv4
    port map (
            O => \N__6373\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__6368\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__6363\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__6358\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__6355\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1150\ : IoInMux
    port map (
            O => \N__6342\,
            I => \N__6339\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__6339\,
            I => \N__6335\
        );

    \I__1148\ : IoInMux
    port map (
            O => \N__6338\,
            I => \N__6332\
        );

    \I__1147\ : Span4Mux_s2_v
    port map (
            O => \N__6335\,
            I => \N__6329\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__6332\,
            I => \N__6326\
        );

    \I__1145\ : Span4Mux_h
    port map (
            O => \N__6329\,
            I => \N__6323\
        );

    \I__1144\ : Span4Mux_s2_v
    port map (
            O => \N__6326\,
            I => \N__6320\
        );

    \I__1143\ : Sp12to4
    port map (
            O => \N__6323\,
            I => \N__6317\
        );

    \I__1142\ : Sp12to4
    port map (
            O => \N__6320\,
            I => \N__6314\
        );

    \I__1141\ : Span12Mux_h
    port map (
            O => \N__6317\,
            I => \N__6309\
        );

    \I__1140\ : Span12Mux_h
    port map (
            O => \N__6314\,
            I => \N__6309\
        );

    \I__1139\ : Odrv12
    port map (
            O => \N__6309\,
            I => \ASn_c\
        );

    \I__1138\ : CEMux
    port map (
            O => \N__6306\,
            I => \N__6303\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__6303\,
            I => \U712_REG_SM.N_239_0_0\
        );

    \I__1136\ : InMux
    port map (
            O => \N__6300\,
            I => \N__6295\
        );

    \I__1135\ : InMux
    port map (
            O => \N__6299\,
            I => \N__6292\
        );

    \I__1134\ : InMux
    port map (
            O => \N__6298\,
            I => \N__6289\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__6295\,
            I => \N__6284\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__6292\,
            I => \N__6284\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__6289\,
            I => \N__6280\
        );

    \I__1130\ : Span4Mux_v
    port map (
            O => \N__6284\,
            I => \N__6277\
        );

    \I__1129\ : InMux
    port map (
            O => \N__6283\,
            I => \N__6274\
        );

    \I__1128\ : Span4Mux_v
    port map (
            O => \N__6280\,
            I => \N__6271\
        );

    \I__1127\ : Span4Mux_v
    port map (
            O => \N__6277\,
            I => \N__6266\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__6274\,
            I => \N__6266\
        );

    \I__1125\ : Sp12to4
    port map (
            O => \N__6271\,
            I => \N__6263\
        );

    \I__1124\ : Span4Mux_v
    port map (
            O => \N__6266\,
            I => \N__6260\
        );

    \I__1123\ : Span12Mux_h
    port map (
            O => \N__6263\,
            I => \N__6257\
        );

    \I__1122\ : Sp12to4
    port map (
            O => \N__6260\,
            I => \N__6254\
        );

    \I__1121\ : Span12Mux_v
    port map (
            O => \N__6257\,
            I => \N__6249\
        );

    \I__1120\ : Span12Mux_h
    port map (
            O => \N__6254\,
            I => \N__6249\
        );

    \I__1119\ : Odrv12
    port map (
            O => \N__6249\,
            I => \RnW_c\
        );

    \I__1118\ : InMux
    port map (
            O => \N__6246\,
            I => \N__6243\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__6243\,
            I => \N__6239\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6242\,
            I => \N__6232\
        );

    \I__1115\ : Span4Mux_v
    port map (
            O => \N__6239\,
            I => \N__6229\
        );

    \I__1114\ : InMux
    port map (
            O => \N__6238\,
            I => \N__6226\
        );

    \I__1113\ : InMux
    port map (
            O => \N__6237\,
            I => \N__6223\
        );

    \I__1112\ : InMux
    port map (
            O => \N__6236\,
            I => \N__6218\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6235\,
            I => \N__6218\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6232\,
            I => \N__6214\
        );

    \I__1109\ : Span4Mux_v
    port map (
            O => \N__6229\,
            I => \N__6209\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__6226\,
            I => \N__6209\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__6223\,
            I => \N__6206\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__6218\,
            I => \N__6203\
        );

    \I__1105\ : InMux
    port map (
            O => \N__6217\,
            I => \N__6200\
        );

    \I__1104\ : Span12Mux_s11_v
    port map (
            O => \N__6214\,
            I => \N__6197\
        );

    \I__1103\ : Span4Mux_v
    port map (
            O => \N__6209\,
            I => \N__6188\
        );

    \I__1102\ : Span4Mux_v
    port map (
            O => \N__6206\,
            I => \N__6188\
        );

    \I__1101\ : Span4Mux_h
    port map (
            O => \N__6203\,
            I => \N__6188\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__6200\,
            I => \N__6188\
        );

    \I__1099\ : Odrv12
    port map (
            O => \N__6197\,
            I => \WRITE_CYCLEm\
        );

    \I__1098\ : Odrv4
    port map (
            O => \N__6188\,
            I => \WRITE_CYCLEm\
        );

    \I__1097\ : IoInMux
    port map (
            O => \N__6183\,
            I => \N__6180\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__6180\,
            I => \N__6177\
        );

    \I__1095\ : IoSpan4Mux
    port map (
            O => \N__6177\,
            I => \N__6174\
        );

    \I__1094\ : Span4Mux_s3_h
    port map (
            O => \N__6174\,
            I => \N__6171\
        );

    \I__1093\ : Span4Mux_h
    port map (
            O => \N__6171\,
            I => \N__6168\
        );

    \I__1092\ : Span4Mux_v
    port map (
            O => \N__6168\,
            I => \N__6165\
        );

    \I__1091\ : Sp12to4
    port map (
            O => \N__6165\,
            I => \N__6162\
        );

    \I__1090\ : Odrv12
    port map (
            O => \N__6162\,
            I => \N_259\
        );

    \I__1089\ : InMux
    port map (
            O => \N__6159\,
            I => \N__6151\
        );

    \I__1088\ : InMux
    port map (
            O => \N__6158\,
            I => \N__6148\
        );

    \I__1087\ : InMux
    port map (
            O => \N__6157\,
            I => \N__6144\
        );

    \I__1086\ : InMux
    port map (
            O => \N__6156\,
            I => \N__6141\
        );

    \I__1085\ : InMux
    port map (
            O => \N__6155\,
            I => \N__6136\
        );

    \I__1084\ : InMux
    port map (
            O => \N__6154\,
            I => \N__6136\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__6151\,
            I => \N__6131\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__6148\,
            I => \N__6131\
        );

    \I__1081\ : InMux
    port map (
            O => \N__6147\,
            I => \N__6128\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__6144\,
            I => \N__6123\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__6141\,
            I => \N__6123\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__6136\,
            I => \U712_CHIP_RAM.N_360\
        );

    \I__1077\ : Odrv4
    port map (
            O => \N__6131\,
            I => \U712_CHIP_RAM.N_360\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__6128\,
            I => \U712_CHIP_RAM.N_360\
        );

    \I__1075\ : Odrv4
    port map (
            O => \N__6123\,
            I => \U712_CHIP_RAM.N_360\
        );

    \I__1074\ : CEMux
    port map (
            O => \N__6114\,
            I => \N__6111\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__6111\,
            I => \N__6108\
        );

    \I__1072\ : Span4Mux_h
    port map (
            O => \N__6108\,
            I => \N__6105\
        );

    \I__1071\ : Odrv4
    port map (
            O => \N__6105\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0_0\
        );

    \I__1070\ : CascadeMux
    port map (
            O => \N__6102\,
            I => \N__6099\
        );

    \I__1069\ : InMux
    port map (
            O => \N__6099\,
            I => \N__6096\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__6096\,
            I => \U712_CHIP_RAM.CLK_EN_5_0\
        );

    \I__1067\ : IoInMux
    port map (
            O => \N__6093\,
            I => \N__6090\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__6090\,
            I => \N__6087\
        );

    \I__1065\ : Span4Mux_s3_h
    port map (
            O => \N__6087\,
            I => \N__6084\
        );

    \I__1064\ : Span4Mux_v
    port map (
            O => \N__6084\,
            I => \N__6081\
        );

    \I__1063\ : Sp12to4
    port map (
            O => \N__6081\,
            I => \N__6078\
        );

    \I__1062\ : Span12Mux_h
    port map (
            O => \N__6078\,
            I => \N__6074\
        );

    \I__1061\ : InMux
    port map (
            O => \N__6077\,
            I => \N__6071\
        );

    \I__1060\ : Odrv12
    port map (
            O => \N__6074\,
            I => \CLK_EN_c\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__6071\,
            I => \CLK_EN_c\
        );

    \I__1058\ : InMux
    port map (
            O => \N__6066\,
            I => \N__6062\
        );

    \I__1057\ : InMux
    port map (
            O => \N__6065\,
            I => \N__6059\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__6062\,
            I => \U712_CHIP_RAM.N_404\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__6059\,
            I => \U712_CHIP_RAM.N_404\
        );

    \I__1054\ : InMux
    port map (
            O => \N__6054\,
            I => \N__6048\
        );

    \I__1053\ : InMux
    port map (
            O => \N__6053\,
            I => \N__6048\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__6048\,
            I => \U712_CHIP_RAM.N_313_2\
        );

    \I__1051\ : CascadeMux
    port map (
            O => \N__6045\,
            I => \U712_CHIP_RAM.N_312_cascade_\
        );

    \I__1050\ : CascadeMux
    port map (
            O => \N__6042\,
            I => \N__6037\
        );

    \I__1049\ : InMux
    port map (
            O => \N__6041\,
            I => \N__6026\
        );

    \I__1048\ : InMux
    port map (
            O => \N__6040\,
            I => \N__6026\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6037\,
            I => \N__6023\
        );

    \I__1046\ : InMux
    port map (
            O => \N__6036\,
            I => \N__6018\
        );

    \I__1045\ : InMux
    port map (
            O => \N__6035\,
            I => \N__6015\
        );

    \I__1044\ : CascadeMux
    port map (
            O => \N__6034\,
            I => \N__6008\
        );

    \I__1043\ : CascadeMux
    port map (
            O => \N__6033\,
            I => \N__6002\
        );

    \I__1042\ : InMux
    port map (
            O => \N__6032\,
            I => \N__5996\
        );

    \I__1041\ : InMux
    port map (
            O => \N__6031\,
            I => \N__5996\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__6026\,
            I => \N__5992\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__6023\,
            I => \N__5989\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6022\,
            I => \N__5986\
        );

    \I__1037\ : InMux
    port map (
            O => \N__6021\,
            I => \N__5983\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__6018\,
            I => \N__5978\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__6015\,
            I => \N__5978\
        );

    \I__1034\ : InMux
    port map (
            O => \N__6014\,
            I => \N__5975\
        );

    \I__1033\ : InMux
    port map (
            O => \N__6013\,
            I => \N__5968\
        );

    \I__1032\ : InMux
    port map (
            O => \N__6012\,
            I => \N__5968\
        );

    \I__1031\ : InMux
    port map (
            O => \N__6011\,
            I => \N__5968\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6008\,
            I => \N__5961\
        );

    \I__1029\ : InMux
    port map (
            O => \N__6007\,
            I => \N__5961\
        );

    \I__1028\ : InMux
    port map (
            O => \N__6006\,
            I => \N__5961\
        );

    \I__1027\ : InMux
    port map (
            O => \N__6005\,
            I => \N__5954\
        );

    \I__1026\ : InMux
    port map (
            O => \N__6002\,
            I => \N__5954\
        );

    \I__1025\ : InMux
    port map (
            O => \N__6001\,
            I => \N__5954\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__5996\,
            I => \N__5951\
        );

    \I__1023\ : InMux
    port map (
            O => \N__5995\,
            I => \N__5948\
        );

    \I__1022\ : Odrv4
    port map (
            O => \N__5992\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1021\ : Odrv4
    port map (
            O => \N__5989\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__5986\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__5983\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1018\ : Odrv12
    port map (
            O => \N__5978\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__5975\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__5968\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__5961\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__5954\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1013\ : Odrv4
    port map (
            O => \N__5951\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__5948\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1011\ : InMux
    port map (
            O => \N__5925\,
            I => \N__5918\
        );

    \I__1010\ : InMux
    port map (
            O => \N__5924\,
            I => \N__5911\
        );

    \I__1009\ : InMux
    port map (
            O => \N__5923\,
            I => \N__5911\
        );

    \I__1008\ : InMux
    port map (
            O => \N__5922\,
            I => \N__5911\
        );

    \I__1007\ : InMux
    port map (
            O => \N__5921\,
            I => \N__5904\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__5918\,
            I => \N__5899\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__5911\,
            I => \N__5899\
        );

    \I__1004\ : InMux
    port map (
            O => \N__5910\,
            I => \N__5896\
        );

    \I__1003\ : InMux
    port map (
            O => \N__5909\,
            I => \N__5891\
        );

    \I__1002\ : InMux
    port map (
            O => \N__5908\,
            I => \N__5891\
        );

    \I__1001\ : InMux
    port map (
            O => \N__5907\,
            I => \N__5888\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__5904\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__999\ : Odrv4
    port map (
            O => \N__5899\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__5896\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__5891\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__5888\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__995\ : InMux
    port map (
            O => \N__5877\,
            I => \N__5867\
        );

    \I__994\ : InMux
    port map (
            O => \N__5876\,
            I => \N__5867\
        );

    \I__993\ : InMux
    port map (
            O => \N__5875\,
            I => \N__5864\
        );

    \I__992\ : InMux
    port map (
            O => \N__5874\,
            I => \N__5857\
        );

    \I__991\ : InMux
    port map (
            O => \N__5873\,
            I => \N__5851\
        );

    \I__990\ : InMux
    port map (
            O => \N__5872\,
            I => \N__5851\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__5867\,
            I => \N__5848\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__5864\,
            I => \N__5845\
        );

    \I__987\ : InMux
    port map (
            O => \N__5863\,
            I => \N__5840\
        );

    \I__986\ : InMux
    port map (
            O => \N__5862\,
            I => \N__5840\
        );

    \I__985\ : InMux
    port map (
            O => \N__5861\,
            I => \N__5835\
        );

    \I__984\ : InMux
    port map (
            O => \N__5860\,
            I => \N__5835\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__5857\,
            I => \N__5831\
        );

    \I__982\ : InMux
    port map (
            O => \N__5856\,
            I => \N__5828\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__5851\,
            I => \N__5819\
        );

    \I__980\ : Span4Mux_h
    port map (
            O => \N__5848\,
            I => \N__5819\
        );

    \I__979\ : Span4Mux_v
    port map (
            O => \N__5845\,
            I => \N__5819\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__5840\,
            I => \N__5819\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__5835\,
            I => \N__5816\
        );

    \I__976\ : InMux
    port map (
            O => \N__5834\,
            I => \N__5813\
        );

    \I__975\ : Span4Mux_h
    port map (
            O => \N__5831\,
            I => \N__5810\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__5828\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__973\ : Odrv4
    port map (
            O => \N__5819\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__972\ : Odrv4
    port map (
            O => \N__5816\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__5813\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__970\ : Odrv4
    port map (
            O => \N__5810\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__969\ : InMux
    port map (
            O => \N__5799\,
            I => \N__5794\
        );

    \I__968\ : InMux
    port map (
            O => \N__5798\,
            I => \N__5790\
        );

    \I__967\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5786\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__5794\,
            I => \N__5779\
        );

    \I__965\ : CascadeMux
    port map (
            O => \N__5793\,
            I => \N__5776\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__5790\,
            I => \N__5772\
        );

    \I__963\ : InMux
    port map (
            O => \N__5789\,
            I => \N__5769\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__5786\,
            I => \N__5766\
        );

    \I__961\ : CascadeMux
    port map (
            O => \N__5785\,
            I => \N__5763\
        );

    \I__960\ : CascadeMux
    port map (
            O => \N__5784\,
            I => \N__5757\
        );

    \I__959\ : InMux
    port map (
            O => \N__5783\,
            I => \N__5752\
        );

    \I__958\ : InMux
    port map (
            O => \N__5782\,
            I => \N__5752\
        );

    \I__957\ : Span4Mux_h
    port map (
            O => \N__5779\,
            I => \N__5747\
        );

    \I__956\ : InMux
    port map (
            O => \N__5776\,
            I => \N__5744\
        );

    \I__955\ : InMux
    port map (
            O => \N__5775\,
            I => \N__5741\
        );

    \I__954\ : Span4Mux_h
    port map (
            O => \N__5772\,
            I => \N__5734\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__5769\,
            I => \N__5734\
        );

    \I__952\ : Span4Mux_h
    port map (
            O => \N__5766\,
            I => \N__5734\
        );

    \I__951\ : InMux
    port map (
            O => \N__5763\,
            I => \N__5729\
        );

    \I__950\ : InMux
    port map (
            O => \N__5762\,
            I => \N__5729\
        );

    \I__949\ : InMux
    port map (
            O => \N__5761\,
            I => \N__5722\
        );

    \I__948\ : InMux
    port map (
            O => \N__5760\,
            I => \N__5722\
        );

    \I__947\ : InMux
    port map (
            O => \N__5757\,
            I => \N__5722\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__5752\,
            I => \N__5719\
        );

    \I__945\ : InMux
    port map (
            O => \N__5751\,
            I => \N__5714\
        );

    \I__944\ : InMux
    port map (
            O => \N__5750\,
            I => \N__5714\
        );

    \I__943\ : Odrv4
    port map (
            O => \N__5747\,
            I => \U712_CHIP_RAM.N_352\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__5744\,
            I => \U712_CHIP_RAM.N_352\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__5741\,
            I => \U712_CHIP_RAM.N_352\
        );

    \I__940\ : Odrv4
    port map (
            O => \N__5734\,
            I => \U712_CHIP_RAM.N_352\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__5729\,
            I => \U712_CHIP_RAM.N_352\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__5722\,
            I => \U712_CHIP_RAM.N_352\
        );

    \I__937\ : Odrv4
    port map (
            O => \N__5719\,
            I => \U712_CHIP_RAM.N_352\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__5714\,
            I => \U712_CHIP_RAM.N_352\
        );

    \I__935\ : CascadeMux
    port map (
            O => \N__5697\,
            I => \N__5693\
        );

    \I__934\ : InMux
    port map (
            O => \N__5696\,
            I => \N__5688\
        );

    \I__933\ : InMux
    port map (
            O => \N__5693\,
            I => \N__5685\
        );

    \I__932\ : InMux
    port map (
            O => \N__5692\,
            I => \N__5680\
        );

    \I__931\ : InMux
    port map (
            O => \N__5691\,
            I => \N__5677\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__5688\,
            I => \N__5672\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__5685\,
            I => \N__5672\
        );

    \I__928\ : CascadeMux
    port map (
            O => \N__5684\,
            I => \N__5667\
        );

    \I__927\ : InMux
    port map (
            O => \N__5683\,
            I => \N__5660\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__5680\,
            I => \N__5657\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__5677\,
            I => \N__5652\
        );

    \I__924\ : Span4Mux_v
    port map (
            O => \N__5672\,
            I => \N__5652\
        );

    \I__923\ : InMux
    port map (
            O => \N__5671\,
            I => \N__5643\
        );

    \I__922\ : InMux
    port map (
            O => \N__5670\,
            I => \N__5643\
        );

    \I__921\ : InMux
    port map (
            O => \N__5667\,
            I => \N__5643\
        );

    \I__920\ : InMux
    port map (
            O => \N__5666\,
            I => \N__5643\
        );

    \I__919\ : InMux
    port map (
            O => \N__5665\,
            I => \N__5638\
        );

    \I__918\ : InMux
    port map (
            O => \N__5664\,
            I => \N__5638\
        );

    \I__917\ : InMux
    port map (
            O => \N__5663\,
            I => \N__5635\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__5660\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__915\ : Odrv4
    port map (
            O => \N__5657\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__914\ : Odrv4
    port map (
            O => \N__5652\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__5643\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__5638\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__5635\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__910\ : InMux
    port map (
            O => \N__5622\,
            I => \N__5619\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__5619\,
            I => \N__5615\
        );

    \I__908\ : InMux
    port map (
            O => \N__5618\,
            I => \N__5612\
        );

    \I__907\ : Odrv4
    port map (
            O => \N__5615\,
            I => \U712_REG_SM.N_232\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__5612\,
            I => \U712_REG_SM.N_232\
        );

    \I__905\ : CascadeMux
    port map (
            O => \N__5607\,
            I => \N__5604\
        );

    \I__904\ : InMux
    port map (
            O => \N__5604\,
            I => \N__5600\
        );

    \I__903\ : InMux
    port map (
            O => \N__5603\,
            I => \N__5597\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__5600\,
            I => \REG_TACK\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__5597\,
            I => \REG_TACK\
        );

    \I__900\ : InMux
    port map (
            O => \N__5592\,
            I => \N__5589\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__5589\,
            I => \U712_REG_SM.N_289\
        );

    \I__898\ : InMux
    port map (
            O => \N__5586\,
            I => \N__5583\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__5583\,
            I => \N__5578\
        );

    \I__896\ : InMux
    port map (
            O => \N__5582\,
            I => \N__5567\
        );

    \I__895\ : InMux
    port map (
            O => \N__5581\,
            I => \N__5567\
        );

    \I__894\ : Span4Mux_h
    port map (
            O => \N__5578\,
            I => \N__5564\
        );

    \I__893\ : InMux
    port map (
            O => \N__5577\,
            I => \N__5561\
        );

    \I__892\ : InMux
    port map (
            O => \N__5576\,
            I => \N__5558\
        );

    \I__891\ : InMux
    port map (
            O => \N__5575\,
            I => \N__5555\
        );

    \I__890\ : InMux
    port map (
            O => \N__5574\,
            I => \N__5552\
        );

    \I__889\ : InMux
    port map (
            O => \N__5573\,
            I => \N__5547\
        );

    \I__888\ : InMux
    port map (
            O => \N__5572\,
            I => \N__5547\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__5567\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__886\ : Odrv4
    port map (
            O => \N__5564\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5561\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__5558\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__5555\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__5552\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__5547\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__880\ : InMux
    port map (
            O => \N__5532\,
            I => \N__5529\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__5529\,
            I => \N__5526\
        );

    \I__878\ : Odrv4
    port map (
            O => \N__5526\,
            I => \U712_REG_SM.N_254\
        );

    \I__877\ : CascadeMux
    port map (
            O => \N__5523\,
            I => \U712_REG_SM.N_254_cascade_\
        );

    \I__876\ : InMux
    port map (
            O => \N__5520\,
            I => \N__5517\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__5517\,
            I => \U712_REG_SM.N_26\
        );

    \I__874\ : InMux
    port map (
            O => \N__5514\,
            I => \N__5511\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__5511\,
            I => \N__5507\
        );

    \I__872\ : IoInMux
    port map (
            O => \N__5510\,
            I => \N__5504\
        );

    \I__871\ : Span4Mux_v
    port map (
            O => \N__5507\,
            I => \N__5501\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__5504\,
            I => \N__5498\
        );

    \I__869\ : Sp12to4
    port map (
            O => \N__5501\,
            I => \N__5495\
        );

    \I__868\ : IoSpan4Mux
    port map (
            O => \N__5498\,
            I => \N__5492\
        );

    \I__867\ : Span12Mux_h
    port map (
            O => \N__5495\,
            I => \N__5489\
        );

    \I__866\ : IoSpan4Mux
    port map (
            O => \N__5492\,
            I => \N__5486\
        );

    \I__865\ : Span12Mux_v
    port map (
            O => \N__5489\,
            I => \N__5483\
        );

    \I__864\ : IoSpan4Mux
    port map (
            O => \N__5486\,
            I => \N__5480\
        );

    \I__863\ : Odrv12
    port map (
            O => \N__5483\,
            I => \C1_c\
        );

    \I__862\ : Odrv4
    port map (
            O => \N__5480\,
            I => \C1_c\
        );

    \I__861\ : InMux
    port map (
            O => \N__5475\,
            I => \N__5472\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__5472\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__859\ : InMux
    port map (
            O => \N__5469\,
            I => \N__5466\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5466\,
            I => \N__5463\
        );

    \I__857\ : Span4Mux_h
    port map (
            O => \N__5463\,
            I => \N__5460\
        );

    \I__856\ : Odrv4
    port map (
            O => \N__5460\,
            I => \U712_CHIP_RAM.un3_DMA_CYCLE_START\
        );

    \I__855\ : InMux
    port map (
            O => \N__5457\,
            I => \N__5454\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__5454\,
            I => \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_0\
        );

    \I__853\ : InMux
    port map (
            O => \N__5451\,
            I => \N__5448\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__5448\,
            I => \N__5444\
        );

    \I__851\ : InMux
    port map (
            O => \N__5447\,
            I => \N__5439\
        );

    \I__850\ : Span4Mux_h
    port map (
            O => \N__5444\,
            I => \N__5436\
        );

    \I__849\ : InMux
    port map (
            O => \N__5443\,
            I => \N__5433\
        );

    \I__848\ : InMux
    port map (
            O => \N__5442\,
            I => \N__5430\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__5439\,
            I => \U712_CHIP_RAM.N_207\
        );

    \I__846\ : Odrv4
    port map (
            O => \N__5436\,
            I => \U712_CHIP_RAM.N_207\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__5433\,
            I => \U712_CHIP_RAM.N_207\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__5430\,
            I => \U712_CHIP_RAM.N_207\
        );

    \I__843\ : InMux
    port map (
            O => \N__5421\,
            I => \N__5418\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__5418\,
            I => \N__5415\
        );

    \I__841\ : Odrv4
    port map (
            O => \N__5415\,
            I => \U712_CHIP_RAM.CLK_EN_5_0_a2_1_a2_0\
        );

    \I__840\ : InMux
    port map (
            O => \N__5412\,
            I => \N__5409\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__5409\,
            I => \N__5406\
        );

    \I__838\ : Span4Mux_h
    port map (
            O => \N__5406\,
            I => \N__5403\
        );

    \I__837\ : Odrv4
    port map (
            O => \N__5403\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0_1\
        );

    \I__836\ : InMux
    port map (
            O => \N__5400\,
            I => \N__5393\
        );

    \I__835\ : CascadeMux
    port map (
            O => \N__5399\,
            I => \N__5388\
        );

    \I__834\ : InMux
    port map (
            O => \N__5398\,
            I => \N__5385\
        );

    \I__833\ : InMux
    port map (
            O => \N__5397\,
            I => \N__5379\
        );

    \I__832\ : InMux
    port map (
            O => \N__5396\,
            I => \N__5379\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__5393\,
            I => \N__5376\
        );

    \I__830\ : InMux
    port map (
            O => \N__5392\,
            I => \N__5370\
        );

    \I__829\ : InMux
    port map (
            O => \N__5391\,
            I => \N__5370\
        );

    \I__828\ : InMux
    port map (
            O => \N__5388\,
            I => \N__5367\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__5385\,
            I => \N__5364\
        );

    \I__826\ : InMux
    port map (
            O => \N__5384\,
            I => \N__5361\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__5379\,
            I => \N__5358\
        );

    \I__824\ : Span4Mux_h
    port map (
            O => \N__5376\,
            I => \N__5355\
        );

    \I__823\ : InMux
    port map (
            O => \N__5375\,
            I => \N__5352\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__5370\,
            I => \N__5349\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__5367\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__820\ : Odrv4
    port map (
            O => \N__5364\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__5361\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__818\ : Odrv4
    port map (
            O => \N__5358\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__817\ : Odrv4
    port map (
            O => \N__5355\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__5352\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__815\ : Odrv4
    port map (
            O => \N__5349\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__814\ : CascadeMux
    port map (
            O => \N__5334\,
            I => \N__5328\
        );

    \I__813\ : CascadeMux
    port map (
            O => \N__5333\,
            I => \N__5324\
        );

    \I__812\ : CascadeMux
    port map (
            O => \N__5332\,
            I => \N__5321\
        );

    \I__811\ : CascadeMux
    port map (
            O => \N__5331\,
            I => \N__5318\
        );

    \I__810\ : InMux
    port map (
            O => \N__5328\,
            I => \N__5315\
        );

    \I__809\ : InMux
    port map (
            O => \N__5327\,
            I => \N__5312\
        );

    \I__808\ : InMux
    port map (
            O => \N__5324\,
            I => \N__5307\
        );

    \I__807\ : InMux
    port map (
            O => \N__5321\,
            I => \N__5307\
        );

    \I__806\ : InMux
    port map (
            O => \N__5318\,
            I => \N__5304\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__5315\,
            I => \N__5297\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__5312\,
            I => \N__5297\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__5307\,
            I => \N__5297\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__5304\,
            I => \N__5294\
        );

    \I__801\ : Span4Mux_h
    port map (
            O => \N__5297\,
            I => \N__5291\
        );

    \I__800\ : Odrv4
    port map (
            O => \N__5294\,
            I => \U712_CHIP_RAM.N_370\
        );

    \I__799\ : Odrv4
    port map (
            O => \N__5291\,
            I => \U712_CHIP_RAM.N_370\
        );

    \I__798\ : InMux
    port map (
            O => \N__5286\,
            I => \N__5283\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5283\,
            I => \U712_CHIP_RAM.N_307\
        );

    \I__796\ : InMux
    port map (
            O => \N__5280\,
            I => \N__5277\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__5277\,
            I => \N__5273\
        );

    \I__794\ : InMux
    port map (
            O => \N__5276\,
            I => \N__5270\
        );

    \I__793\ : Span4Mux_h
    port map (
            O => \N__5273\,
            I => \N__5267\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__5270\,
            I => \U712_CHIP_RAM.N_411\
        );

    \I__791\ : Odrv4
    port map (
            O => \N__5267\,
            I => \U712_CHIP_RAM.N_411\
        );

    \I__790\ : InMux
    port map (
            O => \N__5262\,
            I => \N__5257\
        );

    \I__789\ : InMux
    port map (
            O => \N__5261\,
            I => \N__5254\
        );

    \I__788\ : InMux
    port map (
            O => \N__5260\,
            I => \N__5251\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5257\,
            I => \N__5248\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__5254\,
            I => \N__5245\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__5251\,
            I => \U712_CHIP_RAM.N_403\
        );

    \I__784\ : Odrv4
    port map (
            O => \N__5248\,
            I => \U712_CHIP_RAM.N_403\
        );

    \I__783\ : Odrv4
    port map (
            O => \N__5245\,
            I => \U712_CHIP_RAM.N_403\
        );

    \I__782\ : CascadeMux
    port map (
            O => \N__5238\,
            I => \U712_CHIP_RAM.N_411_cascade_\
        );

    \I__781\ : InMux
    port map (
            O => \N__5235\,
            I => \N__5232\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__5232\,
            I => \U712_CHIP_RAM.N_308\
        );

    \I__779\ : InMux
    port map (
            O => \N__5229\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__778\ : InMux
    port map (
            O => \N__5226\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__777\ : InMux
    port map (
            O => \N__5223\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__776\ : InMux
    port map (
            O => \N__5220\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__775\ : InMux
    port map (
            O => \N__5217\,
            I => \N__5208\
        );

    \I__774\ : InMux
    port map (
            O => \N__5216\,
            I => \N__5201\
        );

    \I__773\ : InMux
    port map (
            O => \N__5215\,
            I => \N__5201\
        );

    \I__772\ : InMux
    port map (
            O => \N__5214\,
            I => \N__5201\
        );

    \I__771\ : InMux
    port map (
            O => \N__5213\,
            I => \N__5194\
        );

    \I__770\ : InMux
    port map (
            O => \N__5212\,
            I => \N__5194\
        );

    \I__769\ : InMux
    port map (
            O => \N__5211\,
            I => \N__5194\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__5208\,
            I => \U712_CHIP_RAM.N_49\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__5201\,
            I => \U712_CHIP_RAM.N_49\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__5194\,
            I => \U712_CHIP_RAM.N_49\
        );

    \I__765\ : InMux
    port map (
            O => \N__5187\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__764\ : CEMux
    port map (
            O => \N__5184\,
            I => \N__5181\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__5181\,
            I => \N__5177\
        );

    \I__762\ : CEMux
    port map (
            O => \N__5180\,
            I => \N__5173\
        );

    \I__761\ : Span4Mux_h
    port map (
            O => \N__5177\,
            I => \N__5170\
        );

    \I__760\ : CEMux
    port map (
            O => \N__5176\,
            I => \N__5167\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__5173\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__758\ : Odrv4
    port map (
            O => \N__5170\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__5167\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__756\ : InMux
    port map (
            O => \N__5160\,
            I => \N__5156\
        );

    \I__755\ : InMux
    port map (
            O => \N__5159\,
            I => \N__5153\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__5156\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__5153\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__752\ : InMux
    port map (
            O => \N__5148\,
            I => \N__5144\
        );

    \I__751\ : InMux
    port map (
            O => \N__5147\,
            I => \N__5141\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__5144\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__5141\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__748\ : CascadeMux
    port map (
            O => \N__5136\,
            I => \N__5133\
        );

    \I__747\ : InMux
    port map (
            O => \N__5133\,
            I => \N__5129\
        );

    \I__746\ : InMux
    port map (
            O => \N__5132\,
            I => \N__5126\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__5129\,
            I => \N__5123\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__5126\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__743\ : Odrv4
    port map (
            O => \N__5123\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__742\ : InMux
    port map (
            O => \N__5118\,
            I => \N__5114\
        );

    \I__741\ : InMux
    port map (
            O => \N__5117\,
            I => \N__5111\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__5114\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__5111\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__738\ : CascadeMux
    port map (
            O => \N__5106\,
            I => \U712_CHIP_RAM.N_352_cascade_\
        );

    \I__737\ : CascadeMux
    port map (
            O => \N__5103\,
            I => \U712_CHIP_RAM.N_328_cascade_\
        );

    \I__736\ : InMux
    port map (
            O => \N__5100\,
            I => \N__5097\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__5097\,
            I => \U712_CHIP_RAM.N_323\
        );

    \I__734\ : InMux
    port map (
            O => \N__5094\,
            I => \N__5091\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__5091\,
            I => \U712_CHIP_RAM.N_63\
        );

    \I__732\ : IoInMux
    port map (
            O => \N__5088\,
            I => \N__5085\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__5085\,
            I => \N__5082\
        );

    \I__730\ : IoSpan4Mux
    port map (
            O => \N__5082\,
            I => \N__5079\
        );

    \I__729\ : Span4Mux_s3_v
    port map (
            O => \N__5079\,
            I => \N__5076\
        );

    \I__728\ : Sp12to4
    port map (
            O => \N__5076\,
            I => \N__5073\
        );

    \I__727\ : Span12Mux_s10_v
    port map (
            O => \N__5073\,
            I => \N__5070\
        );

    \I__726\ : Span12Mux_v
    port map (
            O => \N__5070\,
            I => \N__5066\
        );

    \I__725\ : InMux
    port map (
            O => \N__5069\,
            I => \N__5063\
        );

    \I__724\ : Odrv12
    port map (
            O => \N__5066\,
            I => \LATCH_CLK_c\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__5063\,
            I => \LATCH_CLK_c\
        );

    \I__722\ : InMux
    port map (
            O => \N__5058\,
            I => \N__5052\
        );

    \I__721\ : InMux
    port map (
            O => \N__5057\,
            I => \N__5049\
        );

    \I__720\ : InMux
    port map (
            O => \N__5056\,
            I => \N__5046\
        );

    \I__719\ : InMux
    port map (
            O => \N__5055\,
            I => \N__5043\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__5052\,
            I => \N__5040\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__5049\,
            I => \N__5033\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__5046\,
            I => \N__5033\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__5043\,
            I => \N__5033\
        );

    \I__714\ : Span4Mux_h
    port map (
            O => \N__5040\,
            I => \N__5026\
        );

    \I__713\ : Span4Mux_v
    port map (
            O => \N__5033\,
            I => \N__5026\
        );

    \I__712\ : InMux
    port map (
            O => \N__5032\,
            I => \N__5021\
        );

    \I__711\ : InMux
    port map (
            O => \N__5031\,
            I => \N__5021\
        );

    \I__710\ : Odrv4
    port map (
            O => \N__5026\,
            I => \U712_CHIP_RAM.N_363\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__5021\,
            I => \U712_CHIP_RAM.N_363\
        );

    \I__708\ : CascadeMux
    port map (
            O => \N__5016\,
            I => \U712_CHIP_RAM.N_363_cascade_\
        );

    \I__707\ : InMux
    port map (
            O => \N__5013\,
            I => \N__5010\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__5010\,
            I => \U712_CHIP_RAM.N_369\
        );

    \I__705\ : InMux
    port map (
            O => \N__5007\,
            I => \N__5001\
        );

    \I__704\ : InMux
    port map (
            O => \N__5006\,
            I => \N__4996\
        );

    \I__703\ : InMux
    port map (
            O => \N__5005\,
            I => \N__4996\
        );

    \I__702\ : InMux
    port map (
            O => \N__5004\,
            I => \N__4993\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__5001\,
            I => \U712_CHIP_RAM.N_397\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__4996\,
            I => \U712_CHIP_RAM.N_397\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__4993\,
            I => \U712_CHIP_RAM.N_397\
        );

    \I__698\ : InMux
    port map (
            O => \N__4986\,
            I => \N__4983\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__4983\,
            I => \N__4979\
        );

    \I__696\ : InMux
    port map (
            O => \N__4982\,
            I => \N__4976\
        );

    \I__695\ : Odrv4
    port map (
            O => \N__4979\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__4976\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0\
        );

    \I__693\ : InMux
    port map (
            O => \N__4971\,
            I => \N__4968\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__4968\,
            I => \N__4965\
        );

    \I__691\ : Odrv4
    port map (
            O => \N__4965\,
            I => \U712_CHIP_RAM.N_306\
        );

    \I__690\ : InMux
    port map (
            O => \N__4962\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__689\ : InMux
    port map (
            O => \N__4959\,
            I => \N__4956\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__4956\,
            I => \N__4953\
        );

    \I__687\ : Odrv4
    port map (
            O => \N__4953\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__686\ : InMux
    port map (
            O => \N__4950\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__685\ : CascadeMux
    port map (
            O => \N__4947\,
            I => \N__4944\
        );

    \I__684\ : InMux
    port map (
            O => \N__4944\,
            I => \N__4940\
        );

    \I__683\ : InMux
    port map (
            O => \N__4943\,
            I => \N__4937\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__4940\,
            I => \U712_REG_SM.N_255\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__4937\,
            I => \U712_REG_SM.N_255\
        );

    \I__680\ : IoInMux
    port map (
            O => \N__4932\,
            I => \N__4929\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__4929\,
            I => \N__4926\
        );

    \I__678\ : IoSpan4Mux
    port map (
            O => \N__4926\,
            I => \N__4923\
        );

    \I__677\ : Span4Mux_s3_h
    port map (
            O => \N__4923\,
            I => \N__4920\
        );

    \I__676\ : Span4Mux_h
    port map (
            O => \N__4920\,
            I => \N__4917\
        );

    \I__675\ : Sp12to4
    port map (
            O => \N__4917\,
            I => \N__4913\
        );

    \I__674\ : InMux
    port map (
            O => \N__4916\,
            I => \N__4910\
        );

    \I__673\ : Span12Mux_h
    port map (
            O => \N__4913\,
            I => \N__4905\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__4910\,
            I => \N__4905\
        );

    \I__671\ : Span12Mux_h
    port map (
            O => \N__4905\,
            I => \N__4902\
        );

    \I__670\ : Span12Mux_v
    port map (
            O => \N__4902\,
            I => \N__4899\
        );

    \I__669\ : Odrv12
    port map (
            O => \N__4899\,
            I => \C3_c\
        );

    \I__668\ : InMux
    port map (
            O => \N__4896\,
            I => \N__4893\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__4893\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__666\ : CascadeMux
    port map (
            O => \N__4890\,
            I => \N__4887\
        );

    \I__665\ : InMux
    port map (
            O => \N__4887\,
            I => \N__4884\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__4884\,
            I => \U712_REG_SM.STATE_COUNT_srsts_i_0_a2_0_0_0\
        );

    \I__663\ : InMux
    port map (
            O => \N__4881\,
            I => \N__4877\
        );

    \I__662\ : InMux
    port map (
            O => \N__4880\,
            I => \N__4872\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__4877\,
            I => \N__4869\
        );

    \I__660\ : InMux
    port map (
            O => \N__4876\,
            I => \N__4864\
        );

    \I__659\ : InMux
    port map (
            O => \N__4875\,
            I => \N__4864\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__4872\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__657\ : Odrv4
    port map (
            O => \N__4869\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__4864\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__655\ : InMux
    port map (
            O => \N__4857\,
            I => \N__4854\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__4854\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__653\ : InMux
    port map (
            O => \N__4851\,
            I => \N__4846\
        );

    \I__652\ : InMux
    port map (
            O => \N__4850\,
            I => \N__4841\
        );

    \I__651\ : InMux
    port map (
            O => \N__4849\,
            I => \N__4841\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__4846\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__4841\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__648\ : InMux
    port map (
            O => \N__4836\,
            I => \N__4833\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__4833\,
            I => \U712_REG_SM.N_264\
        );

    \I__646\ : InMux
    port map (
            O => \N__4830\,
            I => \N__4827\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__4827\,
            I => \U712_REG_SM.N_24\
        );

    \I__644\ : CascadeMux
    port map (
            O => \N__4824\,
            I => \N__4821\
        );

    \I__643\ : InMux
    port map (
            O => \N__4821\,
            I => \N__4817\
        );

    \I__642\ : CascadeMux
    port map (
            O => \N__4820\,
            I => \N__4814\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__4817\,
            I => \N__4808\
        );

    \I__640\ : InMux
    port map (
            O => \N__4814\,
            I => \N__4805\
        );

    \I__639\ : InMux
    port map (
            O => \N__4813\,
            I => \N__4802\
        );

    \I__638\ : InMux
    port map (
            O => \N__4812\,
            I => \N__4799\
        );

    \I__637\ : InMux
    port map (
            O => \N__4811\,
            I => \N__4796\
        );

    \I__636\ : Odrv4
    port map (
            O => \N__4808\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__4805\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__4802\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__4799\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__4796\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__631\ : InMux
    port map (
            O => \N__4785\,
            I => \N__4782\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__4782\,
            I => \U712_CHIP_RAM.N_262\
        );

    \I__629\ : CascadeMux
    port map (
            O => \N__4779\,
            I => \U712_CHIP_RAM.N_354_cascade_\
        );

    \I__628\ : InMux
    port map (
            O => \N__4776\,
            I => \N__4773\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__4773\,
            I => \U712_CHIP_RAM.N_408\
        );

    \I__626\ : CascadeMux
    port map (
            O => \N__4770\,
            I => \U712_CHIP_RAM.N_408_cascade_\
        );

    \I__625\ : InMux
    port map (
            O => \N__4767\,
            I => \N__4764\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__4764\,
            I => \N__4759\
        );

    \I__623\ : InMux
    port map (
            O => \N__4763\,
            I => \N__4756\
        );

    \I__622\ : InMux
    port map (
            O => \N__4762\,
            I => \N__4753\
        );

    \I__621\ : Odrv12
    port map (
            O => \N__4759\,
            I => \U712_CHIP_RAM.N_359\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__4756\,
            I => \U712_CHIP_RAM.N_359\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__4753\,
            I => \U712_CHIP_RAM.N_359\
        );

    \I__618\ : InMux
    port map (
            O => \N__4746\,
            I => \N__4740\
        );

    \I__617\ : InMux
    port map (
            O => \N__4745\,
            I => \N__4740\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__4740\,
            I => \U712_CHIP_RAM.N_305\
        );

    \I__615\ : CascadeMux
    port map (
            O => \N__4737\,
            I => \U712_CYCLE_TERM.N_236_i_0_en_cascade_\
        );

    \I__614\ : CEMux
    port map (
            O => \N__4734\,
            I => \N__4731\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__4731\,
            I => \U712_CYCLE_TERM.N_236_i_0_en_0\
        );

    \I__612\ : InMux
    port map (
            O => \N__4728\,
            I => \N__4725\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__4725\,
            I => \U712_REG_SM.STATE_COUNTc_1_0\
        );

    \I__610\ : CascadeMux
    port map (
            O => \N__4722\,
            I => \N__4719\
        );

    \I__609\ : InMux
    port map (
            O => \N__4719\,
            I => \N__4714\
        );

    \I__608\ : InMux
    port map (
            O => \N__4718\,
            I => \N__4711\
        );

    \I__607\ : InMux
    port map (
            O => \N__4717\,
            I => \N__4708\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__4714\,
            I => \N__4705\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__4711\,
            I => \N__4702\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__4708\,
            I => \N__4699\
        );

    \I__603\ : Span4Mux_v
    port map (
            O => \N__4705\,
            I => \N__4694\
        );

    \I__602\ : Span4Mux_h
    port map (
            O => \N__4702\,
            I => \N__4689\
        );

    \I__601\ : Span4Mux_h
    port map (
            O => \N__4699\,
            I => \N__4689\
        );

    \I__600\ : InMux
    port map (
            O => \N__4698\,
            I => \N__4684\
        );

    \I__599\ : InMux
    port map (
            O => \N__4697\,
            I => \N__4684\
        );

    \I__598\ : Odrv4
    port map (
            O => \N__4694\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__597\ : Odrv4
    port map (
            O => \N__4689\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__4684\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__595\ : InMux
    port map (
            O => \N__4677\,
            I => \N__4674\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__4674\,
            I => \N__4671\
        );

    \I__593\ : Span4Mux_v
    port map (
            O => \N__4671\,
            I => \N__4668\
        );

    \I__592\ : Span4Mux_v
    port map (
            O => \N__4668\,
            I => \N__4665\
        );

    \I__591\ : Sp12to4
    port map (
            O => \N__4665\,
            I => \N__4662\
        );

    \I__590\ : Odrv12
    port map (
            O => \N__4662\,
            I => \A_c_15\
        );

    \I__589\ : InMux
    port map (
            O => \N__4659\,
            I => \N__4656\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__4656\,
            I => \N__4653\
        );

    \I__587\ : Span4Mux_v
    port map (
            O => \N__4653\,
            I => \N__4650\
        );

    \I__586\ : Span4Mux_h
    port map (
            O => \N__4650\,
            I => \N__4647\
        );

    \I__585\ : Sp12to4
    port map (
            O => \N__4647\,
            I => \N__4644\
        );

    \I__584\ : Odrv12
    port map (
            O => \N__4644\,
            I => \A_c_8\
        );

    \I__583\ : InMux
    port map (
            O => \N__4641\,
            I => \N__4638\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__4638\,
            I => \N__4635\
        );

    \I__581\ : Odrv4
    port map (
            O => \N__4635\,
            I => \U712_CHIP_RAM.N_217\
        );

    \I__580\ : InMux
    port map (
            O => \N__4632\,
            I => \N__4629\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__4629\,
            I => \U712_CHIP_RAM.N_361\
        );

    \I__578\ : CascadeMux
    port map (
            O => \N__4626\,
            I => \U712_CHIP_RAM.N_217_cascade_\
        );

    \I__577\ : CascadeMux
    port map (
            O => \N__4623\,
            I => \N__4619\
        );

    \I__576\ : InMux
    port map (
            O => \N__4622\,
            I => \N__4616\
        );

    \I__575\ : InMux
    port map (
            O => \N__4619\,
            I => \N__4613\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__4616\,
            I => \U712_CHIP_RAM.N_222\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__4613\,
            I => \U712_CHIP_RAM.N_222\
        );

    \I__572\ : CascadeMux
    port map (
            O => \N__4608\,
            I => \N__4602\
        );

    \I__571\ : InMux
    port map (
            O => \N__4607\,
            I => \N__4599\
        );

    \I__570\ : InMux
    port map (
            O => \N__4606\,
            I => \N__4592\
        );

    \I__569\ : InMux
    port map (
            O => \N__4605\,
            I => \N__4592\
        );

    \I__568\ : InMux
    port map (
            O => \N__4602\,
            I => \N__4592\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__4599\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__4592\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__565\ : CascadeMux
    port map (
            O => \N__4587\,
            I => \U712_CHIP_RAM.N_359_cascade_\
        );

    \I__564\ : InMux
    port map (
            O => \N__4584\,
            I => \N__4580\
        );

    \I__563\ : CascadeMux
    port map (
            O => \N__4583\,
            I => \N__4577\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__4580\,
            I => \N__4574\
        );

    \I__561\ : InMux
    port map (
            O => \N__4577\,
            I => \N__4569\
        );

    \I__560\ : Span4Mux_h
    port map (
            O => \N__4574\,
            I => \N__4566\
        );

    \I__559\ : InMux
    port map (
            O => \N__4573\,
            I => \N__4561\
        );

    \I__558\ : InMux
    port map (
            O => \N__4572\,
            I => \N__4561\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__4569\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__556\ : Odrv4
    port map (
            O => \N__4566\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__4561\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__554\ : CascadeMux
    port map (
            O => \N__4554\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_\
        );

    \I__553\ : CascadeMux
    port map (
            O => \N__4551\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_\
        );

    \I__552\ : InMux
    port map (
            O => \N__4548\,
            I => \N__4545\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__4545\,
            I => \N__4542\
        );

    \I__550\ : Sp12to4
    port map (
            O => \N__4542\,
            I => \N__4539\
        );

    \I__549\ : Span12Mux_v
    port map (
            O => \N__4539\,
            I => \N__4536\
        );

    \I__548\ : Span12Mux_h
    port map (
            O => \N__4536\,
            I => \N__4533\
        );

    \I__547\ : Odrv12
    port map (
            O => \N__4533\,
            I => \A_c_20\
        );

    \I__546\ : CascadeMux
    port map (
            O => \N__4530\,
            I => \N__4527\
        );

    \I__545\ : InMux
    port map (
            O => \N__4527\,
            I => \N__4523\
        );

    \I__544\ : InMux
    port map (
            O => \N__4526\,
            I => \N__4519\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__4523\,
            I => \N__4516\
        );

    \I__542\ : InMux
    port map (
            O => \N__4522\,
            I => \N__4511\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__4519\,
            I => \N__4506\
        );

    \I__540\ : Span4Mux_v
    port map (
            O => \N__4516\,
            I => \N__4506\
        );

    \I__539\ : InMux
    port map (
            O => \N__4515\,
            I => \N__4503\
        );

    \I__538\ : InMux
    port map (
            O => \N__4514\,
            I => \N__4500\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__4511\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__536\ : Odrv4
    port map (
            O => \N__4506\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__4503\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__4500\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__533\ : CascadeMux
    port map (
            O => \N__4491\,
            I => \U712_CHIP_RAM.N_330_cascade_\
        );

    \I__532\ : InMux
    port map (
            O => \N__4488\,
            I => \N__4485\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__4485\,
            I => \N__4482\
        );

    \I__530\ : Odrv4
    port map (
            O => \N__4482\,
            I => \U712_CHIP_RAM.N_331\
        );

    \I__529\ : CascadeMux
    port map (
            O => \N__4479\,
            I => \U712_CHIP_RAM.BANK0_9_cascade_\
        );

    \I__528\ : CascadeMux
    port map (
            O => \N__4476\,
            I => \N__4472\
        );

    \I__527\ : InMux
    port map (
            O => \N__4475\,
            I => \N__4469\
        );

    \I__526\ : InMux
    port map (
            O => \N__4472\,
            I => \N__4466\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__4469\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__4466\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__523\ : IoInMux
    port map (
            O => \N__4461\,
            I => \N__4458\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__4458\,
            I => \N__4455\
        );

    \I__521\ : Span4Mux_s3_v
    port map (
            O => \N__4455\,
            I => \N__4452\
        );

    \I__520\ : Span4Mux_v
    port map (
            O => \N__4452\,
            I => \N__4449\
        );

    \I__519\ : Span4Mux_v
    port map (
            O => \N__4449\,
            I => \N__4445\
        );

    \I__518\ : InMux
    port map (
            O => \N__4448\,
            I => \N__4442\
        );

    \I__517\ : Odrv4
    port map (
            O => \N__4445\,
            I => \BANK0_c\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__4442\,
            I => \BANK0_c\
        );

    \I__515\ : InMux
    port map (
            O => \N__4437\,
            I => \N__4434\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__4434\,
            I => \N__4431\
        );

    \I__513\ : Odrv4
    port map (
            O => \N__4431\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_0\
        );

    \I__512\ : InMux
    port map (
            O => \N__4428\,
            I => \N__4425\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__4425\,
            I => \U712_CHIP_RAM.N_16\
        );

    \I__510\ : CascadeMux
    port map (
            O => \N__4422\,
            I => \U712_CHIP_RAM.N_49_cascade_\
        );

    \I__509\ : InMux
    port map (
            O => \N__4419\,
            I => \N__4416\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__4416\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_55_i_a2_0_a2_0_0\
        );

    \I__507\ : InMux
    port map (
            O => \N__4413\,
            I => \N__4410\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__4410\,
            I => \N__4406\
        );

    \I__505\ : InMux
    port map (
            O => \N__4409\,
            I => \N__4403\
        );

    \I__504\ : Span4Mux_v
    port map (
            O => \N__4406\,
            I => \N__4398\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4403\,
            I => \N__4395\
        );

    \I__502\ : InMux
    port map (
            O => \N__4402\,
            I => \N__4392\
        );

    \I__501\ : InMux
    port map (
            O => \N__4401\,
            I => \N__4389\
        );

    \I__500\ : Odrv4
    port map (
            O => \N__4398\,
            I => \REG_CYCLEm\
        );

    \I__499\ : Odrv4
    port map (
            O => \N__4395\,
            I => \REG_CYCLEm\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__4392\,
            I => \REG_CYCLEm\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__4389\,
            I => \REG_CYCLEm\
        );

    \I__496\ : IoInMux
    port map (
            O => \N__4380\,
            I => \N__4376\
        );

    \I__495\ : IoInMux
    port map (
            O => \N__4379\,
            I => \N__4373\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__4376\,
            I => \N__4370\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__4373\,
            I => \N__4367\
        );

    \I__492\ : Sp12to4
    port map (
            O => \N__4370\,
            I => \N__4364\
        );

    \I__491\ : IoSpan4Mux
    port map (
            O => \N__4367\,
            I => \N__4361\
        );

    \I__490\ : Span12Mux_v
    port map (
            O => \N__4364\,
            I => \N__4358\
        );

    \I__489\ : Sp12to4
    port map (
            O => \N__4361\,
            I => \N__4355\
        );

    \I__488\ : Span12Mux_h
    port map (
            O => \N__4358\,
            I => \N__4350\
        );

    \I__487\ : Span12Mux_v
    port map (
            O => \N__4355\,
            I => \N__4350\
        );

    \I__486\ : Odrv12
    port map (
            O => \N__4350\,
            I => \DRDENn_c\
        );

    \I__485\ : CascadeMux
    port map (
            O => \N__4347\,
            I => \U712_CHIP_RAM.LATCH_CLK_8_i_0_0_cascade_\
        );

    \I__484\ : CascadeMux
    port map (
            O => \N__4344\,
            I => \U712_CHIP_RAM.N_368_cascade_\
        );

    \I__483\ : CascadeMux
    port map (
            O => \N__4341\,
            I => \U712_CHIP_RAM.N_323_cascade_\
        );

    \I__482\ : CascadeMux
    port map (
            O => \N__4338\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0_cascade_\
        );

    \I__481\ : InMux
    port map (
            O => \N__4335\,
            I => \N__4332\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__4332\,
            I => \N__4329\
        );

    \I__479\ : Span4Mux_v
    port map (
            O => \N__4329\,
            I => \N__4326\
        );

    \I__478\ : Sp12to4
    port map (
            O => \N__4326\,
            I => \N__4323\
        );

    \I__477\ : Span12Mux_h
    port map (
            O => \N__4323\,
            I => \N__4320\
        );

    \I__476\ : Odrv12
    port map (
            O => \N__4320\,
            I => \A_c_12\
        );

    \I__475\ : InMux
    port map (
            O => \N__4317\,
            I => \N__4314\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__4314\,
            I => \N__4311\
        );

    \I__473\ : Span12Mux_v
    port map (
            O => \N__4311\,
            I => \N__4308\
        );

    \I__472\ : Odrv12
    port map (
            O => \N__4308\,
            I => \A_c_5\
        );

    \I__471\ : InMux
    port map (
            O => \N__4305\,
            I => \N__4302\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__4302\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__469\ : InMux
    port map (
            O => \N__4299\,
            I => \N__4295\
        );

    \I__468\ : InMux
    port map (
            O => \N__4298\,
            I => \N__4292\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__4295\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__4292\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__465\ : InMux
    port map (
            O => \N__4287\,
            I => \N__4284\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__4284\,
            I => \TACK_EN_i_ess\
        );

    \I__463\ : CascadeMux
    port map (
            O => \N__4281\,
            I => \U712_REG_SM.N_294_cascade_\
        );

    \I__462\ : InMux
    port map (
            O => \N__4278\,
            I => \N__4275\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__4275\,
            I => \N__4271\
        );

    \I__460\ : InMux
    port map (
            O => \N__4274\,
            I => \N__4268\
        );

    \I__459\ : Span4Mux_v
    port map (
            O => \N__4271\,
            I => \N__4265\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__4268\,
            I => \N__4262\
        );

    \I__457\ : Sp12to4
    port map (
            O => \N__4265\,
            I => \N__4259\
        );

    \I__456\ : Span12Mux_h
    port map (
            O => \N__4262\,
            I => \N__4256\
        );

    \I__455\ : Span12Mux_h
    port map (
            O => \N__4259\,
            I => \N__4253\
        );

    \I__454\ : Span12Mux_v
    port map (
            O => \N__4256\,
            I => \N__4250\
        );

    \I__453\ : Span12Mux_v
    port map (
            O => \N__4253\,
            I => \N__4247\
        );

    \I__452\ : Odrv12
    port map (
            O => \N__4250\,
            I => \TSn_c\
        );

    \I__451\ : Odrv12
    port map (
            O => \N__4247\,
            I => \TSn_c\
        );

    \I__450\ : CascadeMux
    port map (
            O => \N__4242\,
            I => \N__4239\
        );

    \I__449\ : InMux
    port map (
            O => \N__4239\,
            I => \N__4236\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__4236\,
            I => \N__4233\
        );

    \I__447\ : Span4Mux_v
    port map (
            O => \N__4233\,
            I => \N__4230\
        );

    \I__446\ : Sp12to4
    port map (
            O => \N__4230\,
            I => \N__4227\
        );

    \I__445\ : Span12Mux_h
    port map (
            O => \N__4227\,
            I => \N__4224\
        );

    \I__444\ : Span12Mux_v
    port map (
            O => \N__4224\,
            I => \N__4221\
        );

    \I__443\ : Odrv12
    port map (
            O => \N__4221\,
            I => \REGSPACEn_c\
        );

    \I__442\ : InMux
    port map (
            O => \N__4218\,
            I => \N__4214\
        );

    \I__441\ : InMux
    port map (
            O => \N__4217\,
            I => \N__4211\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__4214\,
            I => \N__4206\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__4211\,
            I => \N__4206\
        );

    \I__438\ : Span12Mux_h
    port map (
            O => \N__4206\,
            I => \N__4203\
        );

    \I__437\ : Span12Mux_v
    port map (
            O => \N__4203\,
            I => \N__4200\
        );

    \I__436\ : Odrv12
    port map (
            O => \N__4200\,
            I => \AWEn_c\
        );

    \I__435\ : InMux
    port map (
            O => \N__4197\,
            I => \N__4192\
        );

    \I__434\ : InMux
    port map (
            O => \N__4196\,
            I => \N__4187\
        );

    \I__433\ : InMux
    port map (
            O => \N__4195\,
            I => \N__4187\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__4192\,
            I => \U712_CHIP_RAM.N_371\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__4187\,
            I => \U712_CHIP_RAM.N_371\
        );

    \I__430\ : IoInMux
    port map (
            O => \N__4182\,
            I => \N__4179\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__4179\,
            I => \N__4176\
        );

    \I__428\ : IoSpan4Mux
    port map (
            O => \N__4176\,
            I => \N__4173\
        );

    \I__427\ : Span4Mux_s2_v
    port map (
            O => \N__4173\,
            I => \N__4169\
        );

    \I__426\ : CascadeMux
    port map (
            O => \N__4172\,
            I => \N__4166\
        );

    \I__425\ : Sp12to4
    port map (
            O => \N__4169\,
            I => \N__4163\
        );

    \I__424\ : InMux
    port map (
            O => \N__4166\,
            I => \N__4160\
        );

    \I__423\ : Odrv12
    port map (
            O => \N__4163\,
            I => \DBDIR_c\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__4160\,
            I => \DBDIR_c\
        );

    \I__421\ : CascadeMux
    port map (
            O => \N__4155\,
            I => \U712_CHIP_RAM.N_285_cascade_\
        );

    \I__420\ : CascadeMux
    port map (
            O => \N__4152\,
            I => \U712_CHIP_RAM.N_309_cascade_\
        );

    \I__419\ : InMux
    port map (
            O => \N__4149\,
            I => \N__4146\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__4146\,
            I => \U712_CHIP_RAM.N_311\
        );

    \I__417\ : CascadeMux
    port map (
            O => \N__4143\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_55_i_a2_0_0_cascade_\
        );

    \I__416\ : InMux
    port map (
            O => \N__4140\,
            I => \N__4134\
        );

    \I__415\ : InMux
    port map (
            O => \N__4139\,
            I => \N__4127\
        );

    \I__414\ : InMux
    port map (
            O => \N__4138\,
            I => \N__4127\
        );

    \I__413\ : InMux
    port map (
            O => \N__4137\,
            I => \N__4127\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__4134\,
            I => \N__4124\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__4127\,
            I => \U712_CHIP_RAM.N_212\
        );

    \I__410\ : Odrv4
    port map (
            O => \N__4124\,
            I => \U712_CHIP_RAM.N_212\
        );

    \I__409\ : CascadeMux
    port map (
            O => \N__4119\,
            I => \U712_CHIP_RAM.N_326_cascade_\
        );

    \I__408\ : CascadeMux
    port map (
            O => \N__4116\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_cascade_\
        );

    \I__407\ : CEMux
    port map (
            O => \N__4113\,
            I => \N__4110\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__4110\,
            I => \N__4107\
        );

    \I__405\ : Odrv4
    port map (
            O => \N__4107\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_0\
        );

    \I__404\ : CascadeMux
    port map (
            O => \N__4104\,
            I => \U712_CHIP_RAM.N_371_cascade_\
        );

    \I__403\ : CascadeMux
    port map (
            O => \N__4101\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_cascade_\
        );

    \I__402\ : CEMux
    port map (
            O => \N__4098\,
            I => \N__4095\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__4095\,
            I => \N__4092\
        );

    \I__400\ : Span4Mux_v
    port map (
            O => \N__4092\,
            I => \N__4089\
        );

    \I__399\ : Odrv4
    port map (
            O => \N__4089\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0\
        );

    \I__398\ : InMux
    port map (
            O => \N__4086\,
            I => \N__4083\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__4083\,
            I => \U712_CHIP_RAM.N_321\
        );

    \I__396\ : InMux
    port map (
            O => \N__4080\,
            I => \N__4077\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__4077\,
            I => \N__4074\
        );

    \I__394\ : Span4Mux_v
    port map (
            O => \N__4074\,
            I => \N__4071\
        );

    \I__393\ : Span4Mux_v
    port map (
            O => \N__4071\,
            I => \N__4068\
        );

    \I__392\ : Sp12to4
    port map (
            O => \N__4068\,
            I => \N__4065\
        );

    \I__391\ : Odrv12
    port map (
            O => \N__4065\,
            I => \A_c_18\
        );

    \I__390\ : InMux
    port map (
            O => \N__4062\,
            I => \N__4059\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__4059\,
            I => \N__4056\
        );

    \I__388\ : Span4Mux_v
    port map (
            O => \N__4056\,
            I => \N__4053\
        );

    \I__387\ : Span4Mux_v
    port map (
            O => \N__4053\,
            I => \N__4050\
        );

    \I__386\ : Sp12to4
    port map (
            O => \N__4050\,
            I => \N__4047\
        );

    \I__385\ : Odrv12
    port map (
            O => \N__4047\,
            I => \A_c_16\
        );

    \I__384\ : IoInMux
    port map (
            O => \N__4044\,
            I => \N__4041\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__4041\,
            I => \N__4038\
        );

    \I__382\ : Span4Mux_s0_h
    port map (
            O => \N__4038\,
            I => \N__4035\
        );

    \I__381\ : Sp12to4
    port map (
            O => \N__4035\,
            I => \N__4032\
        );

    \I__380\ : Span12Mux_v
    port map (
            O => \N__4032\,
            I => \N__4029\
        );

    \I__379\ : Odrv12
    port map (
            O => \N__4029\,
            I => \N_848_i\
        );

    \I__378\ : IoInMux
    port map (
            O => \N__4026\,
            I => \N__4023\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__4023\,
            I => \N__4020\
        );

    \I__376\ : Span12Mux_s8_v
    port map (
            O => \N__4020\,
            I => \N__4017\
        );

    \I__375\ : Odrv12
    port map (
            O => \N__4017\,
            I => \N_336\
        );

    \I__374\ : IoInMux
    port map (
            O => \N__4014\,
            I => \N__4011\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__4011\,
            I => \N__4008\
        );

    \I__372\ : Span12Mux_s3_v
    port map (
            O => \N__4008\,
            I => \N__4005\
        );

    \I__371\ : Odrv12
    port map (
            O => \N__4005\,
            I => \VBENn_c\
        );

    \I__370\ : CascadeMux
    port map (
            O => \N__4002\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER18_cascade_\
        );

    \I__369\ : IoInMux
    port map (
            O => \N__3999\,
            I => \N__3996\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__3996\,
            I => \N__3993\
        );

    \I__367\ : Span4Mux_s2_v
    port map (
            O => \N__3993\,
            I => \N__3990\
        );

    \I__366\ : Span4Mux_v
    port map (
            O => \N__3990\,
            I => \N__3987\
        );

    \I__365\ : Odrv4
    port map (
            O => \N__3987\,
            I => \CLK80_PLL_i_i\
        );

    \I__364\ : IoInMux
    port map (
            O => \N__3984\,
            I => \N__3981\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__3981\,
            I => \N__3978\
        );

    \I__362\ : IoSpan4Mux
    port map (
            O => \N__3978\,
            I => \N__3975\
        );

    \I__361\ : Span4Mux_s3_h
    port map (
            O => \N__3975\,
            I => \N__3972\
        );

    \I__360\ : Odrv4
    port map (
            O => \N__3972\,
            I => \DBRn_c_i_0\
        );

    \I__359\ : InMux
    port map (
            O => \N__3969\,
            I => \N__3966\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__3966\,
            I => \N__3963\
        );

    \I__357\ : Span4Mux_v
    port map (
            O => \N__3963\,
            I => \N__3959\
        );

    \I__356\ : InMux
    port map (
            O => \N__3962\,
            I => \N__3956\
        );

    \I__355\ : Sp12to4
    port map (
            O => \N__3959\,
            I => \N__3951\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__3956\,
            I => \N__3951\
        );

    \I__353\ : Span12Mux_h
    port map (
            O => \N__3951\,
            I => \N__3948\
        );

    \I__352\ : Span12Mux_v
    port map (
            O => \N__3948\,
            I => \N__3945\
        );

    \I__351\ : Odrv12
    port map (
            O => \N__3945\,
            I => \DBRn_c\
        );

    \I__350\ : InMux
    port map (
            O => \N__3942\,
            I => \N__3939\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__3939\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__348\ : InMux
    port map (
            O => \N__3936\,
            I => \N__3933\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__3933\,
            I => \N__3930\
        );

    \I__346\ : Span12Mux_v
    port map (
            O => \N__3930\,
            I => \N__3927\
        );

    \I__345\ : Span12Mux_v
    port map (
            O => \N__3927\,
            I => \N__3924\
        );

    \I__344\ : Odrv12
    port map (
            O => \N__3924\,
            I => \RAMSPACEn_c\
        );

    \I__343\ : IoInMux
    port map (
            O => \N__3921\,
            I => \N__3918\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__3918\,
            I => \N__3915\
        );

    \I__341\ : Span4Mux_s0_v
    port map (
            O => \N__3915\,
            I => \N__3912\
        );

    \I__340\ : Span4Mux_v
    port map (
            O => \N__3912\,
            I => \N__3909\
        );

    \I__339\ : Sp12to4
    port map (
            O => \N__3909\,
            I => \N__3906\
        );

    \I__338\ : Span12Mux_h
    port map (
            O => \N__3906\,
            I => \N__3903\
        );

    \I__337\ : Span12Mux_v
    port map (
            O => \N__3903\,
            I => \N__3900\
        );

    \I__336\ : Odrv12
    port map (
            O => \N__3900\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            I => \N__6864\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            I => \N__6862\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            I => \N__6863\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__6861\
        );

    \INVU712_CHIP_RAM.DMA_A20C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A20C_net\,
            I => \N__6860\
        );

    \IN_MUX_bfv_10_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_6_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_10_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7257\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5510\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3984\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4932\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_3_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8970\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10479\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8648\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBRn_ibuf_RNIBAB_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3962\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBRn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBR_SYNC_1_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3942\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8955\,
            ce => 'H',
            sr => \N__10442\
        );

    \DBR_SYNC_0_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__3969\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8956\,
            ce => 'H',
            sr => \N__10434\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001110011"
        )
    port map (
            in0 => \N__9378\,
            in1 => \N__4274\,
            in2 => \N__4583\,
            in3 => \N__3936\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8943\,
            ce => 'H',
            sr => \N__10451\
        );

    \U712_CHIP_RAM.DBENn_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101111111001100"
        )
    port map (
            in0 => \N__10176\,
            in1 => \N__7693\,
            in2 => \N__4530\,
            in3 => \N__4986\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8943\,
            ce => 'H',
            sr => \N__10451\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4698\,
            in1 => \N__4573\,
            in2 => \N__5334\,
            in3 => \N__4526\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8948\,
            ce => \N__4113\,
            sr => \N__10443\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__4697\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4572\,
            lcout => \U712_CHIP_RAM.N_212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9209\,
            in1 => \N__4080\,
            in2 => \_gnd_net_\,
            in3 => \N__4062\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__4217\,
            in1 => \N__6298\,
            in2 => \_gnd_net_\,
            in3 => \N__5398\,
            lcout => \WRITE_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8952\,
            ce => \N__4098\,
            sr => \N__10435\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4299\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8957\,
            ce => 'H',
            sr => \N__10420\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__7560\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7836\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8961\,
            ce => 'H',
            sr => \N__10413\
        );

    \TACKn_obuft_RNO_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4287\,
            lcout => \N_848_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DMA_LATCH_EN_i_i_a2_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__7553\,
            in1 => \N__7827\,
            in2 => \_gnd_net_\,
            in3 => \N__6242\,
            lcout => \N_336\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_0_a2_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4413\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9423\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5058\,
            in1 => \N__6769\,
            in2 => \N__6042\,
            in3 => \N__5799\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4002\,
            in3 => \N__5856\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8934\,
            ce => 'H',
            sr => \N__10444\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4HBB7_2_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4514\,
            in2 => \_gnd_net_\,
            in3 => \N__6147\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__4137\,
            in1 => \N__4195\,
            in2 => \N__5332\,
            in3 => \N__4086\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10477\,
            in1 => \_gnd_net_\,
            in2 => \N__4116\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIGGM16_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__4139\,
            in1 => \N__7353\,
            in2 => \N__5333\,
            in3 => \N__4196\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_2_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6755\,
            in2 => \_gnd_net_\,
            in3 => \N__6156\,
            lcout => \U712_CHIP_RAM.N_371\,
            ltout => \U712_CHIP_RAM.N_371_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIQ6QH5_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000010000"
        )
    port map (
            in0 => \N__4138\,
            in1 => \N__6542\,
            in2 => \N__4104\,
            in3 => \N__5400\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10478\,
            in1 => \_gnd_net_\,
            in2 => \N__4101\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__5442\,
            in1 => \N__5004\,
            in2 => \_gnd_net_\,
            in3 => \N__6014\,
            lcout => \U712_CHIP_RAM.N_321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__4959\,
            in1 => \N__7354\,
            in2 => \N__4476\,
            in3 => \N__5217\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8944\,
            ce => \N__5176\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__7376\,
            in1 => \N__5396\,
            in2 => \N__6546\,
            in3 => \N__6155\,
            lcout => \U712_CHIP_RAM.N_311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBDIR_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111010011110000"
        )
    port map (
            in0 => \N__4218\,
            in1 => \N__5397\,
            in2 => \N__4172\,
            in3 => \N__4197\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8949\,
            ce => 'H',
            sr => \N__10425\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6768\,
            in2 => \_gnd_net_\,
            in3 => \N__6154\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_285_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111110011"
        )
    port map (
            in0 => \N__4622\,
            in1 => \N__7377\,
            in2 => \N__4155\,
            in3 => \N__5057\,
            lcout => \U712_CHIP_RAM.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4776\,
            in2 => \_gnd_net_\,
            in3 => \N__5280\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_309_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__5873\,
            in1 => \N__5798\,
            in2 => \N__4152\,
            in3 => \N__4419\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_55_i_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000011"
        )
    port map (
            in0 => \N__9198\,
            in1 => \N__4149\,
            in2 => \N__4143\,
            in3 => \N__4607\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8953\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIHOOI5_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6159\,
            in1 => \N__7331\,
            in2 => \N__5331\,
            in3 => \N__4140\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_326_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI77IM9_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__5412\,
            in1 => \N__5872\,
            in2 => \N__4119\,
            in3 => \N__5797\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI12QHH_2_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__6798\,
            in1 => \N__4785\,
            in2 => \N__4338\,
            in3 => \N__7332\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4335\,
            in1 => \N__4317\,
            in2 => \_gnd_net_\,
            in3 => \N__9197\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4305\,
            in2 => \_gnd_net_\,
            in3 => \N__4298\,
            lcout => \U712_CHIP_RAM.un3_DMA_CYCLE_START\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__7330\,
            in1 => \N__6614\,
            in2 => \_gnd_net_\,
            in3 => \N__6648\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8958\,
            ce => \N__4734\,
            sr => \N__10409\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000001111"
        )
    port map (
            in0 => \N__6409\,
            in1 => \N__5577\,
            in2 => \N__4820\,
            in3 => \N__4881\,
            lcout => \U712_REG_SM.STATE_COUNTc_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_0_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4943\,
            in2 => \_gnd_net_\,
            in3 => \N__6410\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_294_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011100100"
        )
    port map (
            in0 => \N__7281\,
            in1 => \N__4402\,
            in2 => \N__4281\,
            in3 => \N__5532\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8962\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011000000110001"
        )
    port map (
            in0 => \N__6500\,
            in1 => \N__5618\,
            in2 => \N__4890\,
            in3 => \N__6467\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8963\,
            ce => 'H',
            sr => \N__10401\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011100000011"
        )
    port map (
            in0 => \N__4401\,
            in1 => \N__4278\,
            in2 => \N__4242\,
            in3 => \N__4851\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8963\,
            ce => 'H',
            sr => \N__10401\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100011111100"
        )
    port map (
            in0 => \N__4880\,
            in1 => \N__5586\,
            in2 => \N__6414\,
            in3 => \N__4836\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8966\,
            ce => 'H',
            sr => \N__10400\
        );

    \U712_BUFFERS.un1_DRDENn_0_a2_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__7527\,
            in1 => \N__7823\,
            in2 => \_gnd_net_\,
            in3 => \N__4409\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_0_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4641\,
            in2 => \_gnd_net_\,
            in3 => \N__5006\,
            lcout => \U712_CHIP_RAM.N_331\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__7898\,
            in1 => \N__5392\,
            in2 => \_gnd_net_\,
            in3 => \N__4515\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.LATCH_CLK_8_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__5032\,
            in1 => \N__5789\,
            in2 => \N__4347\,
            in3 => \N__6036\,
            lcout => \U712_CHIP_RAM.N_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3FV43_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5860\,
            in1 => \N__5782\,
            in2 => \_gnd_net_\,
            in3 => \N__5031\,
            lcout => \U712_CHIP_RAM.N_397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNI7MCB2_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__5391\,
            in1 => \N__6754\,
            in2 => \_gnd_net_\,
            in3 => \N__4763\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_368_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIGK316_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__5861\,
            in1 => \N__5783\,
            in2 => \N__4344\,
            in3 => \N__5013\,
            lcout => \U712_CHIP_RAM.N_323\,
            ltout => \U712_CHIP_RAM.N_323_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIHBKDA_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__5262\,
            in1 => \N__6237\,
            in2 => \N__4341\,
            in3 => \N__5005\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5907\,
            in1 => \N__5995\,
            in2 => \_gnd_net_\,
            in3 => \N__5663\,
            lcout => \U712_CHIP_RAM.N_359\,
            ltout => \U712_CHIP_RAM.N_359_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__5751\,
            in1 => \_gnd_net_\,
            in2 => \N__4587\,
            in3 => \N__6746\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER15\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIVLD65_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5327\,
            in1 => \N__4584\,
            in2 => \N__4554\,
            in3 => \N__4718\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_2_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__10710\,
            in1 => \_gnd_net_\,
            in2 => \N__4551\,
            in3 => \N__4548\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_330_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_1_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__4522\,
            in1 => \N__5384\,
            in2 => \N__4491\,
            in3 => \N__8628\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.BANK0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__4488\,
            in1 => \N__4448\,
            in2 => \N__4479\,
            in3 => \N__4475\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8935\,
            ce => 'H',
            sr => \N__10426\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI05TJ3_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5834\,
            in1 => \N__4762\,
            in2 => \_gnd_net_\,
            in3 => \N__5750\,
            lcout => \U712_CHIP_RAM.N_360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5OHEF_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101110111011"
        )
    port map (
            in0 => \N__4437\,
            in1 => \N__7375\,
            in2 => \N__4623\,
            in3 => \N__5056\,
            lcout => \U712_CHIP_RAM.N_49\,
            ltout => \U712_CHIP_RAM.N_49_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001101011100"
        )
    port map (
            in0 => \N__4428\,
            in1 => \N__7136\,
            in2 => \N__4422\,
            in3 => \N__6005\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8945\,
            ce => \N__5180\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6742\,
            in1 => \N__5683\,
            in2 => \N__6033\,
            in3 => \N__7374\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_55_i_a2_0_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_2_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6740\,
            in2 => \_gnd_net_\,
            in3 => \N__6001\,
            lcout => \U712_CHIP_RAM.N_403\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1IJO_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__6741\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6217\,
            lcout => \U712_CHIP_RAM.N_207\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011010001"
        )
    port map (
            in0 => \N__5286\,
            in1 => \N__4605\,
            in2 => \N__8101\,
            in3 => \N__5235\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8950\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000100000001"
        )
    port map (
            in0 => \N__4746\,
            in1 => \N__6672\,
            in2 => \N__4608\,
            in3 => \N__8346\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8950\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI1DV43_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__5862\,
            in1 => \N__6006\,
            in2 => \N__5784\,
            in3 => \N__6792\,
            lcout => \U712_CHIP_RAM.N_361\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4677\,
            in1 => \N__4659\,
            in2 => \_gnd_net_\,
            in3 => \N__9199\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI71B91_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7897\,
            in1 => \N__6007\,
            in2 => \_gnd_net_\,
            in3 => \N__5443\,
            lcout => \U712_CHIP_RAM.N_217\,
            ltout => \U712_CHIP_RAM.N_217_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIDDEL6_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__4632\,
            in1 => \N__5760\,
            in2 => \N__4626\,
            in3 => \N__5863\,
            lcout => \U712_CHIP_RAM.N_222\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011010001"
        )
    port map (
            in0 => \N__4971\,
            in1 => \N__4606\,
            in2 => \N__8433\,
            in3 => \N__4745\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8950\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5PDS6_0_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__5055\,
            in1 => \N__5761\,
            in2 => \N__6034\,
            in3 => \N__6158\,
            lcout => \U712_CHIP_RAM.N_262\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__6784\,
            in1 => \N__5925\,
            in2 => \N__5697\,
            in3 => \N__6035\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_354_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIFJSJ3_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__5696\,
            in1 => \N__5261\,
            in2 => \N__4779\,
            in3 => \N__5875\,
            lcout => \U712_CHIP_RAM.N_408\,
            ltout => \U712_CHIP_RAM.N_408_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI997R7_2_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010100000"
        )
    port map (
            in0 => \N__5276\,
            in1 => \N__6785\,
            in2 => \N__4770\,
            in3 => \N__4767\,
            lcout => \U712_CHIP_RAM.N_305\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101010"
        )
    port map (
            in0 => \N__6519\,
            in1 => \N__7329\,
            in2 => \N__6615\,
            in3 => \N__6636\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_236_i_0_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10474\,
            in1 => \_gnd_net_\,
            in2 => \N__4737\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.N_236_i_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNITI8N_2_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__4812\,
            in1 => \N__5575\,
            in2 => \_gnd_net_\,
            in3 => \N__4717\,
            lcout => \U712_REG_SM.N_255\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_1_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4896\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8959\,
            ce => 'H',
            sr => \N__10402\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__5581\,
            in1 => \N__4728\,
            in2 => \N__4722\,
            in3 => \N__6398\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8959\,
            ce => 'H',
            sr => \N__10402\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100001011"
        )
    port map (
            in0 => \N__6397\,
            in1 => \N__5582\,
            in2 => \N__4947\,
            in3 => \N__6501\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8959\,
            ce => 'H',
            sr => \N__10402\
        );

    \U712_REG_SM.C3_SYNC_0_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4916\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8959\,
            ce => 'H',
            sr => \N__10402\
        );

    \U712_REG_SM.STATE_COUNT_RNIVCF31_1_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011011111"
        )
    port map (
            in0 => \N__6451\,
            in1 => \N__5572\,
            in2 => \N__6399\,
            in3 => \N__4875\,
            lcout => \U712_REG_SM.N_239\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_0_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__6299\,
            in1 => \N__4813\,
            in2 => \_gnd_net_\,
            in3 => \N__6453\,
            lcout => \U712_REG_SM.N_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4850\,
            in1 => \N__6455\,
            in2 => \_gnd_net_\,
            in3 => \N__6498\,
            lcout => \U712_REG_SM.STATE_COUNT_srsts_i_0_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4811\,
            in2 => \_gnd_net_\,
            in3 => \N__4876\,
            lcout => \U712_REG_SM.N_232\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__6393\,
            in1 => \N__4857\,
            in2 => \_gnd_net_\,
            in3 => \N__4849\,
            lcout => \U712_REG_SM.N_264\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__6452\,
            in1 => \N__5573\,
            in2 => \_gnd_net_\,
            in3 => \N__6392\,
            lcout => \U712_REG_SM.N_216\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110101010001"
        )
    port map (
            in0 => \N__4830\,
            in1 => \N__6426\,
            in2 => \N__4824\,
            in3 => \N__9863\,
            lcout => \DS_ENm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8964\,
            ce => 'H',
            sr => \N__10398\
        );

    \U712_CHIP_RAM.LATCH_CLK_LC_10_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010011111110"
        )
    port map (
            in0 => \N__5100\,
            in1 => \N__5069\,
            in2 => \N__6840\,
            in3 => \N__5094\,
            lcout => \LATCH_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8925\,
            ce => 'H',
            sr => \N__10436\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5908\,
            in2 => \_gnd_net_\,
            in3 => \N__5664\,
            lcout => \U712_CHIP_RAM.N_363\,
            ltout => \U712_CHIP_RAM.N_363_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI4VIE1_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7864\,
            in2 => \N__5016\,
            in3 => \N__6031\,
            lcout => \U712_CHIP_RAM.N_369\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__9424\,
            in1 => \N__5909\,
            in2 => \_gnd_net_\,
            in3 => \N__5665\,
            lcout => \U712_CHIP_RAM.CLK_EN_5_0_a2_1_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI1NGC4_0_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__5451\,
            in1 => \N__5007\,
            in2 => \_gnd_net_\,
            in3 => \N__6032\,
            lcout => \U712_CHIP_RAM.N_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10476\,
            in2 => \_gnd_net_\,
            in3 => \N__4982\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6021\,
            in2 => \_gnd_net_\,
            in3 => \N__6665\,
            lcout => \U712_CHIP_RAM.N_306\,
            ltout => OPEN,
            carryin => \bfn_10_6_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5214\,
            in1 => \N__5691\,
            in2 => \_gnd_net_\,
            in3 => \N__4962\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__8929\,
            ce => \N__5184\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6786\,
            in2 => \_gnd_net_\,
            in3 => \N__4950\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5215\,
            in1 => \N__5921\,
            in2 => \_gnd_net_\,
            in3 => \N__5229\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__8929\,
            ce => \N__5184\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5211\,
            in1 => \N__5148\,
            in2 => \_gnd_net_\,
            in3 => \N__5226\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__8929\,
            ce => \N__5184\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5216\,
            in1 => \N__5132\,
            in2 => \_gnd_net_\,
            in3 => \N__5223\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__8929\,
            ce => \N__5184\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5212\,
            in1 => \N__5160\,
            in2 => \_gnd_net_\,
            in3 => \N__5220\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__8929\,
            ce => \N__5184\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__5118\,
            in1 => \N__5213\,
            in2 => \_gnd_net_\,
            in3 => \N__5187\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8929\,
            ce => \N__5184\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5159\,
            in1 => \N__5147\,
            in2 => \N__5136\,
            in3 => \N__5117\,
            lcout => \U712_CHIP_RAM.N_352\,
            ltout => \U712_CHIP_RAM.N_352_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3M1M2_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__5666\,
            in1 => \_gnd_net_\,
            in2 => \N__5106\,
            in3 => \N__5874\,
            lcout => \U712_CHIP_RAM.N_396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6065\,
            in1 => \N__5457\,
            in2 => \N__9512\,
            in3 => \N__5775\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_328_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__5671\,
            in1 => \N__6236\,
            in2 => \N__5103\,
            in3 => \N__9483\,
            lcout => \U712_CHIP_RAM.N_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011111000"
        )
    port map (
            in0 => \N__5469\,
            in1 => \N__7372\,
            in2 => \N__5399\,
            in3 => \N__7876\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__5670\,
            in1 => \N__6235\,
            in2 => \_gnd_net_\,
            in3 => \N__6012\,
            lcout => \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__6013\,
            in1 => \N__5447\,
            in2 => \N__5793\,
            in3 => \N__5421\,
            lcout => \U712_CHIP_RAM.CLK_EN_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIHFLS1_3_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__7373\,
            in1 => \N__5910\,
            in2 => \N__5684\,
            in3 => \N__6011\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIRILU_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6530\,
            in2 => \_gnd_net_\,
            in3 => \N__5375\,
            lcout => \U712_CHIP_RAM.N_370\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__6238\,
            in1 => \N__6664\,
            in2 => \_gnd_net_\,
            in3 => \N__6022\,
            lcout => \U712_CHIP_RAM.N_307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__7342\,
            in1 => \N__5762\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_411\,
            ltout => \U712_CHIP_RAM.N_411_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5924\,
            in1 => \N__5260\,
            in2 => \N__5238\,
            in3 => \N__5877\,
            lcout => \U712_CHIP_RAM.N_308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6793\,
            in2 => \_gnd_net_\,
            in3 => \N__5922\,
            lcout => \U712_CHIP_RAM.N_404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_3_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5923\,
            in1 => \N__5876\,
            in2 => \N__5785\,
            in3 => \N__5692\,
            lcout => \U712_CHIP_RAM.N_313_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8337\,
            in1 => \N__8404\,
            in2 => \N__8076\,
            in3 => \N__9235\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__6813\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5603\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__5622\,
            in1 => \N__5520\,
            in2 => \N__5607\,
            in3 => \N__5592\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8954\,
            ce => 'H',
            sr => \N__10403\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__6391\,
            in1 => \N__5576\,
            in2 => \_gnd_net_\,
            in3 => \N__6497\,
            lcout => \U712_REG_SM.N_289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__6454\,
            in1 => \N__5574\,
            in2 => \_gnd_net_\,
            in3 => \N__6390\,
            lcout => \U712_REG_SM.N_254\,
            ltout => \U712_REG_SM.N_254_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6300\,
            in2 => \N__5523\,
            in3 => \N__6496\,
            lcout => \U712_REG_SM.N_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_1_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5475\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8960\,
            ce => 'H',
            sr => \N__10399\
        );

    \U712_REG_SM.C1_SYNC_0_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5514\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8960\,
            ce => 'H',
            sr => \N__10399\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__6499\,
            in1 => \N__6468\,
            in2 => \_gnd_net_\,
            in3 => \N__6456\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8960\,
            ce => 'H',
            sr => \N__10399\
        );

    \U712_REG_SM.ASn_ess_RNO_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10473\,
            in2 => \_gnd_net_\,
            in3 => \N__6425\,
            lcout => \U712_REG_SM.N_239_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_ess_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6405\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8965\,
            ce => \N__6306\,
            sr => \N__10394\
        );

    \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001111111"
        )
    port map (
            in0 => \N__6283\,
            in1 => \N__7793\,
            in2 => \N__7552\,
            in3 => \N__6246\,
            lcout => \N_259\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6797\,
            in2 => \_gnd_net_\,
            in3 => \N__6157\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8926\,
            ce => \N__6114\,
            sr => \N__10414\
        );

    \U712_CHIP_RAM.CLK_EN_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111111100001000"
        )
    port map (
            in0 => \N__6054\,
            in1 => \N__6041\,
            in2 => \N__6102\,
            in3 => \N__6077\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8930\,
            ce => 'H',
            sr => \N__10410\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6681\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6066\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_312_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__6053\,
            in1 => \N__6791\,
            in2 => \N__6045\,
            in3 => \N__6040\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__6812\,
            in1 => \N__6839\,
            in2 => \N__6822\,
            in3 => \N__6819\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8930\,
            ce => 'H',
            sr => \N__10410\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIONRK3_2_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7356\,
            in1 => \N__6790\,
            in2 => \_gnd_net_\,
            in3 => \N__6680\,
            lcout => \U712_CHIP_RAM.N_400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100011111000"
        )
    port map (
            in0 => \N__7062\,
            in1 => \N__6584\,
            in2 => \N__6610\,
            in3 => \N__6643\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8937\,
            ce => 'H',
            sr => \N__10405\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__6583\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7063\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8937\,
            ce => 'H',
            sr => \N__10405\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001100100000"
        )
    port map (
            in0 => \N__6945\,
            in1 => \N__6582\,
            in2 => \N__6647\,
            in3 => \N__6515\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8937\,
            ce => 'H',
            sr => \N__10405\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6959\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8937\,
            ce => 'H',
            sr => \N__10405\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110100010"
        )
    port map (
            in0 => \N__6557\,
            in1 => \N__6585\,
            in2 => \N__7068\,
            in3 => \N__6974\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8946\,
            ce => 'H',
            sr => \N__10404\
        );

    \U712_CHIP_RAM.REFRESH_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6896\,
            in1 => \N__6911\,
            in2 => \N__6879\,
            in3 => \N__7152\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8946\,
            ce => 'H',
            sr => \N__10404\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6975\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8946\,
            ce => 'H',
            sr => \N__10404\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6939\,
            in2 => \_gnd_net_\,
            in3 => \N__6933\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__6859\,
            ce => 'H',
            sr => \N__7194\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6930\,
            in2 => \_gnd_net_\,
            in3 => \N__6924\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__6859\,
            ce => 'H',
            sr => \N__7194\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7164\,
            in2 => \_gnd_net_\,
            in3 => \N__6921\,
            lcout => \U712_CHIP_RAM.REFRESH5lto2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__6859\,
            ce => 'H',
            sr => \N__7194\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7176\,
            in2 => \_gnd_net_\,
            in3 => \N__6918\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__6859\,
            ce => 'H',
            sr => \N__7194\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7188\,
            in2 => \_gnd_net_\,
            in3 => \N__6915\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__6859\,
            ce => 'H',
            sr => \N__7194\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6912\,
            in2 => \_gnd_net_\,
            in3 => \N__6900\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__6859\,
            ce => 'H',
            sr => \N__7194\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6897\,
            in2 => \_gnd_net_\,
            in3 => \N__6885\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__6859\,
            ce => 'H',
            sr => \N__7194\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6875\,
            in2 => \_gnd_net_\,
            in3 => \N__6882\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6859\,
            ce => 'H',
            sr => \N__7194\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7187\,
            in1 => \N__7175\,
            in2 => \_gnd_net_\,
            in3 => \N__7163\,
            lcout => \U712_CHIP_RAM.REFRESH5lt7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIHMEA_1_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9396\,
            in2 => \_gnd_net_\,
            in3 => \N__9273\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_RNIHMEAZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7113\,
            in1 => \N__9422\,
            in2 => \_gnd_net_\,
            in3 => \N__10161\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_231_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9073\,
            in2 => \N__7098\,
            in3 => \N__9274\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__8137\,
            in1 => \N__7091\,
            in2 => \N__9513\,
            in3 => \N__9950\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110111011"
        )
    port map (
            in0 => \N__9951\,
            in1 => \N__8138\,
            in2 => \N__7095\,
            in3 => \N__9487\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_RNI8MQ3_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__7067\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6973\,
            in2 => \_gnd_net_\,
            in3 => \N__6960\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9475\,
            in1 => \N__7446\,
            in2 => \N__9272\,
            in3 => \N__10293\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__9250\,
            in1 => \N__8423\,
            in2 => \_gnd_net_\,
            in3 => \N__8089\,
            lcout => \U712_CHIP_RAM.CMA_5_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7437\,
            in1 => \N__7416\,
            in2 => \_gnd_net_\,
            in3 => \N__9251\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_180_i_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101010101"
        )
    port map (
            in0 => \N__8265\,
            in1 => \N__7724\,
            in2 => \N__7832\,
            in3 => \N__7899\,
            lcout => \N_180_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7355\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__9075\,
            in1 => \N__9621\,
            in2 => \N__9031\,
            in3 => \N__7245\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8927\,
            ce => \N__8836\,
            sr => \N__10415\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100001000"
        )
    port map (
            in0 => \N__8760\,
            in1 => \N__9279\,
            in2 => \N__9516\,
            in3 => \N__9074\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7656\,
            in2 => \N__7215\,
            in3 => \N__7605\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8931\,
            ce => \N__8815\,
            sr => \N__10411\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8437\,
            in2 => \_gnd_net_\,
            in3 => \N__8097\,
            lcout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\,
            ltout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101011101"
        )
    port map (
            in0 => \N__9278\,
            in1 => \N__8759\,
            in2 => \N__7659\,
            in3 => \N__9494\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7650\,
            in1 => \N__7644\,
            in2 => \_gnd_net_\,
            in3 => \N__7638\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8931\,
            ce => \N__8815\,
            sr => \N__10411\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000010011"
        )
    port map (
            in0 => \N__8422\,
            in1 => \N__8347\,
            in2 => \N__9244\,
            in3 => \N__8093\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9214\,
            in1 => \N__7611\,
            in2 => \N__9511\,
            in3 => \N__9549\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7599\,
            in1 => \N__7578\,
            in2 => \_gnd_net_\,
            in3 => \N__9213\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__7725\,
            in1 => \N__7550\,
            in2 => \_gnd_net_\,
            in3 => \N__7900\,
            lcout => \U712_BYTE_ENABLE.N_342\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7726\,
            in1 => \N__7551\,
            in2 => \_gnd_net_\,
            in3 => \N__7901\,
            lcout => \U712_BYTE_ENABLE.N_320\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000000000"
        )
    port map (
            in0 => \N__8594\,
            in1 => \N__9851\,
            in2 => \N__9759\,
            in3 => \N__9503\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_341_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_55_i_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__9502\,
            in1 => \N__7476\,
            in2 => \N__7470\,
            in3 => \N__8285\,
            lcout => \N_55_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100000000"
        )
    port map (
            in0 => \N__9758\,
            in1 => \N__9852\,
            in2 => \N__8598\,
            in3 => \N__9504\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_318_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_105_i_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__9501\,
            in1 => \N__8010\,
            in2 => \N__8004\,
            in3 => \N__8284\,
            lcout => \N_105_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_x2_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9743\,
            in2 => \_gnd_net_\,
            in3 => \N__8516\,
            lcout => \U712_BYTE_ENABLE.N_206_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__9084\,
            in1 => \N__9633\,
            in2 => \N__9042\,
            in3 => \N__7917\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8932\,
            ce => \N__8835\,
            sr => \N__10421\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10475\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7959\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7953\,
            in1 => \N__7938\,
            in2 => \_gnd_net_\,
            in3 => \N__9280\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9281\,
            in1 => \N__9476\,
            in2 => \N__7920\,
            in3 => \N__10254\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9282\,
            in1 => \N__7908\,
            in2 => \N__9517\,
            in3 => \N__9912\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_57_i_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110001"
        )
    port map (
            in0 => \N__7902\,
            in1 => \N__8301\,
            in2 => \N__7831\,
            in3 => \N__7733\,
            lcout => \N_57_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110000"
        )
    port map (
            in0 => \N__9849\,
            in1 => \N__8592\,
            in2 => \N__9518\,
            in3 => \N__8294\,
            lcout => \U712_BYTE_ENABLE.N_339\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011110000"
        )
    port map (
            in0 => \N__9850\,
            in1 => \N__8593\,
            in2 => \N__9519\,
            in3 => \N__8295\,
            lcout => \U712_BYTE_ENABLE.N_316\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_277_i_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010010101000"
        )
    port map (
            in0 => \N__9733\,
            in1 => \N__9833\,
            in2 => \N__8581\,
            in3 => \N__8495\,
            lcout => \N_277_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LLBE_i_o2_i_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100110000"
        )
    port map (
            in0 => \N__9832\,
            in1 => \N__8570\,
            in2 => \N__8505\,
            in3 => \N__9732\,
            lcout => \LLBE_i_o2_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WEn_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8103\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8928\,
            ce => 'H',
            sr => \N__10445\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__8147\,
            in1 => \N__8205\,
            in2 => \N__9515\,
            in3 => \N__9642\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8938\,
            ce => \N__8837\,
            sr => \N__10427\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__8166\,
            in1 => \N__8769\,
            in2 => \N__9514\,
            in3 => \N__8148\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8938\,
            ce => \N__8837\,
            sr => \N__10427\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8444\,
            in1 => \N__9294\,
            in2 => \N__8361\,
            in3 => \N__8102\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8947\,
            ce => \N__8831\,
            sr => \N__10422\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__9085\,
            in1 => \N__9918\,
            in2 => \N__9043\,
            in3 => \N__8733\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8947\,
            ce => \N__8831\,
            sr => \N__10422\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9473\,
            in1 => \N__8706\,
            in2 => \N__9295\,
            in3 => \N__10098\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8694\,
            in1 => \N__8676\,
            in2 => \_gnd_net_\,
            in3 => \N__9283\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9284\,
            in1 => \N__9474\,
            in2 => \N__8655\,
            in3 => \N__10146\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_A20_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__8652\,
            in1 => \N__10680\,
            in2 => \N__10766\,
            in3 => \N__8624\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A20C_net\,
            ce => 'H',
            sr => \N__10412\
        );

    \U712_BYTE_ENABLE.UMBE_0_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110100000"
        )
    port map (
            in0 => \N__8544\,
            in1 => \N__9834\,
            in2 => \N__8520\,
            in3 => \N__9749\,
            lcout => \UMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_276_i_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000110100010"
        )
    port map (
            in0 => \N__9747\,
            in1 => \N__8574\,
            in2 => \N__9848\,
            in3 => \N__8515\,
            lcout => \N_276_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RASn_LC_16_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8445\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8933\,
            ce => 'H',
            sr => \N__10452\
        );

    \U712_CHIP_RAM.CRCSn_LC_16_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8357\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8933\,
            ce => 'H',
            sr => \N__10452\
        );

    \U712_CHIP_RAM.CASn_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9299\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8939\,
            ce => 'H',
            sr => \N__10446\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9472\,
            in1 => \N__9312\,
            in2 => \N__9300\,
            in3 => \N__10521\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__9094\,
            in1 => \N__10038\,
            in2 => \N__9044\,
            in3 => \N__9141\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8951\,
            ce => \N__8841\,
            sr => \N__10428\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__9095\,
            in1 => \N__9609\,
            in2 => \N__9045\,
            in3 => \N__9120\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8951\,
            ce => \N__8841\,
            sr => \N__10428\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__9096\,
            in1 => \N__9041\,
            in2 => \N__8742\,
            in3 => \N__8994\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8951\,
            ce => \N__8841\,
            sr => \N__10428\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10767\,
            in1 => \N__10660\,
            in2 => \_gnd_net_\,
            in3 => \N__8781\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9934\,
            ce => \N__10503\,
            sr => \N__10423\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__10245\,
            in1 => \_gnd_net_\,
            in2 => \N__10693\,
            in3 => \N__9603\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9934\,
            ce => \N__10503\,
            sr => \N__10423\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__10026\,
            in1 => \_gnd_net_\,
            in2 => \N__10694\,
            in3 => \N__10133\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9934\,
            ce => \N__10503\,
            sr => \N__10423\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10200\,
            in1 => \N__10653\,
            in2 => \_gnd_net_\,
            in3 => \N__10244\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9934\,
            ce => \N__10503\,
            sr => \N__10423\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9597\,
            in1 => \N__10679\,
            in2 => \_gnd_net_\,
            in3 => \N__10235\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__10502\,
            sr => \N__10416\
        );

    \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011111111"
        )
    port map (
            in0 => \N__9830\,
            in1 => \N__9712\,
            in2 => \_gnd_net_\,
            in3 => \N__9881\,
            lcout => \un1_LDSn_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__9882\,
            in1 => \N__9831\,
            in2 => \_gnd_net_\,
            in3 => \N__9748\,
            lcout => \N_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10554\,
            in1 => \N__10703\,
            in2 => \_gnd_net_\,
            in3 => \N__10753\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9936\,
            ce => \N__10509\,
            sr => \N__10447\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9599\,
            in1 => \N__10688\,
            in2 => \_gnd_net_\,
            in3 => \N__10283\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9935\,
            ce => \N__10507\,
            sr => \N__10437\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__10284\,
            in1 => \_gnd_net_\,
            in2 => \N__10708\,
            in3 => \N__10084\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9935\,
            ce => \N__10507\,
            sr => \N__10437\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10692\,
            in1 => \N__10553\,
            in2 => \_gnd_net_\,
            in3 => \N__10134\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9935\,
            ce => \N__10507\,
            sr => \N__10437\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10276\,
            in1 => \N__10697\,
            in2 => \_gnd_net_\,
            in3 => \N__9598\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__10505\,
            sr => \N__10429\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__10086\,
            in1 => \_gnd_net_\,
            in2 => \N__10709\,
            in3 => \N__9984\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__10505\,
            sr => \N__10429\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10277\,
            in1 => \N__10698\,
            in2 => \_gnd_net_\,
            in3 => \N__10085\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__10505\,
            sr => \N__10429\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10696\,
            in1 => \N__10234\,
            in2 => \_gnd_net_\,
            in3 => \N__10199\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__10505\,
            sr => \N__10429\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10132\,
            in1 => \N__10022\,
            in2 => \_gnd_net_\,
            in3 => \N__10702\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__10505\,
            sr => \N__10429\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10020\,
            in1 => \N__10661\,
            in2 => \_gnd_net_\,
            in3 => \N__9980\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__10504\,
            sr => \N__10424\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__10546\,
            in1 => \_gnd_net_\,
            in2 => \N__10695\,
            in3 => \N__10131\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__10504\,
            sr => \N__10424\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9978\,
            in1 => \N__10684\,
            in2 => \_gnd_net_\,
            in3 => \N__10075\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9933\,
            ce => \N__10508\,
            sr => \N__10438\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__10021\,
            in1 => \_gnd_net_\,
            in2 => \N__10707\,
            in3 => \N__9979\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9933\,
            ce => \N__10508\,
            sr => \N__10438\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10744\,
            in1 => \N__10621\,
            in2 => \_gnd_net_\,
            in3 => \N__10537\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__10506\,
            sr => \N__10430\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     May 8 2025 19:39:33

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    DA : out std_logic_vector(2 downto 0);
    A : in std_logic_vector(20 downto 0);
    DBRn : in std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    TCIn : out std_logic;
    TBIn : out std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__12710\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10629\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10380\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7827\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7434\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7344\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \bfn_6_6_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_7\ : std_logic;
signal \A_c_8\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_CHIP_RAM.m93_i_a2_4_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto7_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lt7\ : std_logic;
signal \U712_CHIP_RAM.N_430_cascade_\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.N_428\ : std_logic;
signal \U712_CHIP_RAM.N_307_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_467_cascade_\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_0\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \TSn_c\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \U712_CHIP_RAM.N_419\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_5_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDs_0_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_1_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_396_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_0_2\ : std_logic;
signal \U712_CHIP_RAM.N_397\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_1_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDs_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_194_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_1\ : std_logic;
signal \U712_CHIP_RAM.N_305_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\ : std_logic;
signal \U712_CHIP_RAM.N_325\ : std_logic;
signal \U712_CHIP_RAM.N_325_cascade_\ : std_logic;
signal \U712_CHIP_RAM.m101_i_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.m101_i_1\ : std_logic;
signal \U712_CHIP_RAM.N_376\ : std_logic;
signal \U712_CHIP_RAM.m101_i_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_436\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_378\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_551_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER41_0_a3_0_a2_0\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \U712_REG_SM.N_412\ : std_logic;
signal \U712_REG_SM.N_402\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_0\ : std_logic;
signal \REGENn_c\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.REGENn_e_1\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.N_555\ : std_logic;
signal \U712_CHIP_RAM.N_555_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_194\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_2_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_449\ : std_logic;
signal \U712_CHIP_RAM.N_476\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_304_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_312_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_326_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_467\ : std_logic;
signal \U712_CHIP_RAM.N_39\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \U712_CHIP_RAM.N_440\ : std_logic;
signal \U712_CHIP_RAM.N_39_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_326\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.DBENn_7_0_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_344_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_551\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER41_2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.LATCH_CLK_6\ : std_logic;
signal \LATCH_CLK_c\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_435\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_413_cascade_\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \U712_REG_SM.N_308\ : std_logic;
signal \U712_REG_SM.N_308_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ1Z_2\ : std_logic;
signal \U712_REG_SM.N_410_cascade_\ : std_logic;
signal \U712_REG_SM.N_331\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U712_REG_SM.N_404\ : std_logic;
signal \LDSn_c\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_459\ : std_logic;
signal \UDSn_c\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_0\ : std_logic;
signal \bfn_10_5_0_\ : std_logic;
signal \U712_CHIP_RAM.un3_DBR_COUNT_cry_1\ : std_logic;
signal \U712_CHIP_RAM.un3_DBR_COUNT_cry_2\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.un3_DBR_COUNT_cry_3\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.un3_DBR_COUNT_cry_4\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.un3_DBR_COUNT_cry_5\ : std_logic;
signal \U712_CHIP_RAM.un3_DBR_COUNT_cry_6\ : std_logic;
signal \A_c_12\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DBR_COUNTZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.m93_i_a2_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.N_304\ : std_logic;
signal \U712_CHIP_RAM.N_305\ : std_logic;
signal \U712_CHIP_RAM.m123_i_2_cascade_\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_2_0\ : std_logic;
signal \U712_CHIP_RAM.N_390\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_2_3\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\ : std_logic;
signal \A_c_6\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \N_167_i\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.N_321\ : std_logic;
signal \U712_CHIP_RAM.N_321_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_20_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.m77_0_a2_0_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_307\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_6\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \N_202_i\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \U712_REG_SM.N_328\ : std_logic;
signal \U712_REG_SM.N_406\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_330_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_2\ : std_logic;
signal \U712_REG_SM.STATE_COUNTc_0_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_373\ : std_logic;
signal \U712_REG_SM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.N_373_cascade_\ : std_logic;
signal \U712_REG_SM.N_130\ : std_logic;
signal \U712_REG_SM.un1_REGENn_0_sqmuxa_0\ : std_logic;
signal \U712_CHIP_RAM.N_335\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.un1_REGENn_0_sqmuxa_0_0_0\ : std_logic;
signal \N_165_i\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \RASn_c\ : std_logic;
signal \WEn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_314_cascade_\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA25_0_i\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_190\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\ : std_logic;
signal \U712_CYCLE_TERM.N_332\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.N_455_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_1\ : std_logic;
signal \U712_REG_SM.START_RSTZ0\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.N_361\ : std_logic;
signal \U712_CHIP_RAM.N_367\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \A_c_9\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_314\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.m50_i_a2_0_0\ : std_logic;
signal \N_200_i\ : std_logic;
signal \U712_CHIP_RAM.N_337\ : std_logic;
signal \CLK40_PLL_i\ : std_logic;
signal \CLK40_PLL_i_i\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_i_0_9\ : std_logic;
signal \A_c_19\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA25_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_0\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_2\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \N_334_cascade_\ : std_logic;
signal \N_177_i\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0\ : std_logic;
signal \N_336_cascade_\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \N_175_i\ : std_logic;
signal \N_337_i\ : std_logic;
signal \N_336_i\ : std_logic;
signal \N_335_i\ : std_logic;
signal \A_c_1\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \N_334_i\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \RnW_c\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \DMA_WRITE_CYCLE\ : std_logic;
signal \N_379\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \DA_wire\ : std_logic_vector(2 downto 0);
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    TBIn <= \TBIn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    ASn <= \ASn_wire\;
    DA <= \DA_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    TCIn <= \TCIn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    \C3_wire\ <= C3;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL_i\,
            REFERENCECLK => \N__4330\,
            RESETB => \N__7834\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12710\,
            DIN => \N__12709\,
            DOUT => \N__12708\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12710\,
            PADOUT => \N__12709\,
            PADIN => \N__12708\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5815\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12701\,
            DIN => \N__12700\,
            DOUT => \N__12699\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12701\,
            PADOUT => \N__12700\,
            PADIN => \N__12699\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12692\,
            DIN => \N__12691\,
            DOUT => \N__12690\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12692\,
            PADOUT => \N__12691\,
            PADIN => \N__12690\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8452\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12683\,
            DIN => \N__12682\,
            DOUT => \N__12681\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12683\,
            PADOUT => \N__12682\,
            PADIN => \N__12681\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11722\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12674\,
            DIN => \N__12673\,
            DOUT => \N__12672\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12674\,
            PADOUT => \N__12673\,
            PADIN => \N__12672\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12665\,
            DIN => \N__12664\,
            DOUT => \N__12663\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12665\,
            PADOUT => \N__12664\,
            PADIN => \N__12663\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12656\,
            DIN => \N__12655\,
            DOUT => \N__12654\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12656\,
            PADOUT => \N__12655\,
            PADIN => \N__12654\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12647\,
            DIN => \N__12646\,
            DOUT => \N__12645\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12647\,
            PADOUT => \N__12646\,
            PADIN => \N__12645\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12638\,
            DIN => \N__12637\,
            DOUT => \N__12636\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12638\,
            PADOUT => \N__12637\,
            PADIN => \N__12636\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12629\,
            DIN => \N__12628\,
            DOUT => \N__12627\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12629\,
            PADOUT => \N__12628\,
            PADIN => \N__12627\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12620\,
            DIN => \N__12619\,
            DOUT => \N__12618\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12620\,
            PADOUT => \N__12619\,
            PADIN => \N__12618\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12611\,
            DIN => \N__12610\,
            DOUT => \N__12609\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12611\,
            PADOUT => \N__12610\,
            PADIN => \N__12609\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9046\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12602\,
            DIN => \N__12601\,
            DOUT => \N__12600\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12602\,
            PADOUT => \N__12601\,
            PADIN => \N__12600\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11473\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12593\,
            DIN => \N__12592\,
            DOUT => \N__12591\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12593\,
            PADOUT => \N__12592\,
            PADIN => \N__12591\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12584\,
            DIN => \N__12583\,
            DOUT => \N__12582\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12584\,
            PADOUT => \N__12583\,
            PADIN => \N__12582\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12575\,
            DIN => \N__12574\,
            DOUT => \N__12573\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12575\,
            PADOUT => \N__12574\,
            PADIN => \N__12573\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12566\,
            DIN => \N__12565\,
            DOUT => \N__12564\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12566\,
            PADOUT => \N__12565\,
            PADIN => \N__12564\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4627\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12557\,
            DIN => \N__12556\,
            DOUT => \N__12555\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12557\,
            PADOUT => \N__12556\,
            PADIN => \N__12555\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12548\,
            DIN => \N__12547\,
            DOUT => \N__12546\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12548\,
            PADOUT => \N__12547\,
            PADIN => \N__12546\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12539\,
            DIN => \N__12538\,
            DOUT => \N__12537\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12539\,
            PADOUT => \N__12538\,
            PADIN => \N__12537\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9070\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12530\,
            DIN => \N__12529\,
            DOUT => \N__12528\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12530\,
            PADOUT => \N__12529\,
            PADIN => \N__12528\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12521\,
            DIN => \N__12520\,
            DOUT => \N__12519\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12521\,
            PADOUT => \N__12520\,
            PADIN => \N__12519\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9541\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12512\,
            DIN => \N__12511\,
            DOUT => \N__12510\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12512\,
            PADOUT => \N__12511\,
            PADIN => \N__12510\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12503\,
            DIN => \N__12502\,
            DOUT => \N__12501\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12503\,
            PADOUT => \N__12502\,
            PADIN => \N__12501\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11461\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12494\,
            DIN => \N__12493\,
            DOUT => \N__12492\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12494\,
            PADOUT => \N__12493\,
            PADIN => \N__12492\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7749\,
            DIN0 => OPEN,
            DOUT0 => \N__6113\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12485\,
            DIN => \N__12484\,
            DOUT => \N__12483\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12485\,
            PADOUT => \N__12484\,
            PADIN => \N__12483\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12476\,
            DIN => \N__12475\,
            DOUT => \N__12474\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12476\,
            PADOUT => \N__12475\,
            PADIN => \N__12474\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12467\,
            DIN => \N__12466\,
            DOUT => \N__12465\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12467\,
            PADOUT => \N__12466\,
            PADIN => \N__12465\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12458\,
            DIN => \N__12457\,
            DOUT => \N__12456\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12458\,
            PADOUT => \N__12457\,
            PADIN => \N__12456\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12449\,
            DIN => \N__12448\,
            DOUT => \N__12447\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12449\,
            PADOUT => \N__12448\,
            PADIN => \N__12447\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12440\,
            DIN => \N__12439\,
            DOUT => \N__12438\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12440\,
            PADOUT => \N__12439\,
            PADIN => \N__12438\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7852\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12431\,
            DIN => \N__12430\,
            DOUT => \N__12429\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12431\,
            PADOUT => \N__12430\,
            PADIN => \N__12429\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12422\,
            DIN => \N__12421\,
            DOUT => \N__12420\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12422\,
            PADOUT => \N__12421\,
            PADIN => \N__12420\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12413\,
            DIN => \N__12412\,
            DOUT => \N__12411\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12413\,
            PADOUT => \N__12412\,
            PADIN => \N__12411\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12404\,
            DIN => \N__12403\,
            DOUT => \N__12402\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12404\,
            PADOUT => \N__12403\,
            PADIN => \N__12402\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12395\,
            DIN => \N__12394\,
            DOUT => \N__12393\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12395\,
            PADOUT => \N__12394\,
            PADIN => \N__12393\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12386\,
            DIN => \N__12385\,
            DOUT => \N__12384\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12386\,
            PADOUT => \N__12385\,
            PADIN => \N__12384\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7810\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12377\,
            DIN => \N__12376\,
            DOUT => \N__12375\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12377\,
            PADOUT => \N__12376\,
            PADIN => \N__12375\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12368\,
            DIN => \N__12367\,
            DOUT => \N__12366\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12368\,
            PADOUT => \N__12367\,
            PADIN => \N__12366\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12359\,
            DIN => \N__12358\,
            DOUT => \N__12357\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12359\,
            PADOUT => \N__12358\,
            PADIN => \N__12357\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7879\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12350\,
            DIN => \N__12349\,
            DOUT => \N__12348\,
            PACKAGEPIN => \DA_wire\(0)
        );

    \DA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12350\,
            PADOUT => \N__12349\,
            PADIN => \N__12348\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9025\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12341\,
            DIN => \N__12340\,
            DOUT => \N__12339\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12341\,
            PADOUT => \N__12340\,
            PADIN => \N__12339\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12332\,
            DIN => \N__12331\,
            DOUT => \N__12330\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12332\,
            PADOUT => \N__12331\,
            PADIN => \N__12330\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8404\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12323\,
            DIN => \N__12322\,
            DOUT => \N__12321\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12323\,
            PADOUT => \N__12322\,
            PADIN => \N__12321\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8329\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12314\,
            DIN => \N__12313\,
            DOUT => \N__12312\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12314\,
            PADOUT => \N__12313\,
            PADIN => \N__12312\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5227\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12305\,
            DIN => \N__12304\,
            DOUT => \N__12303\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12305\,
            PADOUT => \N__12304\,
            PADIN => \N__12303\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12296\,
            DIN => \N__12295\,
            DOUT => \N__12294\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12296\,
            PADOUT => \N__12295\,
            PADIN => \N__12294\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12287\,
            DIN => \N__12286\,
            DOUT => \N__12285\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12287\,
            PADOUT => \N__12286\,
            PADIN => \N__12285\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9238\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12278\,
            DIN => \N__12277\,
            DOUT => \N__12276\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12278\,
            PADOUT => \N__12277\,
            PADIN => \N__12276\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7750\,
            DIN0 => OPEN,
            DOUT0 => \N__6127\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12269\,
            DIN => \N__12268\,
            DOUT => \N__12267\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12269\,
            PADOUT => \N__12268\,
            PADIN => \N__12267\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7789\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12260\,
            DIN => \N__12259\,
            DOUT => \N__12258\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12260\,
            PADOUT => \N__12259\,
            PADIN => \N__12258\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5077\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12251\,
            DIN => \N__12250\,
            DOUT => \N__12249\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12251\,
            PADOUT => \N__12250\,
            PADIN => \N__12249\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9736\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12242\,
            DIN => \N__12241\,
            DOUT => \N__12240\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12242\,
            PADOUT => \N__12241\,
            PADIN => \N__12240\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12233\,
            DIN => \N__12232\,
            DOUT => \N__12231\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12233\,
            PADOUT => \N__12232\,
            PADIN => \N__12231\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12224\,
            DIN => \N__12223\,
            DOUT => \N__12222\,
            PACKAGEPIN => \DA_wire\(2)
        );

    \DA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12224\,
            PADOUT => \N__12223\,
            PADIN => \N__12222\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6532\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12215\,
            DIN => \N__12214\,
            DOUT => \N__12213\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12215\,
            PADOUT => \N__12214\,
            PADIN => \N__12213\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12206\,
            DIN => \N__12205\,
            DOUT => \N__12204\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12206\,
            PADOUT => \N__12205\,
            PADIN => \N__12204\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12197\,
            DIN => \N__12196\,
            DOUT => \N__12195\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12197\,
            PADOUT => \N__12196\,
            PADIN => \N__12195\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8365\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12188\,
            DIN => \N__12187\,
            DOUT => \N__12186\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12188\,
            PADOUT => \N__12187\,
            PADIN => \N__12186\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11488\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12179\,
            DIN => \N__12178\,
            DOUT => \N__12177\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12179\,
            PADOUT => \N__12178\,
            PADIN => \N__12177\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12170\,
            DIN => \N__12169\,
            DOUT => \N__12168\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12170\,
            PADOUT => \N__12169\,
            PADIN => \N__12168\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11509\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12161\,
            DIN => \N__12160\,
            DOUT => \N__12159\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12161\,
            PADOUT => \N__12160\,
            PADIN => \N__12159\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7742\,
            DIN0 => OPEN,
            DOUT0 => \N__6123\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12152\,
            DIN => \N__12151\,
            DOUT => \N__12150\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12152\,
            PADOUT => \N__12151\,
            PADIN => \N__12150\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8704\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12143\,
            DIN => \N__12142\,
            DOUT => \N__12141\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12143\,
            PADOUT => \N__12142\,
            PADIN => \N__12141\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12134\,
            DIN => \N__12133\,
            DOUT => \N__12132\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12134\,
            PADOUT => \N__12133\,
            PADIN => \N__12132\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12125\,
            DIN => \N__12124\,
            DOUT => \N__12123\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12125\,
            PADOUT => \N__12124\,
            PADIN => \N__12123\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9094\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12116\,
            DIN => \N__12115\,
            DOUT => \N__12114\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12116\,
            PADOUT => \N__12115\,
            PADIN => \N__12114\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12107\,
            DIN => \N__12106\,
            DOUT => \N__12105\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12107\,
            PADOUT => \N__12106\,
            PADIN => \N__12105\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12098\,
            DIN => \N__12097\,
            DOUT => \N__12096\,
            PACKAGEPIN => \DA_wire\(1)
        );

    \DA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12098\,
            PADOUT => \N__12097\,
            PADIN => \N__12096\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6292\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12089\,
            DIN => \N__12088\,
            DOUT => \N__12087\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12089\,
            PADOUT => \N__12088\,
            PADIN => \N__12087\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12080\,
            DIN => \N__12079\,
            DOUT => \N__12078\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12080\,
            PADOUT => \N__12079\,
            PADIN => \N__12078\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12071\,
            DIN => \N__12070\,
            DOUT => \N__12069\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12071\,
            PADOUT => \N__12070\,
            PADIN => \N__12069\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8425\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12062\,
            DIN => \N__12061\,
            DOUT => \N__12060\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12062\,
            PADOUT => \N__12061\,
            PADIN => \N__12060\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5977\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12053\,
            DIN => \N__12052\,
            DOUT => \N__12051\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12053\,
            PADOUT => \N__12052\,
            PADIN => \N__12051\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11029\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12044\,
            DIN => \N__12043\,
            DOUT => \N__12042\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12044\,
            PADOUT => \N__12043\,
            PADIN => \N__12042\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5116\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12035\,
            DIN => \N__12034\,
            DOUT => \N__12033\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12035\,
            PADOUT => \N__12034\,
            PADIN => \N__12033\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12026\,
            DIN => \N__12025\,
            DOUT => \N__12024\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12026\,
            PADOUT => \N__12025\,
            PADIN => \N__12024\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12017\,
            DIN => \N__12016\,
            DOUT => \N__12015\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12017\,
            PADOUT => \N__12016\,
            PADIN => \N__12015\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8302\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12008\,
            DIN => \N__12007\,
            DOUT => \N__12006\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12008\,
            PADOUT => \N__12007\,
            PADIN => \N__12006\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11999\,
            DIN => \N__11998\,
            DOUT => \N__11997\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11999\,
            PADOUT => \N__11998\,
            PADIN => \N__11997\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11990\,
            DIN => \N__11989\,
            DOUT => \N__11988\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11990\,
            PADOUT => \N__11989\,
            PADIN => \N__11988\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5626\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11981\,
            DIN => \N__11980\,
            DOUT => \N__11979\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11981\,
            PADOUT => \N__11980\,
            PADIN => \N__11979\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6058\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11972\,
            DIN => \N__11971\,
            DOUT => \N__11970\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11972\,
            PADOUT => \N__11971\,
            PADIN => \N__11970\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9151\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11963\,
            DIN => \N__11962\,
            DOUT => \N__11961\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11963\,
            PADOUT => \N__11962\,
            PADIN => \N__11961\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11954\,
            DIN => \N__11953\,
            DOUT => \N__11952\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11954\,
            PADOUT => \N__11953\,
            PADIN => \N__11952\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9147\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11945\,
            DIN => \N__11944\,
            DOUT => \N__11943\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11945\,
            PADOUT => \N__11944\,
            PADIN => \N__11943\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4420\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11936\,
            DIN => \N__11935\,
            DOUT => \N__11934\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11936\,
            PADOUT => \N__11935\,
            PADIN => \N__11934\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8353\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11927\,
            DIN => \N__11926\,
            DOUT => \N__11925\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11927\,
            PADOUT => \N__11926\,
            PADIN => \N__11925\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11918\,
            DIN => \N__11917\,
            DOUT => \N__11916\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11918\,
            PADOUT => \N__11917\,
            PADIN => \N__11916\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11909\,
            DIN => \N__11908\,
            DOUT => \N__11907\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11909\,
            PADOUT => \N__11908\,
            PADIN => \N__11907\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11900\,
            DIN => \N__11899\,
            DOUT => \N__11898\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11900\,
            PADOUT => \N__11899\,
            PADIN => \N__11898\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11891\,
            DIN => \N__11890\,
            DOUT => \N__11889\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11891\,
            PADOUT => \N__11890\,
            PADIN => \N__11889\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9146\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11882\,
            DIN => \N__11881\,
            DOUT => \N__11880\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11882\,
            PADOUT => \N__11881\,
            PADIN => \N__11880\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7411\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11873\,
            DIN => \N__11872\,
            DOUT => \N__11871\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11873\,
            PADOUT => \N__11872\,
            PADIN => \N__11871\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6634\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11864\,
            DIN => \N__11863\,
            DOUT => \N__11862\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11864\,
            PADOUT => \N__11863\,
            PADIN => \N__11862\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9481\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2884\ : InMux
    port map (
            O => \N__11845\,
            I => \N__11842\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__11842\,
            I => \N__11837\
        );

    \I__2882\ : CascadeMux
    port map (
            O => \N__11841\,
            I => \N__11832\
        );

    \I__2881\ : CascadeMux
    port map (
            O => \N__11840\,
            I => \N__11828\
        );

    \I__2880\ : Span4Mux_h
    port map (
            O => \N__11837\,
            I => \N__11825\
        );

    \I__2879\ : InMux
    port map (
            O => \N__11836\,
            I => \N__11822\
        );

    \I__2878\ : InMux
    port map (
            O => \N__11835\,
            I => \N__11819\
        );

    \I__2877\ : InMux
    port map (
            O => \N__11832\,
            I => \N__11816\
        );

    \I__2876\ : InMux
    port map (
            O => \N__11831\,
            I => \N__11813\
        );

    \I__2875\ : InMux
    port map (
            O => \N__11828\,
            I => \N__11810\
        );

    \I__2874\ : Sp12to4
    port map (
            O => \N__11825\,
            I => \N__11805\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__11822\,
            I => \N__11805\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__11819\,
            I => \N__11800\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__11816\,
            I => \N__11800\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__11813\,
            I => \N__11797\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__11810\,
            I => \N__11794\
        );

    \I__2868\ : Span12Mux_v
    port map (
            O => \N__11805\,
            I => \N__11791\
        );

    \I__2867\ : Span12Mux_h
    port map (
            O => \N__11800\,
            I => \N__11788\
        );

    \I__2866\ : Span12Mux_v
    port map (
            O => \N__11797\,
            I => \N__11785\
        );

    \I__2865\ : Span4Mux_h
    port map (
            O => \N__11794\,
            I => \N__11782\
        );

    \I__2864\ : Span12Mux_h
    port map (
            O => \N__11791\,
            I => \N__11779\
        );

    \I__2863\ : Span12Mux_v
    port map (
            O => \N__11788\,
            I => \N__11774\
        );

    \I__2862\ : Span12Mux_h
    port map (
            O => \N__11785\,
            I => \N__11774\
        );

    \I__2861\ : Span4Mux_v
    port map (
            O => \N__11782\,
            I => \N__11771\
        );

    \I__2860\ : Odrv12
    port map (
            O => \N__11779\,
            I => \CASUn_c\
        );

    \I__2859\ : Odrv12
    port map (
            O => \N__11774\,
            I => \CASUn_c\
        );

    \I__2858\ : Odrv4
    port map (
            O => \N__11771\,
            I => \CASUn_c\
        );

    \I__2857\ : InMux
    port map (
            O => \N__11764\,
            I => \N__11761\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__11761\,
            I => \N__11758\
        );

    \I__2855\ : Span4Mux_v
    port map (
            O => \N__11758\,
            I => \N__11754\
        );

    \I__2854\ : InMux
    port map (
            O => \N__11757\,
            I => \N__11751\
        );

    \I__2853\ : Span4Mux_h
    port map (
            O => \N__11754\,
            I => \N__11748\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__11751\,
            I => \N__11745\
        );

    \I__2851\ : Sp12to4
    port map (
            O => \N__11748\,
            I => \N__11742\
        );

    \I__2850\ : Span4Mux_v
    port map (
            O => \N__11745\,
            I => \N__11739\
        );

    \I__2849\ : Span12Mux_h
    port map (
            O => \N__11742\,
            I => \N__11735\
        );

    \I__2848\ : Span4Mux_v
    port map (
            O => \N__11739\,
            I => \N__11732\
        );

    \I__2847\ : InMux
    port map (
            O => \N__11738\,
            I => \N__11729\
        );

    \I__2846\ : Odrv12
    port map (
            O => \N__11735\,
            I => \DMA_WRITE_CYCLE\
        );

    \I__2845\ : Odrv4
    port map (
            O => \N__11732\,
            I => \DMA_WRITE_CYCLE\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__11729\,
            I => \DMA_WRITE_CYCLE\
        );

    \I__2843\ : IoInMux
    port map (
            O => \N__11722\,
            I => \N__11719\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__11719\,
            I => \N__11716\
        );

    \I__2841\ : Span4Mux_s3_h
    port map (
            O => \N__11716\,
            I => \N__11713\
        );

    \I__2840\ : Span4Mux_v
    port map (
            O => \N__11713\,
            I => \N__11710\
        );

    \I__2839\ : Odrv4
    port map (
            O => \N__11710\,
            I => \N_379\
        );

    \I__2838\ : InMux
    port map (
            O => \N__11707\,
            I => \N__11704\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__11704\,
            I => \N__11700\
        );

    \I__2836\ : InMux
    port map (
            O => \N__11703\,
            I => \N__11697\
        );

    \I__2835\ : Span4Mux_v
    port map (
            O => \N__11700\,
            I => \N__11694\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__11697\,
            I => \N__11691\
        );

    \I__2833\ : Span4Mux_h
    port map (
            O => \N__11694\,
            I => \N__11688\
        );

    \I__2832\ : Span4Mux_v
    port map (
            O => \N__11691\,
            I => \N__11685\
        );

    \I__2831\ : Odrv4
    port map (
            O => \N__11688\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0\
        );

    \I__2830\ : Odrv4
    port map (
            O => \N__11685\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0\
        );

    \I__2829\ : CascadeMux
    port map (
            O => \N__11680\,
            I => \N_336_cascade_\
        );

    \I__2828\ : CascadeMux
    port map (
            O => \N__11677\,
            I => \N__11672\
        );

    \I__2827\ : InMux
    port map (
            O => \N__11676\,
            I => \N__11668\
        );

    \I__2826\ : InMux
    port map (
            O => \N__11675\,
            I => \N__11665\
        );

    \I__2825\ : InMux
    port map (
            O => \N__11672\,
            I => \N__11662\
        );

    \I__2824\ : InMux
    port map (
            O => \N__11671\,
            I => \N__11650\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__11668\,
            I => \N__11643\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__11665\,
            I => \N__11640\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__11662\,
            I => \N__11637\
        );

    \I__2820\ : InMux
    port map (
            O => \N__11661\,
            I => \N__11630\
        );

    \I__2819\ : InMux
    port map (
            O => \N__11660\,
            I => \N__11630\
        );

    \I__2818\ : InMux
    port map (
            O => \N__11659\,
            I => \N__11630\
        );

    \I__2817\ : InMux
    port map (
            O => \N__11658\,
            I => \N__11625\
        );

    \I__2816\ : InMux
    port map (
            O => \N__11657\,
            I => \N__11625\
        );

    \I__2815\ : InMux
    port map (
            O => \N__11656\,
            I => \N__11618\
        );

    \I__2814\ : InMux
    port map (
            O => \N__11655\,
            I => \N__11618\
        );

    \I__2813\ : InMux
    port map (
            O => \N__11654\,
            I => \N__11618\
        );

    \I__2812\ : InMux
    port map (
            O => \N__11653\,
            I => \N__11615\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__11650\,
            I => \N__11612\
        );

    \I__2810\ : InMux
    port map (
            O => \N__11649\,
            I => \N__11607\
        );

    \I__2809\ : InMux
    port map (
            O => \N__11648\,
            I => \N__11601\
        );

    \I__2808\ : InMux
    port map (
            O => \N__11647\,
            I => \N__11601\
        );

    \I__2807\ : InMux
    port map (
            O => \N__11646\,
            I => \N__11598\
        );

    \I__2806\ : Span4Mux_v
    port map (
            O => \N__11643\,
            I => \N__11587\
        );

    \I__2805\ : Span4Mux_v
    port map (
            O => \N__11640\,
            I => \N__11587\
        );

    \I__2804\ : Span4Mux_h
    port map (
            O => \N__11637\,
            I => \N__11587\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__11630\,
            I => \N__11587\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__11625\,
            I => \N__11587\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__11618\,
            I => \N__11584\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__11615\,
            I => \N__11581\
        );

    \I__2799\ : Span4Mux_v
    port map (
            O => \N__11612\,
            I => \N__11577\
        );

    \I__2798\ : InMux
    port map (
            O => \N__11611\,
            I => \N__11574\
        );

    \I__2797\ : InMux
    port map (
            O => \N__11610\,
            I => \N__11569\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__11607\,
            I => \N__11565\
        );

    \I__2795\ : InMux
    port map (
            O => \N__11606\,
            I => \N__11562\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__11601\,
            I => \N__11553\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__11598\,
            I => \N__11553\
        );

    \I__2792\ : Span4Mux_h
    port map (
            O => \N__11587\,
            I => \N__11553\
        );

    \I__2791\ : Span4Mux_v
    port map (
            O => \N__11584\,
            I => \N__11553\
        );

    \I__2790\ : Span4Mux_v
    port map (
            O => \N__11581\,
            I => \N__11550\
        );

    \I__2789\ : InMux
    port map (
            O => \N__11580\,
            I => \N__11547\
        );

    \I__2788\ : Span4Mux_h
    port map (
            O => \N__11577\,
            I => \N__11542\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__11574\,
            I => \N__11542\
        );

    \I__2786\ : InMux
    port map (
            O => \N__11573\,
            I => \N__11537\
        );

    \I__2785\ : InMux
    port map (
            O => \N__11572\,
            I => \N__11537\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__11569\,
            I => \N__11534\
        );

    \I__2783\ : InMux
    port map (
            O => \N__11568\,
            I => \N__11531\
        );

    \I__2782\ : Span4Mux_v
    port map (
            O => \N__11565\,
            I => \N__11524\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__11562\,
            I => \N__11524\
        );

    \I__2780\ : Span4Mux_v
    port map (
            O => \N__11553\,
            I => \N__11524\
        );

    \I__2779\ : Odrv4
    port map (
            O => \N__11550\,
            I => \CPU_CYCLEm\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__11547\,
            I => \CPU_CYCLEm\
        );

    \I__2777\ : Odrv4
    port map (
            O => \N__11542\,
            I => \CPU_CYCLEm\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__11537\,
            I => \CPU_CYCLEm\
        );

    \I__2775\ : Odrv12
    port map (
            O => \N__11534\,
            I => \CPU_CYCLEm\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__11531\,
            I => \CPU_CYCLEm\
        );

    \I__2773\ : Odrv4
    port map (
            O => \N__11524\,
            I => \CPU_CYCLEm\
        );

    \I__2772\ : IoInMux
    port map (
            O => \N__11509\,
            I => \N__11506\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__11506\,
            I => \N__11503\
        );

    \I__2770\ : Span4Mux_s2_h
    port map (
            O => \N__11503\,
            I => \N__11500\
        );

    \I__2769\ : Span4Mux_v
    port map (
            O => \N__11500\,
            I => \N__11497\
        );

    \I__2768\ : Sp12to4
    port map (
            O => \N__11497\,
            I => \N__11494\
        );

    \I__2767\ : Span12Mux_h
    port map (
            O => \N__11494\,
            I => \N__11491\
        );

    \I__2766\ : Odrv12
    port map (
            O => \N__11491\,
            I => \N_175_i\
        );

    \I__2765\ : IoInMux
    port map (
            O => \N__11488\,
            I => \N__11485\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__11485\,
            I => \N__11482\
        );

    \I__2763\ : IoSpan4Mux
    port map (
            O => \N__11482\,
            I => \N__11479\
        );

    \I__2762\ : Span4Mux_s3_v
    port map (
            O => \N__11479\,
            I => \N__11476\
        );

    \I__2761\ : Odrv4
    port map (
            O => \N__11476\,
            I => \N_337_i\
        );

    \I__2760\ : IoInMux
    port map (
            O => \N__11473\,
            I => \N__11470\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__11470\,
            I => \N__11467\
        );

    \I__2758\ : Span4Mux_s3_v
    port map (
            O => \N__11467\,
            I => \N__11464\
        );

    \I__2757\ : Odrv4
    port map (
            O => \N__11464\,
            I => \N_336_i\
        );

    \I__2756\ : IoInMux
    port map (
            O => \N__11461\,
            I => \N__11458\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__11458\,
            I => \N__11455\
        );

    \I__2754\ : Span12Mux_s6_v
    port map (
            O => \N__11455\,
            I => \N__11452\
        );

    \I__2753\ : Odrv12
    port map (
            O => \N__11452\,
            I => \N_335_i\
        );

    \I__2752\ : InMux
    port map (
            O => \N__11449\,
            I => \N__11444\
        );

    \I__2751\ : InMux
    port map (
            O => \N__11448\,
            I => \N__11441\
        );

    \I__2750\ : InMux
    port map (
            O => \N__11447\,
            I => \N__11438\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__11444\,
            I => \N__11431\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__11441\,
            I => \N__11427\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__11438\,
            I => \N__11424\
        );

    \I__2746\ : InMux
    port map (
            O => \N__11437\,
            I => \N__11415\
        );

    \I__2745\ : InMux
    port map (
            O => \N__11436\,
            I => \N__11415\
        );

    \I__2744\ : InMux
    port map (
            O => \N__11435\,
            I => \N__11415\
        );

    \I__2743\ : InMux
    port map (
            O => \N__11434\,
            I => \N__11415\
        );

    \I__2742\ : Span4Mux_v
    port map (
            O => \N__11431\,
            I => \N__11412\
        );

    \I__2741\ : InMux
    port map (
            O => \N__11430\,
            I => \N__11409\
        );

    \I__2740\ : Span4Mux_v
    port map (
            O => \N__11427\,
            I => \N__11406\
        );

    \I__2739\ : Span4Mux_v
    port map (
            O => \N__11424\,
            I => \N__11403\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__11415\,
            I => \N__11400\
        );

    \I__2737\ : Span4Mux_v
    port map (
            O => \N__11412\,
            I => \N__11397\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__11409\,
            I => \N__11394\
        );

    \I__2735\ : Span4Mux_v
    port map (
            O => \N__11406\,
            I => \N__11387\
        );

    \I__2734\ : Span4Mux_v
    port map (
            O => \N__11403\,
            I => \N__11387\
        );

    \I__2733\ : Span4Mux_v
    port map (
            O => \N__11400\,
            I => \N__11387\
        );

    \I__2732\ : Sp12to4
    port map (
            O => \N__11397\,
            I => \N__11382\
        );

    \I__2731\ : Span12Mux_v
    port map (
            O => \N__11394\,
            I => \N__11382\
        );

    \I__2730\ : Sp12to4
    port map (
            O => \N__11387\,
            I => \N__11379\
        );

    \I__2729\ : Span12Mux_h
    port map (
            O => \N__11382\,
            I => \N__11376\
        );

    \I__2728\ : Span12Mux_h
    port map (
            O => \N__11379\,
            I => \N__11373\
        );

    \I__2727\ : Odrv12
    port map (
            O => \N__11376\,
            I => \A_c_1\
        );

    \I__2726\ : Odrv12
    port map (
            O => \N__11373\,
            I => \A_c_1\
        );

    \I__2725\ : InMux
    port map (
            O => \N__11368\,
            I => \N__11353\
        );

    \I__2724\ : InMux
    port map (
            O => \N__11367\,
            I => \N__11353\
        );

    \I__2723\ : InMux
    port map (
            O => \N__11366\,
            I => \N__11353\
        );

    \I__2722\ : InMux
    port map (
            O => \N__11365\,
            I => \N__11353\
        );

    \I__2721\ : InMux
    port map (
            O => \N__11364\,
            I => \N__11350\
        );

    \I__2720\ : InMux
    port map (
            O => \N__11363\,
            I => \N__11346\
        );

    \I__2719\ : CascadeMux
    port map (
            O => \N__11362\,
            I => \N__11343\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__11353\,
            I => \N__11339\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__11350\,
            I => \N__11336\
        );

    \I__2716\ : InMux
    port map (
            O => \N__11349\,
            I => \N__11333\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__11346\,
            I => \N__11329\
        );

    \I__2714\ : InMux
    port map (
            O => \N__11343\,
            I => \N__11326\
        );

    \I__2713\ : InMux
    port map (
            O => \N__11342\,
            I => \N__11323\
        );

    \I__2712\ : Span4Mux_v
    port map (
            O => \N__11339\,
            I => \N__11318\
        );

    \I__2711\ : Span4Mux_v
    port map (
            O => \N__11336\,
            I => \N__11318\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__11333\,
            I => \N__11315\
        );

    \I__2709\ : InMux
    port map (
            O => \N__11332\,
            I => \N__11312\
        );

    \I__2708\ : Span4Mux_v
    port map (
            O => \N__11329\,
            I => \N__11309\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__11326\,
            I => \N__11306\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__11323\,
            I => \N__11303\
        );

    \I__2705\ : Span4Mux_h
    port map (
            O => \N__11318\,
            I => \N__11298\
        );

    \I__2704\ : Span4Mux_v
    port map (
            O => \N__11315\,
            I => \N__11298\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__11312\,
            I => \N__11295\
        );

    \I__2702\ : Sp12to4
    port map (
            O => \N__11309\,
            I => \N__11290\
        );

    \I__2701\ : Span12Mux_v
    port map (
            O => \N__11306\,
            I => \N__11290\
        );

    \I__2700\ : Span4Mux_v
    port map (
            O => \N__11303\,
            I => \N__11287\
        );

    \I__2699\ : Span4Mux_h
    port map (
            O => \N__11298\,
            I => \N__11282\
        );

    \I__2698\ : Span4Mux_v
    port map (
            O => \N__11295\,
            I => \N__11282\
        );

    \I__2697\ : Span12Mux_h
    port map (
            O => \N__11290\,
            I => \N__11279\
        );

    \I__2696\ : Sp12to4
    port map (
            O => \N__11287\,
            I => \N__11274\
        );

    \I__2695\ : Sp12to4
    port map (
            O => \N__11282\,
            I => \N__11274\
        );

    \I__2694\ : Odrv12
    port map (
            O => \N__11279\,
            I => \A_c_0\
        );

    \I__2693\ : Odrv12
    port map (
            O => \N__11274\,
            I => \A_c_0\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__11269\,
            I => \N__11266\
        );

    \I__2691\ : InMux
    port map (
            O => \N__11266\,
            I => \N__11259\
        );

    \I__2690\ : InMux
    port map (
            O => \N__11265\,
            I => \N__11256\
        );

    \I__2689\ : CascadeMux
    port map (
            O => \N__11264\,
            I => \N__11250\
        );

    \I__2688\ : CascadeMux
    port map (
            O => \N__11263\,
            I => \N__11247\
        );

    \I__2687\ : CascadeMux
    port map (
            O => \N__11262\,
            I => \N__11244\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__11259\,
            I => \N__11241\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__11256\,
            I => \N__11238\
        );

    \I__2684\ : InMux
    port map (
            O => \N__11255\,
            I => \N__11229\
        );

    \I__2683\ : InMux
    port map (
            O => \N__11254\,
            I => \N__11229\
        );

    \I__2682\ : InMux
    port map (
            O => \N__11253\,
            I => \N__11229\
        );

    \I__2681\ : InMux
    port map (
            O => \N__11250\,
            I => \N__11229\
        );

    \I__2680\ : InMux
    port map (
            O => \N__11247\,
            I => \N__11226\
        );

    \I__2679\ : InMux
    port map (
            O => \N__11244\,
            I => \N__11223\
        );

    \I__2678\ : Span4Mux_v
    port map (
            O => \N__11241\,
            I => \N__11218\
        );

    \I__2677\ : Span4Mux_v
    port map (
            O => \N__11238\,
            I => \N__11218\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__11229\,
            I => \N__11215\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__11226\,
            I => \N__11212\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__11223\,
            I => \N__11209\
        );

    \I__2673\ : Span4Mux_v
    port map (
            O => \N__11218\,
            I => \N__11202\
        );

    \I__2672\ : Span4Mux_h
    port map (
            O => \N__11215\,
            I => \N__11202\
        );

    \I__2671\ : Span4Mux_v
    port map (
            O => \N__11212\,
            I => \N__11199\
        );

    \I__2670\ : Span4Mux_v
    port map (
            O => \N__11209\,
            I => \N__11196\
        );

    \I__2669\ : InMux
    port map (
            O => \N__11208\,
            I => \N__11193\
        );

    \I__2668\ : InMux
    port map (
            O => \N__11207\,
            I => \N__11190\
        );

    \I__2667\ : Span4Mux_h
    port map (
            O => \N__11202\,
            I => \N__11185\
        );

    \I__2666\ : Span4Mux_v
    port map (
            O => \N__11199\,
            I => \N__11185\
        );

    \I__2665\ : Span4Mux_h
    port map (
            O => \N__11196\,
            I => \N__11180\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__11193\,
            I => \N__11180\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__11190\,
            I => \N__11177\
        );

    \I__2662\ : Span4Mux_v
    port map (
            O => \N__11185\,
            I => \N__11174\
        );

    \I__2661\ : Span4Mux_h
    port map (
            O => \N__11180\,
            I => \N__11171\
        );

    \I__2660\ : Span12Mux_v
    port map (
            O => \N__11177\,
            I => \N__11168\
        );

    \I__2659\ : Span4Mux_h
    port map (
            O => \N__11174\,
            I => \N__11165\
        );

    \I__2658\ : Sp12to4
    port map (
            O => \N__11171\,
            I => \N__11162\
        );

    \I__2657\ : Span12Mux_h
    port map (
            O => \N__11168\,
            I => \N__11159\
        );

    \I__2656\ : Sp12to4
    port map (
            O => \N__11165\,
            I => \N__11154\
        );

    \I__2655\ : Span12Mux_v
    port map (
            O => \N__11162\,
            I => \N__11154\
        );

    \I__2654\ : Odrv12
    port map (
            O => \N__11159\,
            I => \SIZ_c_1\
        );

    \I__2653\ : Odrv12
    port map (
            O => \N__11154\,
            I => \SIZ_c_1\
        );

    \I__2652\ : CascadeMux
    port map (
            O => \N__11149\,
            I => \N__11144\
        );

    \I__2651\ : InMux
    port map (
            O => \N__11148\,
            I => \N__11141\
        );

    \I__2650\ : InMux
    port map (
            O => \N__11147\,
            I => \N__11135\
        );

    \I__2649\ : InMux
    port map (
            O => \N__11144\,
            I => \N__11132\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__11141\,
            I => \N__11129\
        );

    \I__2647\ : CascadeMux
    port map (
            O => \N__11140\,
            I => \N__11126\
        );

    \I__2646\ : CascadeMux
    port map (
            O => \N__11139\,
            I => \N__11123\
        );

    \I__2645\ : CascadeMux
    port map (
            O => \N__11138\,
            I => \N__11120\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__11135\,
            I => \N__11116\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__11132\,
            I => \N__11113\
        );

    \I__2642\ : Span4Mux_v
    port map (
            O => \N__11129\,
            I => \N__11110\
        );

    \I__2641\ : InMux
    port map (
            O => \N__11126\,
            I => \N__11101\
        );

    \I__2640\ : InMux
    port map (
            O => \N__11123\,
            I => \N__11101\
        );

    \I__2639\ : InMux
    port map (
            O => \N__11120\,
            I => \N__11101\
        );

    \I__2638\ : InMux
    port map (
            O => \N__11119\,
            I => \N__11101\
        );

    \I__2637\ : Span4Mux_v
    port map (
            O => \N__11116\,
            I => \N__11097\
        );

    \I__2636\ : Span4Mux_v
    port map (
            O => \N__11113\,
            I => \N__11093\
        );

    \I__2635\ : Span4Mux_v
    port map (
            O => \N__11110\,
            I => \N__11088\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__11101\,
            I => \N__11088\
        );

    \I__2633\ : CascadeMux
    port map (
            O => \N__11100\,
            I => \N__11084\
        );

    \I__2632\ : Span4Mux_v
    port map (
            O => \N__11097\,
            I => \N__11081\
        );

    \I__2631\ : InMux
    port map (
            O => \N__11096\,
            I => \N__11078\
        );

    \I__2630\ : Span4Mux_v
    port map (
            O => \N__11093\,
            I => \N__11073\
        );

    \I__2629\ : Span4Mux_h
    port map (
            O => \N__11088\,
            I => \N__11073\
        );

    \I__2628\ : InMux
    port map (
            O => \N__11087\,
            I => \N__11070\
        );

    \I__2627\ : InMux
    port map (
            O => \N__11084\,
            I => \N__11067\
        );

    \I__2626\ : Span4Mux_v
    port map (
            O => \N__11081\,
            I => \N__11064\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__11078\,
            I => \N__11061\
        );

    \I__2624\ : Span4Mux_v
    port map (
            O => \N__11073\,
            I => \N__11058\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__11070\,
            I => \N__11053\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__11067\,
            I => \N__11053\
        );

    \I__2621\ : Sp12to4
    port map (
            O => \N__11064\,
            I => \N__11048\
        );

    \I__2620\ : Span12Mux_v
    port map (
            O => \N__11061\,
            I => \N__11048\
        );

    \I__2619\ : Span4Mux_h
    port map (
            O => \N__11058\,
            I => \N__11045\
        );

    \I__2618\ : Sp12to4
    port map (
            O => \N__11053\,
            I => \N__11042\
        );

    \I__2617\ : Span12Mux_h
    port map (
            O => \N__11048\,
            I => \N__11039\
        );

    \I__2616\ : Sp12to4
    port map (
            O => \N__11045\,
            I => \N__11034\
        );

    \I__2615\ : Span12Mux_v
    port map (
            O => \N__11042\,
            I => \N__11034\
        );

    \I__2614\ : Odrv12
    port map (
            O => \N__11039\,
            I => \SIZ_c_0\
        );

    \I__2613\ : Odrv12
    port map (
            O => \N__11034\,
            I => \SIZ_c_0\
        );

    \I__2612\ : IoInMux
    port map (
            O => \N__11029\,
            I => \N__11026\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__11026\,
            I => \N__11023\
        );

    \I__2610\ : Span4Mux_s2_v
    port map (
            O => \N__11023\,
            I => \N__11020\
        );

    \I__2609\ : Span4Mux_h
    port map (
            O => \N__11020\,
            I => \N__11017\
        );

    \I__2608\ : Span4Mux_v
    port map (
            O => \N__11017\,
            I => \N__11014\
        );

    \I__2607\ : Odrv4
    port map (
            O => \N__11014\,
            I => \N_334_i\
        );

    \I__2606\ : InMux
    port map (
            O => \N__11011\,
            I => \N__11007\
        );

    \I__2605\ : InMux
    port map (
            O => \N__11010\,
            I => \N__11003\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__11007\,
            I => \N__11000\
        );

    \I__2603\ : InMux
    port map (
            O => \N__11006\,
            I => \N__10997\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__11003\,
            I => \N__10989\
        );

    \I__2601\ : Span4Mux_h
    port map (
            O => \N__11000\,
            I => \N__10989\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__10997\,
            I => \N__10989\
        );

    \I__2599\ : InMux
    port map (
            O => \N__10996\,
            I => \N__10986\
        );

    \I__2598\ : Span4Mux_v
    port map (
            O => \N__10989\,
            I => \N__10983\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__10986\,
            I => \N__10980\
        );

    \I__2596\ : Span4Mux_v
    port map (
            O => \N__10983\,
            I => \N__10977\
        );

    \I__2595\ : Sp12to4
    port map (
            O => \N__10980\,
            I => \N__10974\
        );

    \I__2594\ : Sp12to4
    port map (
            O => \N__10977\,
            I => \N__10971\
        );

    \I__2593\ : Span12Mux_v
    port map (
            O => \N__10974\,
            I => \N__10968\
        );

    \I__2592\ : Span12Mux_h
    port map (
            O => \N__10971\,
            I => \N__10965\
        );

    \I__2591\ : Span12Mux_h
    port map (
            O => \N__10968\,
            I => \N__10962\
        );

    \I__2590\ : Odrv12
    port map (
            O => \N__10965\,
            I => \DRA_c_4\
        );

    \I__2589\ : Odrv12
    port map (
            O => \N__10962\,
            I => \DRA_c_4\
        );

    \I__2588\ : InMux
    port map (
            O => \N__10957\,
            I => \N__10951\
        );

    \I__2587\ : InMux
    port map (
            O => \N__10956\,
            I => \N__10951\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__10951\,
            I => \N__10946\
        );

    \I__2585\ : InMux
    port map (
            O => \N__10950\,
            I => \N__10943\
        );

    \I__2584\ : InMux
    port map (
            O => \N__10949\,
            I => \N__10940\
        );

    \I__2583\ : Span4Mux_h
    port map (
            O => \N__10946\,
            I => \N__10933\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__10943\,
            I => \N__10933\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__10940\,
            I => \N__10933\
        );

    \I__2580\ : Span4Mux_h
    port map (
            O => \N__10933\,
            I => \N__10930\
        );

    \I__2579\ : Sp12to4
    port map (
            O => \N__10930\,
            I => \N__10927\
        );

    \I__2578\ : Span12Mux_v
    port map (
            O => \N__10927\,
            I => \N__10924\
        );

    \I__2577\ : Odrv12
    port map (
            O => \N__10924\,
            I => \DRA_c_3\
        );

    \I__2576\ : InMux
    port map (
            O => \N__10921\,
            I => \N__10918\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__10918\,
            I => \N__10915\
        );

    \I__2574\ : Odrv12
    port map (
            O => \N__10915\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__2573\ : InMux
    port map (
            O => \N__10912\,
            I => \N__10908\
        );

    \I__2572\ : InMux
    port map (
            O => \N__10911\,
            I => \N__10905\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__10908\,
            I => \N__10899\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__10905\,
            I => \N__10899\
        );

    \I__2569\ : InMux
    port map (
            O => \N__10904\,
            I => \N__10896\
        );

    \I__2568\ : Span4Mux_v
    port map (
            O => \N__10899\,
            I => \N__10892\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__10896\,
            I => \N__10889\
        );

    \I__2566\ : InMux
    port map (
            O => \N__10895\,
            I => \N__10886\
        );

    \I__2565\ : Span4Mux_v
    port map (
            O => \N__10892\,
            I => \N__10883\
        );

    \I__2564\ : Sp12to4
    port map (
            O => \N__10889\,
            I => \N__10878\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__10886\,
            I => \N__10878\
        );

    \I__2562\ : Sp12to4
    port map (
            O => \N__10883\,
            I => \N__10873\
        );

    \I__2561\ : Span12Mux_v
    port map (
            O => \N__10878\,
            I => \N__10873\
        );

    \I__2560\ : Span12Mux_h
    port map (
            O => \N__10873\,
            I => \N__10870\
        );

    \I__2559\ : Odrv12
    port map (
            O => \N__10870\,
            I => \DRA_c_6\
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__10867\,
            I => \N__10864\
        );

    \I__2557\ : InMux
    port map (
            O => \N__10864\,
            I => \N__10858\
        );

    \I__2556\ : CascadeMux
    port map (
            O => \N__10863\,
            I => \N__10854\
        );

    \I__2555\ : InMux
    port map (
            O => \N__10862\,
            I => \N__10843\
        );

    \I__2554\ : InMux
    port map (
            O => \N__10861\,
            I => \N__10840\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__10858\,
            I => \N__10834\
        );

    \I__2552\ : InMux
    port map (
            O => \N__10857\,
            I => \N__10825\
        );

    \I__2551\ : InMux
    port map (
            O => \N__10854\,
            I => \N__10825\
        );

    \I__2550\ : InMux
    port map (
            O => \N__10853\,
            I => \N__10825\
        );

    \I__2549\ : InMux
    port map (
            O => \N__10852\,
            I => \N__10825\
        );

    \I__2548\ : InMux
    port map (
            O => \N__10851\,
            I => \N__10822\
        );

    \I__2547\ : InMux
    port map (
            O => \N__10850\,
            I => \N__10817\
        );

    \I__2546\ : InMux
    port map (
            O => \N__10849\,
            I => \N__10817\
        );

    \I__2545\ : InMux
    port map (
            O => \N__10848\,
            I => \N__10814\
        );

    \I__2544\ : InMux
    port map (
            O => \N__10847\,
            I => \N__10809\
        );

    \I__2543\ : InMux
    port map (
            O => \N__10846\,
            I => \N__10809\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__10843\,
            I => \N__10804\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__10840\,
            I => \N__10804\
        );

    \I__2540\ : InMux
    port map (
            O => \N__10839\,
            I => \N__10801\
        );

    \I__2539\ : InMux
    port map (
            O => \N__10838\,
            I => \N__10796\
        );

    \I__2538\ : InMux
    port map (
            O => \N__10837\,
            I => \N__10796\
        );

    \I__2537\ : Span4Mux_v
    port map (
            O => \N__10834\,
            I => \N__10792\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__10825\,
            I => \N__10781\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__10822\,
            I => \N__10781\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__10817\,
            I => \N__10781\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__10814\,
            I => \N__10781\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__10809\,
            I => \N__10781\
        );

    \I__2531\ : Span4Mux_v
    port map (
            O => \N__10804\,
            I => \N__10778\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__10801\,
            I => \N__10775\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__10796\,
            I => \N__10768\
        );

    \I__2528\ : InMux
    port map (
            O => \N__10795\,
            I => \N__10765\
        );

    \I__2527\ : Span4Mux_h
    port map (
            O => \N__10792\,
            I => \N__10760\
        );

    \I__2526\ : Span4Mux_v
    port map (
            O => \N__10781\,
            I => \N__10760\
        );

    \I__2525\ : Span4Mux_h
    port map (
            O => \N__10778\,
            I => \N__10755\
        );

    \I__2524\ : Span4Mux_v
    port map (
            O => \N__10775\,
            I => \N__10755\
        );

    \I__2523\ : InMux
    port map (
            O => \N__10774\,
            I => \N__10752\
        );

    \I__2522\ : InMux
    port map (
            O => \N__10773\,
            I => \N__10749\
        );

    \I__2521\ : InMux
    port map (
            O => \N__10772\,
            I => \N__10746\
        );

    \I__2520\ : InMux
    port map (
            O => \N__10771\,
            I => \N__10743\
        );

    \I__2519\ : Span4Mux_v
    port map (
            O => \N__10768\,
            I => \N__10738\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__10765\,
            I => \N__10738\
        );

    \I__2517\ : Sp12to4
    port map (
            O => \N__10760\,
            I => \N__10733\
        );

    \I__2516\ : Sp12to4
    port map (
            O => \N__10755\,
            I => \N__10733\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__10752\,
            I => \N__10728\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__10749\,
            I => \N__10728\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__10746\,
            I => \N__10723\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__10743\,
            I => \N__10723\
        );

    \I__2511\ : Sp12to4
    port map (
            O => \N__10738\,
            I => \N__10720\
        );

    \I__2510\ : Span12Mux_h
    port map (
            O => \N__10733\,
            I => \N__10717\
        );

    \I__2509\ : Span12Mux_h
    port map (
            O => \N__10728\,
            I => \N__10714\
        );

    \I__2508\ : Span12Mux_v
    port map (
            O => \N__10723\,
            I => \N__10711\
        );

    \I__2507\ : Span12Mux_v
    port map (
            O => \N__10720\,
            I => \N__10708\
        );

    \I__2506\ : Span12Mux_v
    port map (
            O => \N__10717\,
            I => \N__10705\
        );

    \I__2505\ : Span12Mux_v
    port map (
            O => \N__10714\,
            I => \N__10700\
        );

    \I__2504\ : Span12Mux_h
    port map (
            O => \N__10711\,
            I => \N__10700\
        );

    \I__2503\ : Span12Mux_h
    port map (
            O => \N__10708\,
            I => \N__10697\
        );

    \I__2502\ : Odrv12
    port map (
            O => \N__10705\,
            I => \AGNUS_REV_c\
        );

    \I__2501\ : Odrv12
    port map (
            O => \N__10700\,
            I => \AGNUS_REV_c\
        );

    \I__2500\ : Odrv12
    port map (
            O => \N__10697\,
            I => \AGNUS_REV_c\
        );

    \I__2499\ : InMux
    port map (
            O => \N__10690\,
            I => \N__10684\
        );

    \I__2498\ : InMux
    port map (
            O => \N__10689\,
            I => \N__10681\
        );

    \I__2497\ : InMux
    port map (
            O => \N__10688\,
            I => \N__10678\
        );

    \I__2496\ : InMux
    port map (
            O => \N__10687\,
            I => \N__10675\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__10684\,
            I => \N__10668\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__10681\,
            I => \N__10668\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__10678\,
            I => \N__10668\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__10675\,
            I => \N__10665\
        );

    \I__2491\ : Span4Mux_v
    port map (
            O => \N__10668\,
            I => \N__10662\
        );

    \I__2490\ : Span4Mux_v
    port map (
            O => \N__10665\,
            I => \N__10659\
        );

    \I__2489\ : Sp12to4
    port map (
            O => \N__10662\,
            I => \N__10656\
        );

    \I__2488\ : Span4Mux_h
    port map (
            O => \N__10659\,
            I => \N__10653\
        );

    \I__2487\ : Span12Mux_h
    port map (
            O => \N__10656\,
            I => \N__10648\
        );

    \I__2486\ : Sp12to4
    port map (
            O => \N__10653\,
            I => \N__10648\
        );

    \I__2485\ : Odrv12
    port map (
            O => \N__10648\,
            I => \DRA_c_7\
        );

    \I__2484\ : InMux
    port map (
            O => \N__10645\,
            I => \N__10642\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__10642\,
            I => \N__10639\
        );

    \I__2482\ : Span4Mux_h
    port map (
            O => \N__10639\,
            I => \N__10636\
        );

    \I__2481\ : Odrv4
    port map (
            O => \N__10636\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2480\ : ClkMux
    port map (
            O => \N__10633\,
            I => \N__10615\
        );

    \I__2479\ : ClkMux
    port map (
            O => \N__10632\,
            I => \N__10615\
        );

    \I__2478\ : ClkMux
    port map (
            O => \N__10631\,
            I => \N__10615\
        );

    \I__2477\ : ClkMux
    port map (
            O => \N__10630\,
            I => \N__10615\
        );

    \I__2476\ : ClkMux
    port map (
            O => \N__10629\,
            I => \N__10615\
        );

    \I__2475\ : ClkMux
    port map (
            O => \N__10628\,
            I => \N__10615\
        );

    \I__2474\ : GlobalMux
    port map (
            O => \N__10615\,
            I => \N__10612\
        );

    \I__2473\ : gio2CtrlBuf
    port map (
            O => \N__10612\,
            I => \C3_c_g\
        );

    \I__2472\ : CEMux
    port map (
            O => \N__10609\,
            I => \N__10573\
        );

    \I__2471\ : CEMux
    port map (
            O => \N__10608\,
            I => \N__10573\
        );

    \I__2470\ : CEMux
    port map (
            O => \N__10607\,
            I => \N__10573\
        );

    \I__2469\ : CEMux
    port map (
            O => \N__10606\,
            I => \N__10573\
        );

    \I__2468\ : CEMux
    port map (
            O => \N__10605\,
            I => \N__10573\
        );

    \I__2467\ : CEMux
    port map (
            O => \N__10604\,
            I => \N__10573\
        );

    \I__2466\ : CEMux
    port map (
            O => \N__10603\,
            I => \N__10573\
        );

    \I__2465\ : CEMux
    port map (
            O => \N__10602\,
            I => \N__10573\
        );

    \I__2464\ : CEMux
    port map (
            O => \N__10601\,
            I => \N__10573\
        );

    \I__2463\ : CEMux
    port map (
            O => \N__10600\,
            I => \N__10573\
        );

    \I__2462\ : CEMux
    port map (
            O => \N__10599\,
            I => \N__10573\
        );

    \I__2461\ : CEMux
    port map (
            O => \N__10598\,
            I => \N__10573\
        );

    \I__2460\ : GlobalMux
    port map (
            O => \N__10573\,
            I => \N__10570\
        );

    \I__2459\ : gio2CtrlBuf
    port map (
            O => \N__10570\,
            I => \DBRn_c_i_0_g\
        );

    \I__2458\ : InMux
    port map (
            O => \N__10567\,
            I => \N__10559\
        );

    \I__2457\ : InMux
    port map (
            O => \N__10566\,
            I => \N__10556\
        );

    \I__2456\ : InMux
    port map (
            O => \N__10565\,
            I => \N__10553\
        );

    \I__2455\ : InMux
    port map (
            O => \N__10564\,
            I => \N__10550\
        );

    \I__2454\ : InMux
    port map (
            O => \N__10563\,
            I => \N__10547\
        );

    \I__2453\ : InMux
    port map (
            O => \N__10562\,
            I => \N__10544\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__10559\,
            I => \N__10541\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__10556\,
            I => \N__10536\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__10553\,
            I => \N__10532\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__10550\,
            I => \N__10525\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__10547\,
            I => \N__10519\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__10544\,
            I => \N__10490\
        );

    \I__2446\ : Glb2LocalMux
    port map (
            O => \N__10541\,
            I => \N__10396\
        );

    \I__2445\ : SRMux
    port map (
            O => \N__10540\,
            I => \N__10396\
        );

    \I__2444\ : SRMux
    port map (
            O => \N__10539\,
            I => \N__10396\
        );

    \I__2443\ : Glb2LocalMux
    port map (
            O => \N__10536\,
            I => \N__10396\
        );

    \I__2442\ : SRMux
    port map (
            O => \N__10535\,
            I => \N__10396\
        );

    \I__2441\ : Glb2LocalMux
    port map (
            O => \N__10532\,
            I => \N__10396\
        );

    \I__2440\ : SRMux
    port map (
            O => \N__10531\,
            I => \N__10396\
        );

    \I__2439\ : SRMux
    port map (
            O => \N__10530\,
            I => \N__10396\
        );

    \I__2438\ : SRMux
    port map (
            O => \N__10529\,
            I => \N__10396\
        );

    \I__2437\ : SRMux
    port map (
            O => \N__10528\,
            I => \N__10396\
        );

    \I__2436\ : Glb2LocalMux
    port map (
            O => \N__10525\,
            I => \N__10396\
        );

    \I__2435\ : SRMux
    port map (
            O => \N__10524\,
            I => \N__10396\
        );

    \I__2434\ : SRMux
    port map (
            O => \N__10523\,
            I => \N__10396\
        );

    \I__2433\ : SRMux
    port map (
            O => \N__10522\,
            I => \N__10396\
        );

    \I__2432\ : Glb2LocalMux
    port map (
            O => \N__10519\,
            I => \N__10396\
        );

    \I__2431\ : SRMux
    port map (
            O => \N__10518\,
            I => \N__10396\
        );

    \I__2430\ : SRMux
    port map (
            O => \N__10517\,
            I => \N__10396\
        );

    \I__2429\ : SRMux
    port map (
            O => \N__10516\,
            I => \N__10396\
        );

    \I__2428\ : SRMux
    port map (
            O => \N__10515\,
            I => \N__10396\
        );

    \I__2427\ : SRMux
    port map (
            O => \N__10514\,
            I => \N__10396\
        );

    \I__2426\ : SRMux
    port map (
            O => \N__10513\,
            I => \N__10396\
        );

    \I__2425\ : SRMux
    port map (
            O => \N__10512\,
            I => \N__10396\
        );

    \I__2424\ : SRMux
    port map (
            O => \N__10511\,
            I => \N__10396\
        );

    \I__2423\ : SRMux
    port map (
            O => \N__10510\,
            I => \N__10396\
        );

    \I__2422\ : SRMux
    port map (
            O => \N__10509\,
            I => \N__10396\
        );

    \I__2421\ : SRMux
    port map (
            O => \N__10508\,
            I => \N__10396\
        );

    \I__2420\ : SRMux
    port map (
            O => \N__10507\,
            I => \N__10396\
        );

    \I__2419\ : SRMux
    port map (
            O => \N__10506\,
            I => \N__10396\
        );

    \I__2418\ : SRMux
    port map (
            O => \N__10505\,
            I => \N__10396\
        );

    \I__2417\ : SRMux
    port map (
            O => \N__10504\,
            I => \N__10396\
        );

    \I__2416\ : SRMux
    port map (
            O => \N__10503\,
            I => \N__10396\
        );

    \I__2415\ : SRMux
    port map (
            O => \N__10502\,
            I => \N__10396\
        );

    \I__2414\ : SRMux
    port map (
            O => \N__10501\,
            I => \N__10396\
        );

    \I__2413\ : SRMux
    port map (
            O => \N__10500\,
            I => \N__10396\
        );

    \I__2412\ : SRMux
    port map (
            O => \N__10499\,
            I => \N__10396\
        );

    \I__2411\ : SRMux
    port map (
            O => \N__10498\,
            I => \N__10396\
        );

    \I__2410\ : SRMux
    port map (
            O => \N__10497\,
            I => \N__10396\
        );

    \I__2409\ : SRMux
    port map (
            O => \N__10496\,
            I => \N__10396\
        );

    \I__2408\ : SRMux
    port map (
            O => \N__10495\,
            I => \N__10396\
        );

    \I__2407\ : SRMux
    port map (
            O => \N__10494\,
            I => \N__10396\
        );

    \I__2406\ : SRMux
    port map (
            O => \N__10493\,
            I => \N__10396\
        );

    \I__2405\ : Glb2LocalMux
    port map (
            O => \N__10490\,
            I => \N__10396\
        );

    \I__2404\ : SRMux
    port map (
            O => \N__10489\,
            I => \N__10396\
        );

    \I__2403\ : SRMux
    port map (
            O => \N__10488\,
            I => \N__10396\
        );

    \I__2402\ : SRMux
    port map (
            O => \N__10487\,
            I => \N__10396\
        );

    \I__2401\ : GlobalMux
    port map (
            O => \N__10396\,
            I => \N__10393\
        );

    \I__2400\ : gio2CtrlBuf
    port map (
            O => \N__10393\,
            I => \RESETn_c_i_g\
        );

    \I__2399\ : InMux
    port map (
            O => \N__10390\,
            I => \N__10386\
        );

    \I__2398\ : InMux
    port map (
            O => \N__10389\,
            I => \N__10381\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__10386\,
            I => \N__10377\
        );

    \I__2396\ : InMux
    port map (
            O => \N__10385\,
            I => \N__10374\
        );

    \I__2395\ : InMux
    port map (
            O => \N__10384\,
            I => \N__10371\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__10381\,
            I => \N__10368\
        );

    \I__2393\ : InMux
    port map (
            O => \N__10380\,
            I => \N__10365\
        );

    \I__2392\ : Span4Mux_v
    port map (
            O => \N__10377\,
            I => \N__10362\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__10374\,
            I => \N__10357\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__10371\,
            I => \N__10357\
        );

    \I__2389\ : Sp12to4
    port map (
            O => \N__10368\,
            I => \N__10354\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__10365\,
            I => \N__10351\
        );

    \I__2387\ : Sp12to4
    port map (
            O => \N__10362\,
            I => \N__10348\
        );

    \I__2386\ : Span4Mux_v
    port map (
            O => \N__10357\,
            I => \N__10345\
        );

    \I__2385\ : Span12Mux_h
    port map (
            O => \N__10354\,
            I => \N__10342\
        );

    \I__2384\ : Span12Mux_h
    port map (
            O => \N__10351\,
            I => \N__10339\
        );

    \I__2383\ : Span12Mux_h
    port map (
            O => \N__10348\,
            I => \N__10334\
        );

    \I__2382\ : Sp12to4
    port map (
            O => \N__10345\,
            I => \N__10334\
        );

    \I__2381\ : Span12Mux_v
    port map (
            O => \N__10342\,
            I => \N__10331\
        );

    \I__2380\ : Span12Mux_v
    port map (
            O => \N__10339\,
            I => \N__10328\
        );

    \I__2379\ : Span12Mux_h
    port map (
            O => \N__10334\,
            I => \N__10325\
        );

    \I__2378\ : Odrv12
    port map (
            O => \N__10331\,
            I => \RnW_c\
        );

    \I__2377\ : Odrv12
    port map (
            O => \N__10328\,
            I => \RnW_c\
        );

    \I__2376\ : Odrv12
    port map (
            O => \N__10325\,
            I => \RnW_c\
        );

    \I__2375\ : CascadeMux
    port map (
            O => \N__10318\,
            I => \N__10315\
        );

    \I__2374\ : InMux
    port map (
            O => \N__10315\,
            I => \N__10310\
        );

    \I__2373\ : InMux
    port map (
            O => \N__10314\,
            I => \N__10305\
        );

    \I__2372\ : InMux
    port map (
            O => \N__10313\,
            I => \N__10305\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__10310\,
            I => \N__10300\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__10305\,
            I => \N__10300\
        );

    \I__2369\ : Span4Mux_v
    port map (
            O => \N__10300\,
            I => \N__10295\
        );

    \I__2368\ : InMux
    port map (
            O => \N__10299\,
            I => \N__10292\
        );

    \I__2367\ : InMux
    port map (
            O => \N__10298\,
            I => \N__10289\
        );

    \I__2366\ : Span4Mux_v
    port map (
            O => \N__10295\,
            I => \N__10284\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__10292\,
            I => \N__10284\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__10289\,
            I => \N__10281\
        );

    \I__2363\ : Span4Mux_v
    port map (
            O => \N__10284\,
            I => \N__10278\
        );

    \I__2362\ : Span4Mux_v
    port map (
            O => \N__10281\,
            I => \N__10275\
        );

    \I__2361\ : Span4Mux_v
    port map (
            O => \N__10278\,
            I => \N__10271\
        );

    \I__2360\ : Sp12to4
    port map (
            O => \N__10275\,
            I => \N__10268\
        );

    \I__2359\ : InMux
    port map (
            O => \N__10274\,
            I => \N__10265\
        );

    \I__2358\ : Sp12to4
    port map (
            O => \N__10271\,
            I => \N__10262\
        );

    \I__2357\ : Span12Mux_h
    port map (
            O => \N__10268\,
            I => \N__10257\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__10265\,
            I => \N__10257\
        );

    \I__2355\ : Span12Mux_h
    port map (
            O => \N__10262\,
            I => \N__10252\
        );

    \I__2354\ : Span12Mux_v
    port map (
            O => \N__10257\,
            I => \N__10252\
        );

    \I__2353\ : Odrv12
    port map (
            O => \N__10252\,
            I => \CASLn_c\
        );

    \I__2352\ : InMux
    port map (
            O => \N__10249\,
            I => \N__10246\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__10246\,
            I => \N__10243\
        );

    \I__2350\ : Span12Mux_h
    port map (
            O => \N__10243\,
            I => \N__10240\
        );

    \I__2349\ : Odrv12
    port map (
            O => \N__10240\,
            I => \RAS1n_c\
        );

    \I__2348\ : InMux
    port map (
            O => \N__10237\,
            I => \N__10234\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__10234\,
            I => \N__10231\
        );

    \I__2346\ : Span4Mux_v
    port map (
            O => \N__10231\,
            I => \N__10227\
        );

    \I__2345\ : InMux
    port map (
            O => \N__10230\,
            I => \N__10224\
        );

    \I__2344\ : Sp12to4
    port map (
            O => \N__10227\,
            I => \N__10219\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__10224\,
            I => \N__10219\
        );

    \I__2342\ : Span12Mux_h
    port map (
            O => \N__10219\,
            I => \N__10216\
        );

    \I__2341\ : Odrv12
    port map (
            O => \N__10216\,
            I => \RAS0n_c\
        );

    \I__2340\ : InMux
    port map (
            O => \N__10213\,
            I => \N__10210\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__10210\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2338\ : InMux
    port map (
            O => \N__10207\,
            I => \N__10203\
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__10206\,
            I => \N__10194\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__10203\,
            I => \N__10190\
        );

    \I__2335\ : InMux
    port map (
            O => \N__10202\,
            I => \N__10187\
        );

    \I__2334\ : InMux
    port map (
            O => \N__10201\,
            I => \N__10184\
        );

    \I__2333\ : InMux
    port map (
            O => \N__10200\,
            I => \N__10178\
        );

    \I__2332\ : InMux
    port map (
            O => \N__10199\,
            I => \N__10178\
        );

    \I__2331\ : InMux
    port map (
            O => \N__10198\,
            I => \N__10175\
        );

    \I__2330\ : CascadeMux
    port map (
            O => \N__10197\,
            I => \N__10167\
        );

    \I__2329\ : InMux
    port map (
            O => \N__10194\,
            I => \N__10154\
        );

    \I__2328\ : InMux
    port map (
            O => \N__10193\,
            I => \N__10154\
        );

    \I__2327\ : Span4Mux_v
    port map (
            O => \N__10190\,
            I => \N__10145\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__10187\,
            I => \N__10145\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__10184\,
            I => \N__10145\
        );

    \I__2324\ : InMux
    port map (
            O => \N__10183\,
            I => \N__10142\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__10178\,
            I => \N__10136\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__10175\,
            I => \N__10136\
        );

    \I__2321\ : InMux
    port map (
            O => \N__10174\,
            I => \N__10131\
        );

    \I__2320\ : InMux
    port map (
            O => \N__10173\,
            I => \N__10131\
        );

    \I__2319\ : InMux
    port map (
            O => \N__10172\,
            I => \N__10128\
        );

    \I__2318\ : InMux
    port map (
            O => \N__10171\,
            I => \N__10121\
        );

    \I__2317\ : InMux
    port map (
            O => \N__10170\,
            I => \N__10121\
        );

    \I__2316\ : InMux
    port map (
            O => \N__10167\,
            I => \N__10121\
        );

    \I__2315\ : InMux
    port map (
            O => \N__10166\,
            I => \N__10118\
        );

    \I__2314\ : InMux
    port map (
            O => \N__10165\,
            I => \N__10113\
        );

    \I__2313\ : InMux
    port map (
            O => \N__10164\,
            I => \N__10113\
        );

    \I__2312\ : InMux
    port map (
            O => \N__10163\,
            I => \N__10104\
        );

    \I__2311\ : InMux
    port map (
            O => \N__10162\,
            I => \N__10104\
        );

    \I__2310\ : InMux
    port map (
            O => \N__10161\,
            I => \N__10104\
        );

    \I__2309\ : InMux
    port map (
            O => \N__10160\,
            I => \N__10104\
        );

    \I__2308\ : InMux
    port map (
            O => \N__10159\,
            I => \N__10098\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__10154\,
            I => \N__10095\
        );

    \I__2306\ : InMux
    port map (
            O => \N__10153\,
            I => \N__10092\
        );

    \I__2305\ : InMux
    port map (
            O => \N__10152\,
            I => \N__10089\
        );

    \I__2304\ : Span4Mux_v
    port map (
            O => \N__10145\,
            I => \N__10083\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__10142\,
            I => \N__10083\
        );

    \I__2302\ : InMux
    port map (
            O => \N__10141\,
            I => \N__10080\
        );

    \I__2301\ : Span4Mux_h
    port map (
            O => \N__10136\,
            I => \N__10071\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__10131\,
            I => \N__10071\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__10128\,
            I => \N__10071\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__10121\,
            I => \N__10071\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__10118\,
            I => \N__10064\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__10113\,
            I => \N__10064\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__10104\,
            I => \N__10064\
        );

    \I__2294\ : InMux
    port map (
            O => \N__10103\,
            I => \N__10057\
        );

    \I__2293\ : InMux
    port map (
            O => \N__10102\,
            I => \N__10057\
        );

    \I__2292\ : InMux
    port map (
            O => \N__10101\,
            I => \N__10057\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__10098\,
            I => \N__10052\
        );

    \I__2290\ : Span4Mux_h
    port map (
            O => \N__10095\,
            I => \N__10045\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__10092\,
            I => \N__10045\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__10089\,
            I => \N__10045\
        );

    \I__2287\ : InMux
    port map (
            O => \N__10088\,
            I => \N__10042\
        );

    \I__2286\ : Span4Mux_h
    port map (
            O => \N__10083\,
            I => \N__10037\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__10080\,
            I => \N__10037\
        );

    \I__2284\ : Span4Mux_v
    port map (
            O => \N__10071\,
            I => \N__10032\
        );

    \I__2283\ : Span4Mux_v
    port map (
            O => \N__10064\,
            I => \N__10032\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__10057\,
            I => \N__10029\
        );

    \I__2281\ : InMux
    port map (
            O => \N__10056\,
            I => \N__10024\
        );

    \I__2280\ : InMux
    port map (
            O => \N__10055\,
            I => \N__10024\
        );

    \I__2279\ : Span4Mux_v
    port map (
            O => \N__10052\,
            I => \N__10019\
        );

    \I__2278\ : Span4Mux_v
    port map (
            O => \N__10045\,
            I => \N__10019\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__10042\,
            I => \N__10014\
        );

    \I__2276\ : Sp12to4
    port map (
            O => \N__10037\,
            I => \N__10014\
        );

    \I__2275\ : Span4Mux_h
    port map (
            O => \N__10032\,
            I => \N__10009\
        );

    \I__2274\ : Span4Mux_v
    port map (
            O => \N__10029\,
            I => \N__10009\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__10024\,
            I => \N__10006\
        );

    \I__2272\ : Sp12to4
    port map (
            O => \N__10019\,
            I => \N__9999\
        );

    \I__2271\ : Span12Mux_v
    port map (
            O => \N__10014\,
            I => \N__9999\
        );

    \I__2270\ : Sp12to4
    port map (
            O => \N__10009\,
            I => \N__9999\
        );

    \I__2269\ : Span12Mux_h
    port map (
            O => \N__10006\,
            I => \N__9996\
        );

    \I__2268\ : Span12Mux_h
    port map (
            O => \N__9999\,
            I => \N__9993\
        );

    \I__2267\ : Odrv12
    port map (
            O => \N__9996\,
            I => \RESETn_c\
        );

    \I__2266\ : Odrv12
    port map (
            O => \N__9993\,
            I => \RESETn_c\
        );

    \I__2265\ : InMux
    port map (
            O => \N__9988\,
            I => \N__9985\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__9985\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\
        );

    \I__2263\ : InMux
    port map (
            O => \N__9982\,
            I => \N__9979\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__9979\,
            I => \N__9976\
        );

    \I__2261\ : Odrv12
    port map (
            O => \N__9976\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_2\
        );

    \I__2260\ : InMux
    port map (
            O => \N__9973\,
            I => \N__9970\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__9970\,
            I => \N__9931\
        );

    \I__2258\ : ClkMux
    port map (
            O => \N__9969\,
            I => \N__9832\
        );

    \I__2257\ : ClkMux
    port map (
            O => \N__9968\,
            I => \N__9832\
        );

    \I__2256\ : ClkMux
    port map (
            O => \N__9967\,
            I => \N__9832\
        );

    \I__2255\ : ClkMux
    port map (
            O => \N__9966\,
            I => \N__9832\
        );

    \I__2254\ : ClkMux
    port map (
            O => \N__9965\,
            I => \N__9832\
        );

    \I__2253\ : ClkMux
    port map (
            O => \N__9964\,
            I => \N__9832\
        );

    \I__2252\ : ClkMux
    port map (
            O => \N__9963\,
            I => \N__9832\
        );

    \I__2251\ : ClkMux
    port map (
            O => \N__9962\,
            I => \N__9832\
        );

    \I__2250\ : ClkMux
    port map (
            O => \N__9961\,
            I => \N__9832\
        );

    \I__2249\ : ClkMux
    port map (
            O => \N__9960\,
            I => \N__9832\
        );

    \I__2248\ : ClkMux
    port map (
            O => \N__9959\,
            I => \N__9832\
        );

    \I__2247\ : ClkMux
    port map (
            O => \N__9958\,
            I => \N__9832\
        );

    \I__2246\ : ClkMux
    port map (
            O => \N__9957\,
            I => \N__9832\
        );

    \I__2245\ : ClkMux
    port map (
            O => \N__9956\,
            I => \N__9832\
        );

    \I__2244\ : ClkMux
    port map (
            O => \N__9955\,
            I => \N__9832\
        );

    \I__2243\ : ClkMux
    port map (
            O => \N__9954\,
            I => \N__9832\
        );

    \I__2242\ : ClkMux
    port map (
            O => \N__9953\,
            I => \N__9832\
        );

    \I__2241\ : ClkMux
    port map (
            O => \N__9952\,
            I => \N__9832\
        );

    \I__2240\ : ClkMux
    port map (
            O => \N__9951\,
            I => \N__9832\
        );

    \I__2239\ : ClkMux
    port map (
            O => \N__9950\,
            I => \N__9832\
        );

    \I__2238\ : ClkMux
    port map (
            O => \N__9949\,
            I => \N__9832\
        );

    \I__2237\ : ClkMux
    port map (
            O => \N__9948\,
            I => \N__9832\
        );

    \I__2236\ : ClkMux
    port map (
            O => \N__9947\,
            I => \N__9832\
        );

    \I__2235\ : ClkMux
    port map (
            O => \N__9946\,
            I => \N__9832\
        );

    \I__2234\ : ClkMux
    port map (
            O => \N__9945\,
            I => \N__9832\
        );

    \I__2233\ : ClkMux
    port map (
            O => \N__9944\,
            I => \N__9832\
        );

    \I__2232\ : ClkMux
    port map (
            O => \N__9943\,
            I => \N__9832\
        );

    \I__2231\ : ClkMux
    port map (
            O => \N__9942\,
            I => \N__9832\
        );

    \I__2230\ : ClkMux
    port map (
            O => \N__9941\,
            I => \N__9832\
        );

    \I__2229\ : ClkMux
    port map (
            O => \N__9940\,
            I => \N__9832\
        );

    \I__2228\ : ClkMux
    port map (
            O => \N__9939\,
            I => \N__9832\
        );

    \I__2227\ : ClkMux
    port map (
            O => \N__9938\,
            I => \N__9832\
        );

    \I__2226\ : ClkMux
    port map (
            O => \N__9937\,
            I => \N__9832\
        );

    \I__2225\ : ClkMux
    port map (
            O => \N__9936\,
            I => \N__9832\
        );

    \I__2224\ : ClkMux
    port map (
            O => \N__9935\,
            I => \N__9832\
        );

    \I__2223\ : ClkMux
    port map (
            O => \N__9934\,
            I => \N__9832\
        );

    \I__2222\ : Glb2LocalMux
    port map (
            O => \N__9931\,
            I => \N__9832\
        );

    \I__2221\ : ClkMux
    port map (
            O => \N__9930\,
            I => \N__9832\
        );

    \I__2220\ : ClkMux
    port map (
            O => \N__9929\,
            I => \N__9832\
        );

    \I__2219\ : ClkMux
    port map (
            O => \N__9928\,
            I => \N__9832\
        );

    \I__2218\ : ClkMux
    port map (
            O => \N__9927\,
            I => \N__9832\
        );

    \I__2217\ : ClkMux
    port map (
            O => \N__9926\,
            I => \N__9832\
        );

    \I__2216\ : ClkMux
    port map (
            O => \N__9925\,
            I => \N__9832\
        );

    \I__2215\ : ClkMux
    port map (
            O => \N__9924\,
            I => \N__9832\
        );

    \I__2214\ : ClkMux
    port map (
            O => \N__9923\,
            I => \N__9832\
        );

    \I__2213\ : GlobalMux
    port map (
            O => \N__9832\,
            I => \CLK80_PLL\
        );

    \I__2212\ : InMux
    port map (
            O => \N__9829\,
            I => \N__9823\
        );

    \I__2211\ : InMux
    port map (
            O => \N__9828\,
            I => \N__9823\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__9823\,
            I => \N__9818\
        );

    \I__2209\ : InMux
    port map (
            O => \N__9822\,
            I => \N__9815\
        );

    \I__2208\ : InMux
    port map (
            O => \N__9821\,
            I => \N__9812\
        );

    \I__2207\ : Span4Mux_v
    port map (
            O => \N__9818\,
            I => \N__9809\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__9815\,
            I => \N__9806\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__9812\,
            I => \N__9803\
        );

    \I__2204\ : Sp12to4
    port map (
            O => \N__9809\,
            I => \N__9800\
        );

    \I__2203\ : Sp12to4
    port map (
            O => \N__9806\,
            I => \N__9797\
        );

    \I__2202\ : Span12Mux_h
    port map (
            O => \N__9803\,
            I => \N__9794\
        );

    \I__2201\ : Span12Mux_h
    port map (
            O => \N__9800\,
            I => \N__9791\
        );

    \I__2200\ : Span12Mux_v
    port map (
            O => \N__9797\,
            I => \N__9788\
        );

    \I__2199\ : Span12Mux_v
    port map (
            O => \N__9794\,
            I => \N__9785\
        );

    \I__2198\ : Span12Mux_v
    port map (
            O => \N__9791\,
            I => \N__9780\
        );

    \I__2197\ : Span12Mux_h
    port map (
            O => \N__9788\,
            I => \N__9780\
        );

    \I__2196\ : Odrv12
    port map (
            O => \N__9785\,
            I => \DRA_c_1\
        );

    \I__2195\ : Odrv12
    port map (
            O => \N__9780\,
            I => \DRA_c_1\
        );

    \I__2194\ : InMux
    port map (
            O => \N__9775\,
            I => \N__9771\
        );

    \I__2193\ : InMux
    port map (
            O => \N__9774\,
            I => \N__9768\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__9771\,
            I => \N__9763\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__9768\,
            I => \N__9763\
        );

    \I__2190\ : Span12Mux_h
    port map (
            O => \N__9763\,
            I => \N__9760\
        );

    \I__2189\ : Span12Mux_v
    port map (
            O => \N__9760\,
            I => \N__9757\
        );

    \I__2188\ : Odrv12
    port map (
            O => \N__9757\,
            I => \DRA_c_0\
        );

    \I__2187\ : InMux
    port map (
            O => \N__9754\,
            I => \N__9751\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__9751\,
            I => \N__9748\
        );

    \I__2185\ : Span4Mux_v
    port map (
            O => \N__9748\,
            I => \N__9745\
        );

    \I__2184\ : Span4Mux_h
    port map (
            O => \N__9745\,
            I => \N__9742\
        );

    \I__2183\ : Odrv4
    port map (
            O => \N__9742\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__2182\ : CascadeMux
    port map (
            O => \N__9739\,
            I => \N_334_cascade_\
        );

    \I__2181\ : IoInMux
    port map (
            O => \N__9736\,
            I => \N__9733\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__9733\,
            I => \N__9730\
        );

    \I__2179\ : Span4Mux_s3_h
    port map (
            O => \N__9730\,
            I => \N__9727\
        );

    \I__2178\ : Sp12to4
    port map (
            O => \N__9727\,
            I => \N__9724\
        );

    \I__2177\ : Span12Mux_s8_v
    port map (
            O => \N__9724\,
            I => \N__9721\
        );

    \I__2176\ : Span12Mux_h
    port map (
            O => \N__9721\,
            I => \N__9718\
        );

    \I__2175\ : Odrv12
    port map (
            O => \N__9718\,
            I => \N_177_i\
        );

    \I__2174\ : InMux
    port map (
            O => \N__9715\,
            I => \N__9711\
        );

    \I__2173\ : InMux
    port map (
            O => \N__9714\,
            I => \N__9708\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__9711\,
            I => \N__9704\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__9708\,
            I => \N__9701\
        );

    \I__2170\ : InMux
    port map (
            O => \N__9707\,
            I => \N__9698\
        );

    \I__2169\ : Span4Mux_v
    port map (
            O => \N__9704\,
            I => \N__9690\
        );

    \I__2168\ : Span4Mux_h
    port map (
            O => \N__9701\,
            I => \N__9690\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__9698\,
            I => \N__9690\
        );

    \I__2166\ : InMux
    port map (
            O => \N__9697\,
            I => \N__9687\
        );

    \I__2165\ : Span4Mux_v
    port map (
            O => \N__9690\,
            I => \N__9684\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__9687\,
            I => \N__9681\
        );

    \I__2163\ : Span4Mux_v
    port map (
            O => \N__9684\,
            I => \N__9678\
        );

    \I__2162\ : Span12Mux_v
    port map (
            O => \N__9681\,
            I => \N__9673\
        );

    \I__2161\ : Sp12to4
    port map (
            O => \N__9678\,
            I => \N__9673\
        );

    \I__2160\ : Span12Mux_h
    port map (
            O => \N__9673\,
            I => \N__9670\
        );

    \I__2159\ : Odrv12
    port map (
            O => \N__9670\,
            I => \DRA_c_2\
        );

    \I__2158\ : InMux
    port map (
            O => \N__9667\,
            I => \N__9664\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__9664\,
            I => \N__9661\
        );

    \I__2156\ : Odrv4
    port map (
            O => \N__9661\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__2155\ : InMux
    port map (
            O => \N__9658\,
            I => \N__9655\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__9655\,
            I => \N__9652\
        );

    \I__2153\ : Odrv4
    port map (
            O => \N__9652\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__2152\ : InMux
    port map (
            O => \N__9649\,
            I => \N__9646\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__9646\,
            I => \N__9642\
        );

    \I__2150\ : InMux
    port map (
            O => \N__9645\,
            I => \N__9639\
        );

    \I__2149\ : Span4Mux_v
    port map (
            O => \N__9642\,
            I => \N__9634\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__9639\,
            I => \N__9631\
        );

    \I__2147\ : InMux
    port map (
            O => \N__9638\,
            I => \N__9628\
        );

    \I__2146\ : InMux
    port map (
            O => \N__9637\,
            I => \N__9625\
        );

    \I__2145\ : Span4Mux_v
    port map (
            O => \N__9634\,
            I => \N__9622\
        );

    \I__2144\ : Sp12to4
    port map (
            O => \N__9631\,
            I => \N__9615\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__9628\,
            I => \N__9615\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__9625\,
            I => \N__9615\
        );

    \I__2141\ : Sp12to4
    port map (
            O => \N__9622\,
            I => \N__9610\
        );

    \I__2140\ : Span12Mux_v
    port map (
            O => \N__9615\,
            I => \N__9610\
        );

    \I__2139\ : Span12Mux_h
    port map (
            O => \N__9610\,
            I => \N__9607\
        );

    \I__2138\ : Odrv12
    port map (
            O => \N__9607\,
            I => \DRA_c_5\
        );

    \I__2137\ : InMux
    port map (
            O => \N__9604\,
            I => \N__9601\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9601\,
            I => \N__9598\
        );

    \I__2135\ : Span12Mux_v
    port map (
            O => \N__9598\,
            I => \N__9595\
        );

    \I__2134\ : Odrv12
    port map (
            O => \N__9595\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__2133\ : IoInMux
    port map (
            O => \N__9592\,
            I => \N__9589\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__9589\,
            I => \N__9586\
        );

    \I__2131\ : Odrv12
    port map (
            O => \N__9586\,
            I => \RESETn_c_i\
        );

    \I__2130\ : InMux
    port map (
            O => \N__9583\,
            I => \N__9580\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__9580\,
            I => \N__9576\
        );

    \I__2128\ : InMux
    port map (
            O => \N__9579\,
            I => \N__9573\
        );

    \I__2127\ : Span4Mux_h
    port map (
            O => \N__9576\,
            I => \N__9567\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__9573\,
            I => \N__9567\
        );

    \I__2125\ : CascadeMux
    port map (
            O => \N__9572\,
            I => \N__9562\
        );

    \I__2124\ : Span4Mux_h
    port map (
            O => \N__9567\,
            I => \N__9559\
        );

    \I__2123\ : InMux
    port map (
            O => \N__9566\,
            I => \N__9556\
        );

    \I__2122\ : InMux
    port map (
            O => \N__9565\,
            I => \N__9553\
        );

    \I__2121\ : InMux
    port map (
            O => \N__9562\,
            I => \N__9550\
        );

    \I__2120\ : Odrv4
    port map (
            O => \N__9559\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__9556\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__9553\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__9550\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2116\ : IoInMux
    port map (
            O => \N__9541\,
            I => \N__9538\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__9538\,
            I => \N__9535\
        );

    \I__2114\ : Span4Mux_s2_v
    port map (
            O => \N__9535\,
            I => \N__9532\
        );

    \I__2113\ : Span4Mux_v
    port map (
            O => \N__9532\,
            I => \N__9529\
        );

    \I__2112\ : Span4Mux_v
    port map (
            O => \N__9529\,
            I => \N__9526\
        );

    \I__2111\ : Span4Mux_h
    port map (
            O => \N__9526\,
            I => \N__9523\
        );

    \I__2110\ : Odrv4
    port map (
            O => \N__9523\,
            I => \CRCSn_c\
        );

    \I__2109\ : InMux
    port map (
            O => \N__9520\,
            I => \N__9517\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__9517\,
            I => \N__9514\
        );

    \I__2107\ : Odrv12
    port map (
            O => \N__9514\,
            I => \U712_CHIP_RAM.CMA_5_i_0_9\
        );

    \I__2106\ : InMux
    port map (
            O => \N__9511\,
            I => \N__9508\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__9508\,
            I => \N__9505\
        );

    \I__2104\ : Span4Mux_v
    port map (
            O => \N__9505\,
            I => \N__9502\
        );

    \I__2103\ : Span4Mux_v
    port map (
            O => \N__9502\,
            I => \N__9499\
        );

    \I__2102\ : Sp12to4
    port map (
            O => \N__9499\,
            I => \N__9496\
        );

    \I__2101\ : Span12Mux_h
    port map (
            O => \N__9496\,
            I => \N__9493\
        );

    \I__2100\ : Odrv12
    port map (
            O => \N__9493\,
            I => \A_c_19\
        );

    \I__2099\ : InMux
    port map (
            O => \N__9490\,
            I => \N__9487\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__9487\,
            I => \N__9484\
        );

    \I__2097\ : Odrv4
    port map (
            O => \N__9484\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2096\ : IoInMux
    port map (
            O => \N__9481\,
            I => \N__9478\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__9478\,
            I => \N__9475\
        );

    \I__2094\ : Span4Mux_s3_h
    port map (
            O => \N__9475\,
            I => \N__9472\
        );

    \I__2093\ : Sp12to4
    port map (
            O => \N__9472\,
            I => \N__9469\
        );

    \I__2092\ : Span12Mux_s10_v
    port map (
            O => \N__9469\,
            I => \N__9466\
        );

    \I__2091\ : Span12Mux_h
    port map (
            O => \N__9466\,
            I => \N__9463\
        );

    \I__2090\ : Odrv12
    port map (
            O => \N__9463\,
            I => \CMA_c_9\
        );

    \I__2089\ : CEMux
    port map (
            O => \N__9460\,
            I => \N__9455\
        );

    \I__2088\ : CEMux
    port map (
            O => \N__9459\,
            I => \N__9452\
        );

    \I__2087\ : CEMux
    port map (
            O => \N__9458\,
            I => \N__9448\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__9455\,
            I => \N__9445\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__9452\,
            I => \N__9441\
        );

    \I__2084\ : CEMux
    port map (
            O => \N__9451\,
            I => \N__9438\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__9448\,
            I => \N__9435\
        );

    \I__2082\ : Span4Mux_v
    port map (
            O => \N__9445\,
            I => \N__9432\
        );

    \I__2081\ : CEMux
    port map (
            O => \N__9444\,
            I => \N__9429\
        );

    \I__2080\ : Span4Mux_h
    port map (
            O => \N__9441\,
            I => \N__9424\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__9438\,
            I => \N__9424\
        );

    \I__2078\ : Span4Mux_h
    port map (
            O => \N__9435\,
            I => \N__9421\
        );

    \I__2077\ : Span4Mux_h
    port map (
            O => \N__9432\,
            I => \N__9418\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__9429\,
            I => \N__9415\
        );

    \I__2075\ : Sp12to4
    port map (
            O => \N__9424\,
            I => \N__9412\
        );

    \I__2074\ : Odrv4
    port map (
            O => \N__9421\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__2073\ : Odrv4
    port map (
            O => \N__9418\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__2072\ : Odrv4
    port map (
            O => \N__9415\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__2071\ : Odrv12
    port map (
            O => \N__9412\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__2070\ : CascadeMux
    port map (
            O => \N__9403\,
            I => \N__9400\
        );

    \I__2069\ : InMux
    port map (
            O => \N__9400\,
            I => \N__9397\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__9397\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__2067\ : InMux
    port map (
            O => \N__9394\,
            I => \N__9391\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__9391\,
            I => \N__9388\
        );

    \I__2065\ : Span4Mux_h
    port map (
            O => \N__9388\,
            I => \N__9385\
        );

    \I__2064\ : Odrv4
    port map (
            O => \N__9385\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__2063\ : InMux
    port map (
            O => \N__9382\,
            I => \N__9379\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__9379\,
            I => \N__9376\
        );

    \I__2061\ : Span4Mux_v
    port map (
            O => \N__9376\,
            I => \N__9373\
        );

    \I__2060\ : Odrv4
    port map (
            O => \N__9373\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__2059\ : InMux
    port map (
            O => \N__9370\,
            I => \N__9367\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__9367\,
            I => \N__9364\
        );

    \I__2057\ : Span4Mux_h
    port map (
            O => \N__9364\,
            I => \N__9361\
        );

    \I__2056\ : Odrv4
    port map (
            O => \N__9361\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__2055\ : InMux
    port map (
            O => \N__9358\,
            I => \N__9355\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__9355\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2053\ : InMux
    port map (
            O => \N__9352\,
            I => \N__9349\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__9349\,
            I => \N__9346\
        );

    \I__2051\ : Odrv4
    port map (
            O => \N__9346\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2050\ : InMux
    port map (
            O => \N__9343\,
            I => \N__9340\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__9340\,
            I => \N__9337\
        );

    \I__2048\ : Odrv4
    port map (
            O => \N__9337\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__2047\ : InMux
    port map (
            O => \N__9334\,
            I => \N__9326\
        );

    \I__2046\ : InMux
    port map (
            O => \N__9333\,
            I => \N__9326\
        );

    \I__2045\ : InMux
    port map (
            O => \N__9332\,
            I => \N__9323\
        );

    \I__2044\ : InMux
    port map (
            O => \N__9331\,
            I => \N__9320\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__9326\,
            I => \N__9317\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__9323\,
            I => \N__9312\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__9320\,
            I => \N__9312\
        );

    \I__2040\ : Span4Mux_v
    port map (
            O => \N__9317\,
            I => \N__9309\
        );

    \I__2039\ : Span4Mux_h
    port map (
            O => \N__9312\,
            I => \N__9306\
        );

    \I__2038\ : Span4Mux_h
    port map (
            O => \N__9309\,
            I => \N__9303\
        );

    \I__2037\ : Span4Mux_h
    port map (
            O => \N__9306\,
            I => \N__9300\
        );

    \I__2036\ : Sp12to4
    port map (
            O => \N__9303\,
            I => \N__9295\
        );

    \I__2035\ : Sp12to4
    port map (
            O => \N__9300\,
            I => \N__9295\
        );

    \I__2034\ : Odrv12
    port map (
            O => \N__9295\,
            I => \DRA_c_8\
        );

    \I__2033\ : InMux
    port map (
            O => \N__9292\,
            I => \N__9289\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__9289\,
            I => \N__9286\
        );

    \I__2031\ : Span4Mux_h
    port map (
            O => \N__9286\,
            I => \N__9283\
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__9283\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__2029\ : InMux
    port map (
            O => \N__9280\,
            I => \N__9277\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__9277\,
            I => \N__9274\
        );

    \I__2027\ : Odrv12
    port map (
            O => \N__9274\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2026\ : InMux
    port map (
            O => \N__9271\,
            I => \N__9265\
        );

    \I__2025\ : InMux
    port map (
            O => \N__9270\,
            I => \N__9265\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__9265\,
            I => \N__9262\
        );

    \I__2023\ : Span4Mux_v
    port map (
            O => \N__9262\,
            I => \N__9259\
        );

    \I__2022\ : Odrv4
    port map (
            O => \N__9259\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__2021\ : InMux
    port map (
            O => \N__9256\,
            I => \N__9252\
        );

    \I__2020\ : CascadeMux
    port map (
            O => \N__9255\,
            I => \N__9249\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__9252\,
            I => \N__9246\
        );

    \I__2018\ : InMux
    port map (
            O => \N__9249\,
            I => \N__9243\
        );

    \I__2017\ : Odrv12
    port map (
            O => \N__9246\,
            I => \U712_CHIP_RAM.m50_i_a2_0_0\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__9243\,
            I => \U712_CHIP_RAM.m50_i_a2_0_0\
        );

    \I__2015\ : IoInMux
    port map (
            O => \N__9238\,
            I => \N__9235\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__9235\,
            I => \N__9232\
        );

    \I__2013\ : Span12Mux_s4_h
    port map (
            O => \N__9232\,
            I => \N__9229\
        );

    \I__2012\ : Span12Mux_v
    port map (
            O => \N__9229\,
            I => \N__9226\
        );

    \I__2011\ : Span12Mux_h
    port map (
            O => \N__9226\,
            I => \N__9223\
        );

    \I__2010\ : Odrv12
    port map (
            O => \N__9223\,
            I => \N_200_i\
        );

    \I__2009\ : InMux
    port map (
            O => \N__9220\,
            I => \N__9217\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__9217\,
            I => \N__9214\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__9214\,
            I => \U712_CHIP_RAM.N_337\
        );

    \I__2006\ : CascadeMux
    port map (
            O => \N__9211\,
            I => \N__9205\
        );

    \I__2005\ : InMux
    port map (
            O => \N__9210\,
            I => \N__9202\
        );

    \I__2004\ : InMux
    port map (
            O => \N__9209\,
            I => \N__9199\
        );

    \I__2003\ : InMux
    port map (
            O => \N__9208\,
            I => \N__9196\
        );

    \I__2002\ : InMux
    port map (
            O => \N__9205\,
            I => \N__9193\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__9202\,
            I => \N__9190\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__9199\,
            I => \N__9185\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__9196\,
            I => \N__9185\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__9193\,
            I => \N__9182\
        );

    \I__1997\ : Span4Mux_v
    port map (
            O => \N__9190\,
            I => \N__9179\
        );

    \I__1996\ : Span4Mux_v
    port map (
            O => \N__9185\,
            I => \N__9176\
        );

    \I__1995\ : Span4Mux_v
    port map (
            O => \N__9182\,
            I => \N__9173\
        );

    \I__1994\ : Span4Mux_h
    port map (
            O => \N__9179\,
            I => \N__9170\
        );

    \I__1993\ : Sp12to4
    port map (
            O => \N__9176\,
            I => \N__9167\
        );

    \I__1992\ : Sp12to4
    port map (
            O => \N__9173\,
            I => \N__9164\
        );

    \I__1991\ : Sp12to4
    port map (
            O => \N__9170\,
            I => \N__9157\
        );

    \I__1990\ : Span12Mux_h
    port map (
            O => \N__9167\,
            I => \N__9157\
        );

    \I__1989\ : Span12Mux_h
    port map (
            O => \N__9164\,
            I => \N__9157\
        );

    \I__1988\ : Span12Mux_v
    port map (
            O => \N__9157\,
            I => \N__9154\
        );

    \I__1987\ : Odrv12
    port map (
            O => \N__9154\,
            I => \CLK40_PLL_i\
        );

    \I__1986\ : IoInMux
    port map (
            O => \N__9151\,
            I => \N__9148\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__9148\,
            I => \N__9143\
        );

    \I__1984\ : IoInMux
    port map (
            O => \N__9147\,
            I => \N__9140\
        );

    \I__1983\ : IoInMux
    port map (
            O => \N__9146\,
            I => \N__9137\
        );

    \I__1982\ : IoSpan4Mux
    port map (
            O => \N__9143\,
            I => \N__9132\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__9140\,
            I => \N__9132\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__9137\,
            I => \N__9129\
        );

    \I__1979\ : IoSpan4Mux
    port map (
            O => \N__9132\,
            I => \N__9126\
        );

    \I__1978\ : Span4Mux_s2_h
    port map (
            O => \N__9129\,
            I => \N__9123\
        );

    \I__1977\ : Span4Mux_s0_v
    port map (
            O => \N__9126\,
            I => \N__9120\
        );

    \I__1976\ : Span4Mux_v
    port map (
            O => \N__9123\,
            I => \N__9117\
        );

    \I__1975\ : Sp12to4
    port map (
            O => \N__9120\,
            I => \N__9114\
        );

    \I__1974\ : Sp12to4
    port map (
            O => \N__9117\,
            I => \N__9111\
        );

    \I__1973\ : Span12Mux_v
    port map (
            O => \N__9114\,
            I => \N__9106\
        );

    \I__1972\ : Span12Mux_h
    port map (
            O => \N__9111\,
            I => \N__9106\
        );

    \I__1971\ : Odrv12
    port map (
            O => \N__9106\,
            I => \CLK40_PLL_i_i\
        );

    \I__1970\ : InMux
    port map (
            O => \N__9103\,
            I => \N__9100\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__9100\,
            I => \N__9097\
        );

    \I__1968\ : Odrv4
    port map (
            O => \N__9097\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\
        );

    \I__1967\ : IoInMux
    port map (
            O => \N__9094\,
            I => \N__9091\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__9091\,
            I => \N__9088\
        );

    \I__1965\ : IoSpan4Mux
    port map (
            O => \N__9088\,
            I => \N__9085\
        );

    \I__1964\ : Span4Mux_s3_h
    port map (
            O => \N__9085\,
            I => \N__9082\
        );

    \I__1963\ : Span4Mux_v
    port map (
            O => \N__9082\,
            I => \N__9079\
        );

    \I__1962\ : Span4Mux_h
    port map (
            O => \N__9079\,
            I => \N__9076\
        );

    \I__1961\ : Sp12to4
    port map (
            O => \N__9076\,
            I => \N__9073\
        );

    \I__1960\ : Odrv12
    port map (
            O => \N__9073\,
            I => \CMA_c_8\
        );

    \I__1959\ : IoInMux
    port map (
            O => \N__9070\,
            I => \N__9067\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__9067\,
            I => \N__9064\
        );

    \I__1957\ : Span4Mux_s0_v
    port map (
            O => \N__9064\,
            I => \N__9061\
        );

    \I__1956\ : Sp12to4
    port map (
            O => \N__9061\,
            I => \N__9058\
        );

    \I__1955\ : Span12Mux_h
    port map (
            O => \N__9058\,
            I => \N__9055\
        );

    \I__1954\ : Odrv12
    port map (
            O => \N__9055\,
            I => \CMA_c_0\
        );

    \I__1953\ : InMux
    port map (
            O => \N__9052\,
            I => \N__9049\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__9049\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__1951\ : IoInMux
    port map (
            O => \N__9046\,
            I => \N__9043\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__9043\,
            I => \N__9040\
        );

    \I__1949\ : IoSpan4Mux
    port map (
            O => \N__9040\,
            I => \N__9037\
        );

    \I__1948\ : Span4Mux_s2_h
    port map (
            O => \N__9037\,
            I => \N__9034\
        );

    \I__1947\ : Sp12to4
    port map (
            O => \N__9034\,
            I => \N__9031\
        );

    \I__1946\ : Span12Mux_h
    port map (
            O => \N__9031\,
            I => \N__9028\
        );

    \I__1945\ : Odrv12
    port map (
            O => \N__9028\,
            I => \CMA_c_7\
        );

    \I__1944\ : IoInMux
    port map (
            O => \N__9025\,
            I => \N__9022\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__9022\,
            I => \N__9018\
        );

    \I__1942\ : InMux
    port map (
            O => \N__9021\,
            I => \N__9015\
        );

    \I__1941\ : Span12Mux_s4_v
    port map (
            O => \N__9018\,
            I => \N__9012\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__9015\,
            I => \N__9009\
        );

    \I__1939\ : Span12Mux_v
    port map (
            O => \N__9012\,
            I => \N__9004\
        );

    \I__1938\ : Span12Mux_v
    port map (
            O => \N__9009\,
            I => \N__9004\
        );

    \I__1937\ : Span12Mux_h
    port map (
            O => \N__9004\,
            I => \N__9001\
        );

    \I__1936\ : Odrv12
    port map (
            O => \N__9001\,
            I => \A_c_9\
        );

    \I__1935\ : InMux
    port map (
            O => \N__8998\,
            I => \N__8995\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__8995\,
            I => \N__8992\
        );

    \I__1933\ : Odrv12
    port map (
            O => \N__8992\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\
        );

    \I__1932\ : CascadeMux
    port map (
            O => \N__8989\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\
        );

    \I__1931\ : InMux
    port map (
            O => \N__8986\,
            I => \N__8983\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__8983\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__1929\ : InMux
    port map (
            O => \N__8980\,
            I => \N__8977\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__8977\,
            I => \N__8974\
        );

    \I__1927\ : Odrv4
    port map (
            O => \N__8974\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\
        );

    \I__1926\ : CascadeMux
    port map (
            O => \N__8971\,
            I => \N__8967\
        );

    \I__1925\ : InMux
    port map (
            O => \N__8970\,
            I => \N__8953\
        );

    \I__1924\ : InMux
    port map (
            O => \N__8967\,
            I => \N__8953\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__8966\,
            I => \N__8946\
        );

    \I__1922\ : CascadeMux
    port map (
            O => \N__8965\,
            I => \N__8943\
        );

    \I__1921\ : CascadeMux
    port map (
            O => \N__8964\,
            I => \N__8939\
        );

    \I__1920\ : InMux
    port map (
            O => \N__8963\,
            I => \N__8933\
        );

    \I__1919\ : InMux
    port map (
            O => \N__8962\,
            I => \N__8933\
        );

    \I__1918\ : InMux
    port map (
            O => \N__8961\,
            I => \N__8926\
        );

    \I__1917\ : InMux
    port map (
            O => \N__8960\,
            I => \N__8926\
        );

    \I__1916\ : InMux
    port map (
            O => \N__8959\,
            I => \N__8926\
        );

    \I__1915\ : InMux
    port map (
            O => \N__8958\,
            I => \N__8923\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__8953\,
            I => \N__8920\
        );

    \I__1913\ : InMux
    port map (
            O => \N__8952\,
            I => \N__8913\
        );

    \I__1912\ : InMux
    port map (
            O => \N__8951\,
            I => \N__8913\
        );

    \I__1911\ : InMux
    port map (
            O => \N__8950\,
            I => \N__8913\
        );

    \I__1910\ : InMux
    port map (
            O => \N__8949\,
            I => \N__8910\
        );

    \I__1909\ : InMux
    port map (
            O => \N__8946\,
            I => \N__8907\
        );

    \I__1908\ : InMux
    port map (
            O => \N__8943\,
            I => \N__8902\
        );

    \I__1907\ : InMux
    port map (
            O => \N__8942\,
            I => \N__8902\
        );

    \I__1906\ : InMux
    port map (
            O => \N__8939\,
            I => \N__8897\
        );

    \I__1905\ : InMux
    port map (
            O => \N__8938\,
            I => \N__8897\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__8933\,
            I => \N__8892\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__8926\,
            I => \N__8892\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__8923\,
            I => \N__8885\
        );

    \I__1901\ : Span4Mux_v
    port map (
            O => \N__8920\,
            I => \N__8880\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__8913\,
            I => \N__8880\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__8910\,
            I => \N__8875\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__8907\,
            I => \N__8875\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__8902\,
            I => \N__8870\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__8897\,
            I => \N__8870\
        );

    \I__1895\ : Span4Mux_v
    port map (
            O => \N__8892\,
            I => \N__8867\
        );

    \I__1894\ : InMux
    port map (
            O => \N__8891\,
            I => \N__8860\
        );

    \I__1893\ : InMux
    port map (
            O => \N__8890\,
            I => \N__8860\
        );

    \I__1892\ : InMux
    port map (
            O => \N__8889\,
            I => \N__8860\
        );

    \I__1891\ : InMux
    port map (
            O => \N__8888\,
            I => \N__8853\
        );

    \I__1890\ : Span4Mux_h
    port map (
            O => \N__8885\,
            I => \N__8848\
        );

    \I__1889\ : Span4Mux_h
    port map (
            O => \N__8880\,
            I => \N__8848\
        );

    \I__1888\ : Span4Mux_v
    port map (
            O => \N__8875\,
            I => \N__8839\
        );

    \I__1887\ : Span4Mux_h
    port map (
            O => \N__8870\,
            I => \N__8839\
        );

    \I__1886\ : Span4Mux_h
    port map (
            O => \N__8867\,
            I => \N__8839\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__8860\,
            I => \N__8839\
        );

    \I__1884\ : InMux
    port map (
            O => \N__8859\,
            I => \N__8830\
        );

    \I__1883\ : InMux
    port map (
            O => \N__8858\,
            I => \N__8830\
        );

    \I__1882\ : InMux
    port map (
            O => \N__8857\,
            I => \N__8830\
        );

    \I__1881\ : InMux
    port map (
            O => \N__8856\,
            I => \N__8830\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__8853\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1879\ : Odrv4
    port map (
            O => \N__8848\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1878\ : Odrv4
    port map (
            O => \N__8839\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__8830\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1876\ : InMux
    port map (
            O => \N__8821\,
            I => \N__8812\
        );

    \I__1875\ : InMux
    port map (
            O => \N__8820\,
            I => \N__8809\
        );

    \I__1874\ : InMux
    port map (
            O => \N__8819\,
            I => \N__8802\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8818\,
            I => \N__8802\
        );

    \I__1872\ : InMux
    port map (
            O => \N__8817\,
            I => \N__8802\
        );

    \I__1871\ : InMux
    port map (
            O => \N__8816\,
            I => \N__8797\
        );

    \I__1870\ : InMux
    port map (
            O => \N__8815\,
            I => \N__8797\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__8812\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__8809\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__8802\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__8797\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0\
        );

    \I__1865\ : CascadeMux
    port map (
            O => \N__8788\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_\
        );

    \I__1864\ : CascadeMux
    port map (
            O => \N__8785\,
            I => \N__8778\
        );

    \I__1863\ : CascadeMux
    port map (
            O => \N__8784\,
            I => \N__8775\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__8783\,
            I => \N__8772\
        );

    \I__1861\ : CascadeMux
    port map (
            O => \N__8782\,
            I => \N__8767\
        );

    \I__1860\ : CascadeMux
    port map (
            O => \N__8781\,
            I => \N__8764\
        );

    \I__1859\ : InMux
    port map (
            O => \N__8778\,
            I => \N__8761\
        );

    \I__1858\ : InMux
    port map (
            O => \N__8775\,
            I => \N__8756\
        );

    \I__1857\ : InMux
    port map (
            O => \N__8772\,
            I => \N__8756\
        );

    \I__1856\ : CascadeMux
    port map (
            O => \N__8771\,
            I => \N__8753\
        );

    \I__1855\ : InMux
    port map (
            O => \N__8770\,
            I => \N__8748\
        );

    \I__1854\ : InMux
    port map (
            O => \N__8767\,
            I => \N__8743\
        );

    \I__1853\ : InMux
    port map (
            O => \N__8764\,
            I => \N__8743\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__8761\,
            I => \N__8738\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__8756\,
            I => \N__8738\
        );

    \I__1850\ : InMux
    port map (
            O => \N__8753\,
            I => \N__8734\
        );

    \I__1849\ : InMux
    port map (
            O => \N__8752\,
            I => \N__8731\
        );

    \I__1848\ : InMux
    port map (
            O => \N__8751\,
            I => \N__8728\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__8748\,
            I => \N__8723\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__8743\,
            I => \N__8723\
        );

    \I__1845\ : Span4Mux_v
    port map (
            O => \N__8738\,
            I => \N__8720\
        );

    \I__1844\ : InMux
    port map (
            O => \N__8737\,
            I => \N__8717\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__8734\,
            I => \U712_CHIP_RAM.N_314\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__8731\,
            I => \U712_CHIP_RAM.N_314\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__8728\,
            I => \U712_CHIP_RAM.N_314\
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__8723\,
            I => \U712_CHIP_RAM.N_314\
        );

    \I__1839\ : Odrv4
    port map (
            O => \N__8720\,
            I => \U712_CHIP_RAM.N_314\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__8717\,
            I => \U712_CHIP_RAM.N_314\
        );

    \I__1837\ : IoInMux
    port map (
            O => \N__8704\,
            I => \N__8701\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__8701\,
            I => \N__8698\
        );

    \I__1835\ : Span12Mux_s0_v
    port map (
            O => \N__8698\,
            I => \N__8695\
        );

    \I__1834\ : Span12Mux_v
    port map (
            O => \N__8695\,
            I => \N__8692\
        );

    \I__1833\ : Odrv12
    port map (
            O => \N__8692\,
            I => \CMA_c_2\
        );

    \I__1832\ : InMux
    port map (
            O => \N__8689\,
            I => \N__8686\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__8686\,
            I => \N__8683\
        );

    \I__1830\ : Odrv4
    port map (
            O => \N__8683\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__1829\ : InMux
    port map (
            O => \N__8680\,
            I => \N__8674\
        );

    \I__1828\ : InMux
    port map (
            O => \N__8679\,
            I => \N__8674\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8674\,
            I => \N__8669\
        );

    \I__1826\ : InMux
    port map (
            O => \N__8673\,
            I => \N__8666\
        );

    \I__1825\ : InMux
    port map (
            O => \N__8672\,
            I => \N__8663\
        );

    \I__1824\ : Span4Mux_h
    port map (
            O => \N__8669\,
            I => \N__8658\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__8666\,
            I => \N__8658\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__8663\,
            I => \N__8655\
        );

    \I__1821\ : Span4Mux_v
    port map (
            O => \N__8658\,
            I => \N__8652\
        );

    \I__1820\ : Span4Mux_h
    port map (
            O => \N__8655\,
            I => \N__8649\
        );

    \I__1819\ : Sp12to4
    port map (
            O => \N__8652\,
            I => \N__8646\
        );

    \I__1818\ : Sp12to4
    port map (
            O => \N__8649\,
            I => \N__8643\
        );

    \I__1817\ : Span12Mux_h
    port map (
            O => \N__8646\,
            I => \N__8640\
        );

    \I__1816\ : Span12Mux_v
    port map (
            O => \N__8643\,
            I => \N__8637\
        );

    \I__1815\ : Span12Mux_v
    port map (
            O => \N__8640\,
            I => \N__8634\
        );

    \I__1814\ : Span12Mux_h
    port map (
            O => \N__8637\,
            I => \N__8631\
        );

    \I__1813\ : Odrv12
    port map (
            O => \N__8634\,
            I => \DRA_c_9\
        );

    \I__1812\ : Odrv12
    port map (
            O => \N__8631\,
            I => \DRA_c_9\
        );

    \I__1811\ : InMux
    port map (
            O => \N__8626\,
            I => \N__8617\
        );

    \I__1810\ : InMux
    port map (
            O => \N__8625\,
            I => \N__8617\
        );

    \I__1809\ : InMux
    port map (
            O => \N__8624\,
            I => \N__8617\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__8617\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__8614\,
            I => \U712_CYCLE_TERM.N_455_cascade_\
        );

    \I__1806\ : InMux
    port map (
            O => \N__8611\,
            I => \N__8606\
        );

    \I__1805\ : InMux
    port map (
            O => \N__8610\,
            I => \N__8602\
        );

    \I__1804\ : CascadeMux
    port map (
            O => \N__8609\,
            I => \N__8599\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__8606\,
            I => \N__8596\
        );

    \I__1802\ : InMux
    port map (
            O => \N__8605\,
            I => \N__8593\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__8602\,
            I => \N__8590\
        );

    \I__1800\ : InMux
    port map (
            O => \N__8599\,
            I => \N__8587\
        );

    \I__1799\ : Span4Mux_h
    port map (
            O => \N__8596\,
            I => \N__8580\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__8593\,
            I => \N__8580\
        );

    \I__1797\ : Span4Mux_v
    port map (
            O => \N__8590\,
            I => \N__8580\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__8587\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1795\ : Odrv4
    port map (
            O => \N__8580\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1794\ : InMux
    port map (
            O => \N__8575\,
            I => \N__8569\
        );

    \I__1793\ : InMux
    port map (
            O => \N__8574\,
            I => \N__8562\
        );

    \I__1792\ : InMux
    port map (
            O => \N__8573\,
            I => \N__8562\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8572\,
            I => \N__8562\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__8569\,
            I => \REG_TACK\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__8562\,
            I => \REG_TACK\
        );

    \I__1788\ : CascadeMux
    port map (
            O => \N__8557\,
            I => \N__8554\
        );

    \I__1787\ : InMux
    port map (
            O => \N__8554\,
            I => \N__8548\
        );

    \I__1786\ : InMux
    port map (
            O => \N__8553\,
            I => \N__8543\
        );

    \I__1785\ : InMux
    port map (
            O => \N__8552\,
            I => \N__8543\
        );

    \I__1784\ : InMux
    port map (
            O => \N__8551\,
            I => \N__8540\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__8548\,
            I => \N__8535\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__8543\,
            I => \N__8535\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__8540\,
            I => \CPU_TACKm\
        );

    \I__1780\ : Odrv12
    port map (
            O => \N__8535\,
            I => \CPU_TACKm\
        );

    \I__1779\ : InMux
    port map (
            O => \N__8530\,
            I => \N__8527\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__8527\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1777\ : CascadeMux
    port map (
            O => \N__8524\,
            I => \N__8519\
        );

    \I__1776\ : InMux
    port map (
            O => \N__8523\,
            I => \N__8516\
        );

    \I__1775\ : InMux
    port map (
            O => \N__8522\,
            I => \N__8513\
        );

    \I__1774\ : InMux
    port map (
            O => \N__8519\,
            I => \N__8510\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__8516\,
            I => \N__8507\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__8513\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__8510\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__1770\ : Odrv12
    port map (
            O => \N__8507\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__1769\ : InMux
    port map (
            O => \N__8500\,
            I => \N__8497\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__8497\,
            I => \N__8489\
        );

    \I__1767\ : InMux
    port map (
            O => \N__8496\,
            I => \N__8486\
        );

    \I__1766\ : InMux
    port map (
            O => \N__8495\,
            I => \N__8483\
        );

    \I__1765\ : InMux
    port map (
            O => \N__8494\,
            I => \N__8476\
        );

    \I__1764\ : InMux
    port map (
            O => \N__8493\,
            I => \N__8476\
        );

    \I__1763\ : InMux
    port map (
            O => \N__8492\,
            I => \N__8476\
        );

    \I__1762\ : Odrv4
    port map (
            O => \N__8489\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__8486\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__8483\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__8476\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__1758\ : InMux
    port map (
            O => \N__8467\,
            I => \N__8464\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__8464\,
            I => \N__8460\
        );

    \I__1756\ : InMux
    port map (
            O => \N__8463\,
            I => \N__8457\
        );

    \I__1755\ : Odrv4
    port map (
            O => \N__8460\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__8457\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__1753\ : IoInMux
    port map (
            O => \N__8452\,
            I => \N__8449\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__8449\,
            I => \N__8446\
        );

    \I__1751\ : Span12Mux_s9_v
    port map (
            O => \N__8446\,
            I => \N__8443\
        );

    \I__1750\ : Span12Mux_h
    port map (
            O => \N__8443\,
            I => \N__8440\
        );

    \I__1749\ : Odrv12
    port map (
            O => \N__8440\,
            I => \CASn_c\
        );

    \I__1748\ : InMux
    port map (
            O => \N__8437\,
            I => \N__8434\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__8434\,
            I => \U712_CHIP_RAM.N_361\
        );

    \I__1746\ : InMux
    port map (
            O => \N__8431\,
            I => \N__8428\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__8428\,
            I => \U712_CHIP_RAM.N_367\
        );

    \I__1744\ : IoInMux
    port map (
            O => \N__8425\,
            I => \N__8422\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__8422\,
            I => \N__8419\
        );

    \I__1742\ : IoSpan4Mux
    port map (
            O => \N__8419\,
            I => \N__8416\
        );

    \I__1741\ : Span4Mux_s2_h
    port map (
            O => \N__8416\,
            I => \N__8413\
        );

    \I__1740\ : Sp12to4
    port map (
            O => \N__8413\,
            I => \N__8410\
        );

    \I__1739\ : Span12Mux_h
    port map (
            O => \N__8410\,
            I => \N__8407\
        );

    \I__1738\ : Odrv12
    port map (
            O => \N__8407\,
            I => \CMA_c_5\
        );

    \I__1737\ : IoInMux
    port map (
            O => \N__8404\,
            I => \N__8401\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__8401\,
            I => \N__8398\
        );

    \I__1735\ : IoSpan4Mux
    port map (
            O => \N__8398\,
            I => \N__8395\
        );

    \I__1734\ : Span4Mux_s3_v
    port map (
            O => \N__8395\,
            I => \N__8392\
        );

    \I__1733\ : Span4Mux_v
    port map (
            O => \N__8392\,
            I => \N__8389\
        );

    \I__1732\ : Span4Mux_h
    port map (
            O => \N__8389\,
            I => \N__8386\
        );

    \I__1731\ : Odrv4
    port map (
            O => \N__8386\,
            I => \CMA_c_10\
        );

    \I__1730\ : InMux
    port map (
            O => \N__8383\,
            I => \N__8380\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__8380\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__1728\ : InMux
    port map (
            O => \N__8377\,
            I => \N__8374\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__8374\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__1726\ : InMux
    port map (
            O => \N__8371\,
            I => \N__8368\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__8368\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\
        );

    \I__1724\ : IoInMux
    port map (
            O => \N__8365\,
            I => \N__8362\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__8362\,
            I => \N__8359\
        );

    \I__1722\ : Span12Mux_s5_v
    port map (
            O => \N__8359\,
            I => \N__8356\
        );

    \I__1721\ : Odrv12
    port map (
            O => \N__8356\,
            I => \CMA_c_1\
        );

    \I__1720\ : IoInMux
    port map (
            O => \N__8353\,
            I => \N__8350\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__8350\,
            I => \N__8347\
        );

    \I__1718\ : IoSpan4Mux
    port map (
            O => \N__8347\,
            I => \N__8344\
        );

    \I__1717\ : Span4Mux_s2_h
    port map (
            O => \N__8344\,
            I => \N__8341\
        );

    \I__1716\ : Sp12to4
    port map (
            O => \N__8341\,
            I => \N__8338\
        );

    \I__1715\ : Span12Mux_s9_h
    port map (
            O => \N__8338\,
            I => \N__8335\
        );

    \I__1714\ : Span12Mux_v
    port map (
            O => \N__8335\,
            I => \N__8332\
        );

    \I__1713\ : Odrv12
    port map (
            O => \N__8332\,
            I => \CMA_c_3\
        );

    \I__1712\ : IoInMux
    port map (
            O => \N__8329\,
            I => \N__8326\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__8326\,
            I => \N__8323\
        );

    \I__1710\ : IoSpan4Mux
    port map (
            O => \N__8323\,
            I => \N__8320\
        );

    \I__1709\ : Span4Mux_s3_h
    port map (
            O => \N__8320\,
            I => \N__8317\
        );

    \I__1708\ : Sp12to4
    port map (
            O => \N__8317\,
            I => \N__8314\
        );

    \I__1707\ : Span12Mux_h
    port map (
            O => \N__8314\,
            I => \N__8311\
        );

    \I__1706\ : Odrv12
    port map (
            O => \N__8311\,
            I => \CMA_c_4\
        );

    \I__1705\ : InMux
    port map (
            O => \N__8308\,
            I => \N__8305\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__8305\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__1703\ : IoInMux
    port map (
            O => \N__8302\,
            I => \N__8299\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__8299\,
            I => \N__8296\
        );

    \I__1701\ : IoSpan4Mux
    port map (
            O => \N__8296\,
            I => \N__8293\
        );

    \I__1700\ : Span4Mux_s2_h
    port map (
            O => \N__8293\,
            I => \N__8290\
        );

    \I__1699\ : Sp12to4
    port map (
            O => \N__8290\,
            I => \N__8287\
        );

    \I__1698\ : Span12Mux_s11_h
    port map (
            O => \N__8287\,
            I => \N__8284\
        );

    \I__1697\ : Span12Mux_v
    port map (
            O => \N__8284\,
            I => \N__8281\
        );

    \I__1696\ : Odrv12
    port map (
            O => \N__8281\,
            I => \CMA_c_6\
        );

    \I__1695\ : CascadeMux
    port map (
            O => \N__8278\,
            I => \N__8275\
        );

    \I__1694\ : InMux
    port map (
            O => \N__8275\,
            I => \N__8272\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__8272\,
            I => \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\
        );

    \I__1692\ : InMux
    port map (
            O => \N__8269\,
            I => \N__8266\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__8266\,
            I => \U712_CHIP_RAM.N_190\
        );

    \I__1690\ : InMux
    port map (
            O => \N__8263\,
            I => \N__8260\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__8260\,
            I => \N__8257\
        );

    \I__1688\ : Sp12to4
    port map (
            O => \N__8257\,
            I => \N__8254\
        );

    \I__1687\ : Span12Mux_v
    port map (
            O => \N__8254\,
            I => \N__8251\
        );

    \I__1686\ : Span12Mux_h
    port map (
            O => \N__8251\,
            I => \N__8248\
        );

    \I__1685\ : Odrv12
    port map (
            O => \N__8248\,
            I => \A_c_13\
        );

    \I__1684\ : InMux
    port map (
            O => \N__8245\,
            I => \N__8242\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__8242\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__8239\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\
        );

    \I__1681\ : InMux
    port map (
            O => \N__8236\,
            I => \N__8233\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__8233\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__1679\ : InMux
    port map (
            O => \N__8230\,
            I => \N__8227\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__8227\,
            I => \N__8224\
        );

    \I__1677\ : Odrv4
    port map (
            O => \N__8224\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__8221\,
            I => \N__8217\
        );

    \I__1675\ : InMux
    port map (
            O => \N__8220\,
            I => \N__8214\
        );

    \I__1674\ : InMux
    port map (
            O => \N__8217\,
            I => \N__8211\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__8214\,
            I => \N__8206\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__8211\,
            I => \N__8206\
        );

    \I__1671\ : Odrv12
    port map (
            O => \N__8206\,
            I => \DBRn_c_i\
        );

    \I__1670\ : InMux
    port map (
            O => \N__8203\,
            I => \N__8200\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__8200\,
            I => \N__8196\
        );

    \I__1668\ : InMux
    port map (
            O => \N__8199\,
            I => \N__8193\
        );

    \I__1667\ : Span4Mux_h
    port map (
            O => \N__8196\,
            I => \N__8190\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__8193\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__1665\ : Odrv4
    port map (
            O => \N__8190\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__1664\ : InMux
    port map (
            O => \N__8185\,
            I => \N__8182\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__8182\,
            I => \U712_CYCLE_TERM.N_332\
        );

    \I__1662\ : InMux
    port map (
            O => \N__8179\,
            I => \N__8174\
        );

    \I__1661\ : InMux
    port map (
            O => \N__8178\,
            I => \N__8171\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__8177\,
            I => \N__8168\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__8174\,
            I => \N__8163\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__8171\,
            I => \N__8163\
        );

    \I__1657\ : InMux
    port map (
            O => \N__8168\,
            I => \N__8160\
        );

    \I__1656\ : Span4Mux_v
    port map (
            O => \N__8163\,
            I => \N__8153\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__8160\,
            I => \N__8153\
        );

    \I__1654\ : InMux
    port map (
            O => \N__8159\,
            I => \N__8148\
        );

    \I__1653\ : InMux
    port map (
            O => \N__8158\,
            I => \N__8148\
        );

    \I__1652\ : Odrv4
    port map (
            O => \N__8153\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__8148\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1650\ : InMux
    port map (
            O => \N__8143\,
            I => \N__8140\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__8140\,
            I => \N__8135\
        );

    \I__1648\ : InMux
    port map (
            O => \N__8139\,
            I => \N__8132\
        );

    \I__1647\ : InMux
    port map (
            O => \N__8138\,
            I => \N__8127\
        );

    \I__1646\ : Span4Mux_v
    port map (
            O => \N__8135\,
            I => \N__8122\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__8132\,
            I => \N__8122\
        );

    \I__1644\ : InMux
    port map (
            O => \N__8131\,
            I => \N__8117\
        );

    \I__1643\ : InMux
    port map (
            O => \N__8130\,
            I => \N__8117\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__8127\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1641\ : Odrv4
    port map (
            O => \N__8122\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__8117\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1639\ : CascadeMux
    port map (
            O => \N__8110\,
            I => \U712_CHIP_RAM.N_314_cascade_\
        );

    \I__1638\ : InMux
    port map (
            O => \N__8107\,
            I => \N__8104\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__8104\,
            I => \N__8101\
        );

    \I__1636\ : Span4Mux_v
    port map (
            O => \N__8101\,
            I => \N__8098\
        );

    \I__1635\ : Span4Mux_v
    port map (
            O => \N__8098\,
            I => \N__8095\
        );

    \I__1634\ : Sp12to4
    port map (
            O => \N__8095\,
            I => \N__8092\
        );

    \I__1633\ : Span12Mux_h
    port map (
            O => \N__8092\,
            I => \N__8089\
        );

    \I__1632\ : Odrv12
    port map (
            O => \N__8089\,
            I => \A_c_14\
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__8086\,
            I => \N__8083\
        );

    \I__1630\ : InMux
    port map (
            O => \N__8083\,
            I => \N__8080\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__8080\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\
        );

    \I__1628\ : InMux
    port map (
            O => \N__8077\,
            I => \N__8074\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__8074\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i\
        );

    \I__1626\ : InMux
    port map (
            O => \N__8071\,
            I => \N__8068\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__8068\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\
        );

    \I__1624\ : InMux
    port map (
            O => \N__8065\,
            I => \N__8062\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__8062\,
            I => \N__8059\
        );

    \I__1622\ : Span12Mux_h
    port map (
            O => \N__8059\,
            I => \N__8056\
        );

    \I__1621\ : Odrv12
    port map (
            O => \N__8056\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\
        );

    \I__1620\ : InMux
    port map (
            O => \N__8053\,
            I => \N__8050\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__8050\,
            I => \N__8047\
        );

    \I__1618\ : Odrv4
    port map (
            O => \N__8047\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__1617\ : InMux
    port map (
            O => \N__8044\,
            I => \N__8041\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__8041\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__1615\ : InMux
    port map (
            O => \N__8038\,
            I => \N__8031\
        );

    \I__1614\ : InMux
    port map (
            O => \N__8037\,
            I => \N__8025\
        );

    \I__1613\ : InMux
    port map (
            O => \N__8036\,
            I => \N__8025\
        );

    \I__1612\ : InMux
    port map (
            O => \N__8035\,
            I => \N__8022\
        );

    \I__1611\ : InMux
    port map (
            O => \N__8034\,
            I => \N__8019\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__8031\,
            I => \N__8016\
        );

    \I__1609\ : InMux
    port map (
            O => \N__8030\,
            I => \N__8013\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__8025\,
            I => \N__8010\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__8022\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__8019\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1605\ : Odrv4
    port map (
            O => \N__8016\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__8013\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1603\ : Odrv4
    port map (
            O => \N__8010\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1602\ : CascadeMux
    port map (
            O => \N__7999\,
            I => \U712_REG_SM.N_373_cascade_\
        );

    \I__1601\ : InMux
    port map (
            O => \N__7996\,
            I => \N__7993\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__7993\,
            I => \U712_REG_SM.N_130\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7990\,
            I => \N__7986\
        );

    \I__1598\ : InMux
    port map (
            O => \N__7989\,
            I => \N__7982\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__7986\,
            I => \N__7979\
        );

    \I__1596\ : InMux
    port map (
            O => \N__7985\,
            I => \N__7976\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__7982\,
            I => \U712_REG_SM.un1_REGENn_0_sqmuxa_0\
        );

    \I__1594\ : Odrv4
    port map (
            O => \N__7979\,
            I => \U712_REG_SM.un1_REGENn_0_sqmuxa_0\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__7976\,
            I => \U712_REG_SM.un1_REGENn_0_sqmuxa_0\
        );

    \I__1592\ : InMux
    port map (
            O => \N__7969\,
            I => \N__7966\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__7966\,
            I => \N__7963\
        );

    \I__1590\ : Odrv4
    port map (
            O => \N__7963\,
            I => \U712_CHIP_RAM.N_335\
        );

    \I__1589\ : CascadeMux
    port map (
            O => \N__7960\,
            I => \N__7952\
        );

    \I__1588\ : InMux
    port map (
            O => \N__7959\,
            I => \N__7948\
        );

    \I__1587\ : InMux
    port map (
            O => \N__7958\,
            I => \N__7945\
        );

    \I__1586\ : InMux
    port map (
            O => \N__7957\,
            I => \N__7937\
        );

    \I__1585\ : CascadeMux
    port map (
            O => \N__7956\,
            I => \N__7932\
        );

    \I__1584\ : InMux
    port map (
            O => \N__7955\,
            I => \N__7929\
        );

    \I__1583\ : InMux
    port map (
            O => \N__7952\,
            I => \N__7926\
        );

    \I__1582\ : InMux
    port map (
            O => \N__7951\,
            I => \N__7923\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__7948\,
            I => \N__7918\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__7945\,
            I => \N__7918\
        );

    \I__1579\ : InMux
    port map (
            O => \N__7944\,
            I => \N__7909\
        );

    \I__1578\ : InMux
    port map (
            O => \N__7943\,
            I => \N__7909\
        );

    \I__1577\ : InMux
    port map (
            O => \N__7942\,
            I => \N__7909\
        );

    \I__1576\ : InMux
    port map (
            O => \N__7941\,
            I => \N__7909\
        );

    \I__1575\ : InMux
    port map (
            O => \N__7940\,
            I => \N__7906\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__7937\,
            I => \N__7903\
        );

    \I__1573\ : InMux
    port map (
            O => \N__7936\,
            I => \N__7896\
        );

    \I__1572\ : InMux
    port map (
            O => \N__7935\,
            I => \N__7896\
        );

    \I__1571\ : InMux
    port map (
            O => \N__7932\,
            I => \N__7896\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__7929\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__7926\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__7923\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1567\ : Odrv4
    port map (
            O => \N__7918\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__7909\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__7906\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1564\ : Odrv4
    port map (
            O => \N__7903\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__7896\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1562\ : IoInMux
    port map (
            O => \N__7879\,
            I => \N__7876\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__7876\,
            I => \N__7873\
        );

    \I__1560\ : Span12Mux_s11_v
    port map (
            O => \N__7873\,
            I => \N__7870\
        );

    \I__1559\ : Span12Mux_h
    port map (
            O => \N__7870\,
            I => \N__7867\
        );

    \I__1558\ : Odrv12
    port map (
            O => \N__7867\,
            I => \ASn_c\
        );

    \I__1557\ : CEMux
    port map (
            O => \N__7864\,
            I => \N__7861\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__7861\,
            I => \N__7858\
        );

    \I__1555\ : Span4Mux_h
    port map (
            O => \N__7858\,
            I => \N__7855\
        );

    \I__1554\ : Odrv4
    port map (
            O => \N__7855\,
            I => \U712_REG_SM.un1_REGENn_0_sqmuxa_0_0_0\
        );

    \I__1553\ : IoInMux
    port map (
            O => \N__7852\,
            I => \N__7849\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__7849\,
            I => \N__7846\
        );

    \I__1551\ : IoSpan4Mux
    port map (
            O => \N__7846\,
            I => \N__7843\
        );

    \I__1550\ : Span4Mux_s3_v
    port map (
            O => \N__7843\,
            I => \N__7840\
        );

    \I__1549\ : Span4Mux_v
    port map (
            O => \N__7840\,
            I => \N__7837\
        );

    \I__1548\ : Odrv4
    port map (
            O => \N__7837\,
            I => \N_165_i\
        );

    \I__1547\ : IoInMux
    port map (
            O => \N__7834\,
            I => \N__7830\
        );

    \I__1546\ : InMux
    port map (
            O => \N__7833\,
            I => \N__7827\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__7830\,
            I => \N__7824\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__7827\,
            I => \N__7821\
        );

    \I__1543\ : Span12Mux_s8_v
    port map (
            O => \N__7824\,
            I => \N__7818\
        );

    \I__1542\ : Span4Mux_h
    port map (
            O => \N__7821\,
            I => \N__7815\
        );

    \I__1541\ : Odrv12
    port map (
            O => \N__7818\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1540\ : Odrv4
    port map (
            O => \N__7815\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1539\ : IoInMux
    port map (
            O => \N__7810\,
            I => \N__7807\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7807\,
            I => \N__7804\
        );

    \I__1537\ : Span4Mux_s2_v
    port map (
            O => \N__7804\,
            I => \N__7801\
        );

    \I__1536\ : Span4Mux_v
    port map (
            O => \N__7801\,
            I => \N__7798\
        );

    \I__1535\ : Sp12to4
    port map (
            O => \N__7798\,
            I => \N__7795\
        );

    \I__1534\ : Span12Mux_h
    port map (
            O => \N__7795\,
            I => \N__7792\
        );

    \I__1533\ : Odrv12
    port map (
            O => \N__7792\,
            I => \RASn_c\
        );

    \I__1532\ : IoInMux
    port map (
            O => \N__7789\,
            I => \N__7786\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__7786\,
            I => \N__7783\
        );

    \I__1530\ : IoSpan4Mux
    port map (
            O => \N__7783\,
            I => \N__7780\
        );

    \I__1529\ : IoSpan4Mux
    port map (
            O => \N__7780\,
            I => \N__7777\
        );

    \I__1528\ : Sp12to4
    port map (
            O => \N__7777\,
            I => \N__7774\
        );

    \I__1527\ : Span12Mux_s7_v
    port map (
            O => \N__7774\,
            I => \N__7771\
        );

    \I__1526\ : Span12Mux_h
    port map (
            O => \N__7771\,
            I => \N__7768\
        );

    \I__1525\ : Odrv12
    port map (
            O => \N__7768\,
            I => \WEn_c\
        );

    \I__1524\ : InMux
    port map (
            O => \N__7765\,
            I => \N__7762\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__7762\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\
        );

    \I__1522\ : InMux
    port map (
            O => \N__7759\,
            I => \N__7753\
        );

    \I__1521\ : InMux
    port map (
            O => \N__7758\,
            I => \N__7753\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__7753\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1519\ : IoInMux
    port map (
            O => \N__7750\,
            I => \N__7746\
        );

    \I__1518\ : IoInMux
    port map (
            O => \N__7749\,
            I => \N__7743\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__7746\,
            I => \N__7739\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__7743\,
            I => \N__7736\
        );

    \I__1515\ : IoInMux
    port map (
            O => \N__7742\,
            I => \N__7733\
        );

    \I__1514\ : Span4Mux_s1_v
    port map (
            O => \N__7739\,
            I => \N__7730\
        );

    \I__1513\ : IoSpan4Mux
    port map (
            O => \N__7736\,
            I => \N__7727\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__7733\,
            I => \N__7724\
        );

    \I__1511\ : Span4Mux_v
    port map (
            O => \N__7730\,
            I => \N__7721\
        );

    \I__1510\ : Span4Mux_s2_v
    port map (
            O => \N__7727\,
            I => \N__7718\
        );

    \I__1509\ : Span4Mux_s2_h
    port map (
            O => \N__7724\,
            I => \N__7715\
        );

    \I__1508\ : Sp12to4
    port map (
            O => \N__7721\,
            I => \N__7712\
        );

    \I__1507\ : Span4Mux_v
    port map (
            O => \N__7718\,
            I => \N__7709\
        );

    \I__1506\ : Span4Mux_h
    port map (
            O => \N__7715\,
            I => \N__7706\
        );

    \I__1505\ : Span12Mux_h
    port map (
            O => \N__7712\,
            I => \N__7703\
        );

    \I__1504\ : Sp12to4
    port map (
            O => \N__7709\,
            I => \N__7700\
        );

    \I__1503\ : Sp12to4
    port map (
            O => \N__7706\,
            I => \N__7697\
        );

    \I__1502\ : Span12Mux_v
    port map (
            O => \N__7703\,
            I => \N__7689\
        );

    \I__1501\ : Span12Mux_v
    port map (
            O => \N__7700\,
            I => \N__7689\
        );

    \I__1500\ : Span12Mux_v
    port map (
            O => \N__7697\,
            I => \N__7689\
        );

    \I__1499\ : InMux
    port map (
            O => \N__7696\,
            I => \N__7686\
        );

    \I__1498\ : Odrv12
    port map (
            O => \N__7689\,
            I => \TACK_EN\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__7686\,
            I => \TACK_EN\
        );

    \I__1496\ : CascadeMux
    port map (
            O => \N__7681\,
            I => \N__7677\
        );

    \I__1495\ : CascadeMux
    port map (
            O => \N__7680\,
            I => \N__7674\
        );

    \I__1494\ : InMux
    port map (
            O => \N__7677\,
            I => \N__7670\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7674\,
            I => \N__7667\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7673\,
            I => \N__7664\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__7670\,
            I => \N__7661\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__7667\,
            I => \U712_REG_SM.N_328\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__7664\,
            I => \U712_REG_SM.N_328\
        );

    \I__1488\ : Odrv4
    port map (
            O => \N__7661\,
            I => \U712_REG_SM.N_328\
        );

    \I__1487\ : CascadeMux
    port map (
            O => \N__7654\,
            I => \N__7651\
        );

    \I__1486\ : InMux
    port map (
            O => \N__7651\,
            I => \N__7648\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__7648\,
            I => \U712_REG_SM.N_406\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7645\,
            I => \N__7642\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__7642\,
            I => \N__7637\
        );

    \I__1482\ : InMux
    port map (
            O => \N__7641\,
            I => \N__7633\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7640\,
            I => \N__7629\
        );

    \I__1480\ : Span4Mux_h
    port map (
            O => \N__7637\,
            I => \N__7626\
        );

    \I__1479\ : InMux
    port map (
            O => \N__7636\,
            I => \N__7623\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__7633\,
            I => \N__7620\
        );

    \I__1477\ : InMux
    port map (
            O => \N__7632\,
            I => \N__7617\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__7629\,
            I => \N__7614\
        );

    \I__1475\ : Odrv4
    port map (
            O => \N__7626\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__7623\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1473\ : Odrv4
    port map (
            O => \N__7620\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__7617\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1471\ : Odrv4
    port map (
            O => \N__7614\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1470\ : CascadeMux
    port map (
            O => \N__7603\,
            I => \U712_REG_SM.N_330_cascade_\
        );

    \I__1469\ : InMux
    port map (
            O => \N__7600\,
            I => \N__7597\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__7597\,
            I => \N__7591\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7596\,
            I => \N__7588\
        );

    \I__1466\ : InMux
    port map (
            O => \N__7595\,
            I => \N__7583\
        );

    \I__1465\ : InMux
    port map (
            O => \N__7594\,
            I => \N__7583\
        );

    \I__1464\ : Odrv4
    port map (
            O => \N__7591\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__7588\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__7583\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1461\ : InMux
    port map (
            O => \N__7576\,
            I => \N__7573\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__7573\,
            I => \U712_REG_SM.STATE_COUNTc_0_0\
        );

    \I__1459\ : InMux
    port map (
            O => \N__7570\,
            I => \N__7563\
        );

    \I__1458\ : InMux
    port map (
            O => \N__7569\,
            I => \N__7558\
        );

    \I__1457\ : InMux
    port map (
            O => \N__7568\,
            I => \N__7558\
        );

    \I__1456\ : InMux
    port map (
            O => \N__7567\,
            I => \N__7555\
        );

    \I__1455\ : InMux
    port map (
            O => \N__7566\,
            I => \N__7552\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__7563\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__7558\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__7555\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__7552\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1450\ : CascadeMux
    port map (
            O => \N__7543\,
            I => \N__7539\
        );

    \I__1449\ : InMux
    port map (
            O => \N__7542\,
            I => \N__7528\
        );

    \I__1448\ : InMux
    port map (
            O => \N__7539\,
            I => \N__7528\
        );

    \I__1447\ : CascadeMux
    port map (
            O => \N__7538\,
            I => \N__7523\
        );

    \I__1446\ : CascadeMux
    port map (
            O => \N__7537\,
            I => \N__7519\
        );

    \I__1445\ : InMux
    port map (
            O => \N__7536\,
            I => \N__7516\
        );

    \I__1444\ : CascadeMux
    port map (
            O => \N__7535\,
            I => \N__7513\
        );

    \I__1443\ : CascadeMux
    port map (
            O => \N__7534\,
            I => \N__7510\
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__7533\,
            I => \N__7507\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__7528\,
            I => \N__7503\
        );

    \I__1440\ : InMux
    port map (
            O => \N__7527\,
            I => \N__7498\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7526\,
            I => \N__7498\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7523\,
            I => \N__7493\
        );

    \I__1437\ : InMux
    port map (
            O => \N__7522\,
            I => \N__7493\
        );

    \I__1436\ : InMux
    port map (
            O => \N__7519\,
            I => \N__7490\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__7516\,
            I => \N__7487\
        );

    \I__1434\ : InMux
    port map (
            O => \N__7513\,
            I => \N__7484\
        );

    \I__1433\ : InMux
    port map (
            O => \N__7510\,
            I => \N__7477\
        );

    \I__1432\ : InMux
    port map (
            O => \N__7507\,
            I => \N__7477\
        );

    \I__1431\ : InMux
    port map (
            O => \N__7506\,
            I => \N__7477\
        );

    \I__1430\ : Odrv12
    port map (
            O => \N__7503\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__7498\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__7493\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__7490\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1426\ : Odrv4
    port map (
            O => \N__7487\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__7484\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__7477\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1423\ : InMux
    port map (
            O => \N__7462\,
            I => \N__7459\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__7459\,
            I => \U712_REG_SM.N_373\
        );

    \I__1421\ : InMux
    port map (
            O => \N__7456\,
            I => \N__7452\
        );

    \I__1420\ : InMux
    port map (
            O => \N__7455\,
            I => \N__7449\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__7452\,
            I => \N__7446\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__7449\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__1417\ : Odrv4
    port map (
            O => \N__7446\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__1416\ : InMux
    port map (
            O => \N__7441\,
            I => \N__7438\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__7438\,
            I => \N__7435\
        );

    \I__1414\ : Span4Mux_h
    port map (
            O => \N__7435\,
            I => \N__7431\
        );

    \I__1413\ : InMux
    port map (
            O => \N__7434\,
            I => \N__7428\
        );

    \I__1412\ : Span4Mux_v
    port map (
            O => \N__7431\,
            I => \N__7423\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__7428\,
            I => \N__7423\
        );

    \I__1410\ : Span4Mux_v
    port map (
            O => \N__7423\,
            I => \N__7419\
        );

    \I__1409\ : InMux
    port map (
            O => \N__7422\,
            I => \N__7416\
        );

    \I__1408\ : Odrv4
    port map (
            O => \N__7419\,
            I => \REG_CYCLEm\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__7416\,
            I => \REG_CYCLEm\
        );

    \I__1406\ : IoInMux
    port map (
            O => \N__7411\,
            I => \N__7408\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__7408\,
            I => \N__7405\
        );

    \I__1404\ : Span4Mux_s1_v
    port map (
            O => \N__7405\,
            I => \N__7402\
        );

    \I__1403\ : Span4Mux_v
    port map (
            O => \N__7402\,
            I => \N__7399\
        );

    \I__1402\ : Sp12to4
    port map (
            O => \N__7399\,
            I => \N__7396\
        );

    \I__1401\ : Span12Mux_s10_h
    port map (
            O => \N__7396\,
            I => \N__7393\
        );

    \I__1400\ : Span12Mux_v
    port map (
            O => \N__7393\,
            I => \N__7390\
        );

    \I__1399\ : Odrv12
    port map (
            O => \N__7390\,
            I => \N_167_i\
        );

    \I__1398\ : InMux
    port map (
            O => \N__7387\,
            I => \N__7381\
        );

    \I__1397\ : InMux
    port map (
            O => \N__7386\,
            I => \N__7376\
        );

    \I__1396\ : InMux
    port map (
            O => \N__7385\,
            I => \N__7376\
        );

    \I__1395\ : InMux
    port map (
            O => \N__7384\,
            I => \N__7373\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__7381\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__7376\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__7373\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1391\ : InMux
    port map (
            O => \N__7366\,
            I => \N__7363\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__7363\,
            I => \U712_CHIP_RAM.N_321\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__7360\,
            I => \U712_CHIP_RAM.N_321_cascade_\
        );

    \I__1388\ : InMux
    port map (
            O => \N__7357\,
            I => \N__7353\
        );

    \I__1387\ : InMux
    port map (
            O => \N__7356\,
            I => \N__7350\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__7353\,
            I => \U712_CHIP_RAM.N_20_0\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__7350\,
            I => \U712_CHIP_RAM.N_20_0\
        );

    \I__1384\ : CascadeMux
    port map (
            O => \N__7345\,
            I => \N__7341\
        );

    \I__1383\ : CascadeMux
    port map (
            O => \N__7344\,
            I => \N__7337\
        );

    \I__1382\ : InMux
    port map (
            O => \N__7341\,
            I => \N__7332\
        );

    \I__1381\ : InMux
    port map (
            O => \N__7340\,
            I => \N__7329\
        );

    \I__1380\ : InMux
    port map (
            O => \N__7337\,
            I => \N__7326\
        );

    \I__1379\ : InMux
    port map (
            O => \N__7336\,
            I => \N__7322\
        );

    \I__1378\ : InMux
    port map (
            O => \N__7335\,
            I => \N__7319\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__7332\,
            I => \N__7316\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__7329\,
            I => \N__7313\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__7326\,
            I => \N__7310\
        );

    \I__1374\ : InMux
    port map (
            O => \N__7325\,
            I => \N__7299\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__7322\,
            I => \N__7294\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__7319\,
            I => \N__7294\
        );

    \I__1371\ : Span4Mux_h
    port map (
            O => \N__7316\,
            I => \N__7291\
        );

    \I__1370\ : Span4Mux_h
    port map (
            O => \N__7313\,
            I => \N__7286\
        );

    \I__1369\ : Span4Mux_h
    port map (
            O => \N__7310\,
            I => \N__7286\
        );

    \I__1368\ : InMux
    port map (
            O => \N__7309\,
            I => \N__7281\
        );

    \I__1367\ : InMux
    port map (
            O => \N__7308\,
            I => \N__7281\
        );

    \I__1366\ : InMux
    port map (
            O => \N__7307\,
            I => \N__7278\
        );

    \I__1365\ : InMux
    port map (
            O => \N__7306\,
            I => \N__7273\
        );

    \I__1364\ : InMux
    port map (
            O => \N__7305\,
            I => \N__7273\
        );

    \I__1363\ : InMux
    port map (
            O => \N__7304\,
            I => \N__7266\
        );

    \I__1362\ : InMux
    port map (
            O => \N__7303\,
            I => \N__7266\
        );

    \I__1361\ : InMux
    port map (
            O => \N__7302\,
            I => \N__7266\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__7299\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1359\ : Odrv4
    port map (
            O => \N__7294\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1358\ : Odrv4
    port map (
            O => \N__7291\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1357\ : Odrv4
    port map (
            O => \N__7286\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__7281\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__7278\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__7273\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__7266\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1352\ : CascadeMux
    port map (
            O => \N__7249\,
            I => \U712_CHIP_RAM.m77_0_a2_0_2_cascade_\
        );

    \I__1351\ : CascadeMux
    port map (
            O => \N__7246\,
            I => \N__7240\
        );

    \I__1350\ : InMux
    port map (
            O => \N__7245\,
            I => \N__7237\
        );

    \I__1349\ : InMux
    port map (
            O => \N__7244\,
            I => \N__7232\
        );

    \I__1348\ : InMux
    port map (
            O => \N__7243\,
            I => \N__7232\
        );

    \I__1347\ : InMux
    port map (
            O => \N__7240\,
            I => \N__7229\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__7237\,
            I => \N__7226\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__7232\,
            I => \N__7223\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__7229\,
            I => \N__7218\
        );

    \I__1343\ : Span4Mux_h
    port map (
            O => \N__7226\,
            I => \N__7215\
        );

    \I__1342\ : Span4Mux_v
    port map (
            O => \N__7223\,
            I => \N__7212\
        );

    \I__1341\ : InMux
    port map (
            O => \N__7222\,
            I => \N__7209\
        );

    \I__1340\ : InMux
    port map (
            O => \N__7221\,
            I => \N__7206\
        );

    \I__1339\ : Odrv4
    port map (
            O => \N__7218\,
            I => \U712_CHIP_RAM.N_307\
        );

    \I__1338\ : Odrv4
    port map (
            O => \N__7215\,
            I => \U712_CHIP_RAM.N_307\
        );

    \I__1337\ : Odrv4
    port map (
            O => \N__7212\,
            I => \U712_CHIP_RAM.N_307\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__7209\,
            I => \U712_CHIP_RAM.N_307\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__7206\,
            I => \U712_CHIP_RAM.N_307\
        );

    \I__1334\ : CascadeMux
    port map (
            O => \N__7195\,
            I => \N__7191\
        );

    \I__1333\ : InMux
    port map (
            O => \N__7194\,
            I => \N__7182\
        );

    \I__1332\ : InMux
    port map (
            O => \N__7191\,
            I => \N__7179\
        );

    \I__1331\ : CascadeMux
    port map (
            O => \N__7190\,
            I => \N__7176\
        );

    \I__1330\ : InMux
    port map (
            O => \N__7189\,
            I => \N__7173\
        );

    \I__1329\ : CascadeMux
    port map (
            O => \N__7188\,
            I => \N__7163\
        );

    \I__1328\ : InMux
    port map (
            O => \N__7187\,
            I => \N__7156\
        );

    \I__1327\ : InMux
    port map (
            O => \N__7186\,
            I => \N__7151\
        );

    \I__1326\ : InMux
    port map (
            O => \N__7185\,
            I => \N__7151\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__7182\,
            I => \N__7148\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__7179\,
            I => \N__7145\
        );

    \I__1323\ : InMux
    port map (
            O => \N__7176\,
            I => \N__7142\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__7173\,
            I => \N__7139\
        );

    \I__1321\ : InMux
    port map (
            O => \N__7172\,
            I => \N__7136\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__7171\,
            I => \N__7133\
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__7170\,
            I => \N__7130\
        );

    \I__1318\ : InMux
    port map (
            O => \N__7169\,
            I => \N__7120\
        );

    \I__1317\ : InMux
    port map (
            O => \N__7168\,
            I => \N__7117\
        );

    \I__1316\ : InMux
    port map (
            O => \N__7167\,
            I => \N__7110\
        );

    \I__1315\ : InMux
    port map (
            O => \N__7166\,
            I => \N__7110\
        );

    \I__1314\ : InMux
    port map (
            O => \N__7163\,
            I => \N__7110\
        );

    \I__1313\ : InMux
    port map (
            O => \N__7162\,
            I => \N__7107\
        );

    \I__1312\ : InMux
    port map (
            O => \N__7161\,
            I => \N__7102\
        );

    \I__1311\ : InMux
    port map (
            O => \N__7160\,
            I => \N__7102\
        );

    \I__1310\ : InMux
    port map (
            O => \N__7159\,
            I => \N__7099\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__7156\,
            I => \N__7096\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__7151\,
            I => \N__7091\
        );

    \I__1307\ : Span4Mux_h
    port map (
            O => \N__7148\,
            I => \N__7091\
        );

    \I__1306\ : Span4Mux_v
    port map (
            O => \N__7145\,
            I => \N__7082\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__7142\,
            I => \N__7082\
        );

    \I__1304\ : Span4Mux_v
    port map (
            O => \N__7139\,
            I => \N__7082\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__7136\,
            I => \N__7082\
        );

    \I__1302\ : InMux
    port map (
            O => \N__7133\,
            I => \N__7075\
        );

    \I__1301\ : InMux
    port map (
            O => \N__7130\,
            I => \N__7075\
        );

    \I__1300\ : InMux
    port map (
            O => \N__7129\,
            I => \N__7075\
        );

    \I__1299\ : InMux
    port map (
            O => \N__7128\,
            I => \N__7062\
        );

    \I__1298\ : InMux
    port map (
            O => \N__7127\,
            I => \N__7062\
        );

    \I__1297\ : InMux
    port map (
            O => \N__7126\,
            I => \N__7062\
        );

    \I__1296\ : InMux
    port map (
            O => \N__7125\,
            I => \N__7062\
        );

    \I__1295\ : InMux
    port map (
            O => \N__7124\,
            I => \N__7062\
        );

    \I__1294\ : InMux
    port map (
            O => \N__7123\,
            I => \N__7062\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__7120\,
            I => \N__7051\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__7117\,
            I => \N__7051\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__7110\,
            I => \N__7051\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__7107\,
            I => \N__7051\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__7102\,
            I => \N__7051\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__7099\,
            I => \N__7048\
        );

    \I__1287\ : Odrv12
    port map (
            O => \N__7096\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1286\ : Odrv4
    port map (
            O => \N__7091\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1285\ : Odrv4
    port map (
            O => \N__7082\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__7075\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__7062\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1282\ : Odrv4
    port map (
            O => \N__7051\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1281\ : Odrv4
    port map (
            O => \N__7048\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1280\ : InMux
    port map (
            O => \N__7033\,
            I => \N__7027\
        );

    \I__1279\ : InMux
    port map (
            O => \N__7032\,
            I => \N__7013\
        );

    \I__1278\ : InMux
    port map (
            O => \N__7031\,
            I => \N__7008\
        );

    \I__1277\ : InMux
    port map (
            O => \N__7030\,
            I => \N__7008\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__7027\,
            I => \N__7005\
        );

    \I__1275\ : InMux
    port map (
            O => \N__7026\,
            I => \N__6990\
        );

    \I__1274\ : InMux
    port map (
            O => \N__7025\,
            I => \N__6990\
        );

    \I__1273\ : InMux
    port map (
            O => \N__7024\,
            I => \N__6990\
        );

    \I__1272\ : InMux
    port map (
            O => \N__7023\,
            I => \N__6990\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__7022\,
            I => \N__6987\
        );

    \I__1270\ : CascadeMux
    port map (
            O => \N__7021\,
            I => \N__6979\
        );

    \I__1269\ : InMux
    port map (
            O => \N__7020\,
            I => \N__6972\
        );

    \I__1268\ : InMux
    port map (
            O => \N__7019\,
            I => \N__6972\
        );

    \I__1267\ : InMux
    port map (
            O => \N__7018\,
            I => \N__6969\
        );

    \I__1266\ : InMux
    port map (
            O => \N__7017\,
            I => \N__6966\
        );

    \I__1265\ : InMux
    port map (
            O => \N__7016\,
            I => \N__6963\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__7013\,
            I => \N__6960\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__7008\,
            I => \N__6955\
        );

    \I__1262\ : Span4Mux_h
    port map (
            O => \N__7005\,
            I => \N__6955\
        );

    \I__1261\ : InMux
    port map (
            O => \N__7004\,
            I => \N__6948\
        );

    \I__1260\ : InMux
    port map (
            O => \N__7003\,
            I => \N__6948\
        );

    \I__1259\ : InMux
    port map (
            O => \N__7002\,
            I => \N__6948\
        );

    \I__1258\ : InMux
    port map (
            O => \N__7001\,
            I => \N__6945\
        );

    \I__1257\ : InMux
    port map (
            O => \N__7000\,
            I => \N__6940\
        );

    \I__1256\ : InMux
    port map (
            O => \N__6999\,
            I => \N__6940\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__6990\,
            I => \N__6937\
        );

    \I__1254\ : InMux
    port map (
            O => \N__6987\,
            I => \N__6926\
        );

    \I__1253\ : InMux
    port map (
            O => \N__6986\,
            I => \N__6926\
        );

    \I__1252\ : InMux
    port map (
            O => \N__6985\,
            I => \N__6926\
        );

    \I__1251\ : InMux
    port map (
            O => \N__6984\,
            I => \N__6926\
        );

    \I__1250\ : InMux
    port map (
            O => \N__6983\,
            I => \N__6926\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6982\,
            I => \N__6917\
        );

    \I__1248\ : InMux
    port map (
            O => \N__6979\,
            I => \N__6917\
        );

    \I__1247\ : InMux
    port map (
            O => \N__6978\,
            I => \N__6917\
        );

    \I__1246\ : InMux
    port map (
            O => \N__6977\,
            I => \N__6917\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__6972\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__6969\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__6966\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__6963\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1241\ : Odrv4
    port map (
            O => \N__6960\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1240\ : Odrv4
    port map (
            O => \N__6955\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__6948\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6945\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__6940\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1236\ : Odrv4
    port map (
            O => \N__6937\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__6926\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__6917\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1233\ : CascadeMux
    port map (
            O => \N__6892\,
            I => \N__6887\
        );

    \I__1232\ : InMux
    port map (
            O => \N__6891\,
            I => \N__6882\
        );

    \I__1231\ : InMux
    port map (
            O => \N__6890\,
            I => \N__6877\
        );

    \I__1230\ : InMux
    port map (
            O => \N__6887\,
            I => \N__6877\
        );

    \I__1229\ : InMux
    port map (
            O => \N__6886\,
            I => \N__6874\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6885\,
            I => \N__6870\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__6882\,
            I => \N__6867\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__6877\,
            I => \N__6860\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__6874\,
            I => \N__6852\
        );

    \I__1224\ : InMux
    port map (
            O => \N__6873\,
            I => \N__6849\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__6870\,
            I => \N__6846\
        );

    \I__1222\ : Span4Mux_v
    port map (
            O => \N__6867\,
            I => \N__6843\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6866\,
            I => \N__6840\
        );

    \I__1220\ : InMux
    port map (
            O => \N__6865\,
            I => \N__6833\
        );

    \I__1219\ : InMux
    port map (
            O => \N__6864\,
            I => \N__6833\
        );

    \I__1218\ : InMux
    port map (
            O => \N__6863\,
            I => \N__6833\
        );

    \I__1217\ : Span4Mux_h
    port map (
            O => \N__6860\,
            I => \N__6830\
        );

    \I__1216\ : InMux
    port map (
            O => \N__6859\,
            I => \N__6827\
        );

    \I__1215\ : InMux
    port map (
            O => \N__6858\,
            I => \N__6822\
        );

    \I__1214\ : InMux
    port map (
            O => \N__6857\,
            I => \N__6822\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6856\,
            I => \N__6819\
        );

    \I__1212\ : InMux
    port map (
            O => \N__6855\,
            I => \N__6816\
        );

    \I__1211\ : Odrv4
    port map (
            O => \N__6852\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__6849\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1209\ : Odrv4
    port map (
            O => \N__6846\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1208\ : Odrv4
    port map (
            O => \N__6843\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__6840\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__6833\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1205\ : Odrv4
    port map (
            O => \N__6830\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__6827\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__6822\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__6819\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__6816\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1200\ : CascadeMux
    port map (
            O => \N__6793\,
            I => \N__6788\
        );

    \I__1199\ : CascadeMux
    port map (
            O => \N__6792\,
            I => \N__6785\
        );

    \I__1198\ : InMux
    port map (
            O => \N__6791\,
            I => \N__6779\
        );

    \I__1197\ : InMux
    port map (
            O => \N__6788\,
            I => \N__6779\
        );

    \I__1196\ : InMux
    port map (
            O => \N__6785\,
            I => \N__6774\
        );

    \I__1195\ : InMux
    port map (
            O => \N__6784\,
            I => \N__6768\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__6779\,
            I => \N__6765\
        );

    \I__1193\ : CascadeMux
    port map (
            O => \N__6778\,
            I => \N__6761\
        );

    \I__1192\ : InMux
    port map (
            O => \N__6777\,
            I => \N__6755\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__6774\,
            I => \N__6749\
        );

    \I__1190\ : InMux
    port map (
            O => \N__6773\,
            I => \N__6746\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6772\,
            I => \N__6741\
        );

    \I__1188\ : InMux
    port map (
            O => \N__6771\,
            I => \N__6741\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__6768\,
            I => \N__6736\
        );

    \I__1186\ : Span4Mux_h
    port map (
            O => \N__6765\,
            I => \N__6736\
        );

    \I__1185\ : InMux
    port map (
            O => \N__6764\,
            I => \N__6731\
        );

    \I__1184\ : InMux
    port map (
            O => \N__6761\,
            I => \N__6731\
        );

    \I__1183\ : InMux
    port map (
            O => \N__6760\,
            I => \N__6726\
        );

    \I__1182\ : InMux
    port map (
            O => \N__6759\,
            I => \N__6726\
        );

    \I__1181\ : InMux
    port map (
            O => \N__6758\,
            I => \N__6723\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6755\,
            I => \N__6720\
        );

    \I__1179\ : InMux
    port map (
            O => \N__6754\,
            I => \N__6715\
        );

    \I__1178\ : InMux
    port map (
            O => \N__6753\,
            I => \N__6715\
        );

    \I__1177\ : InMux
    port map (
            O => \N__6752\,
            I => \N__6712\
        );

    \I__1176\ : Odrv4
    port map (
            O => \N__6749\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6746\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__6741\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1173\ : Odrv4
    port map (
            O => \N__6736\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__6731\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__6726\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__6723\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1169\ : Odrv4
    port map (
            O => \N__6720\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__6715\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__6712\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1166\ : InMux
    port map (
            O => \N__6691\,
            I => \N__6688\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__6688\,
            I => \N__6685\
        );

    \I__1164\ : Span4Mux_h
    port map (
            O => \N__6685\,
            I => \N__6682\
        );

    \I__1163\ : Span4Mux_v
    port map (
            O => \N__6682\,
            I => \N__6679\
        );

    \I__1162\ : Odrv4
    port map (
            O => \N__6679\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_6\
        );

    \I__1161\ : SRMux
    port map (
            O => \N__6676\,
            I => \N__6672\
        );

    \I__1160\ : SRMux
    port map (
            O => \N__6675\,
            I => \N__6669\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__6672\,
            I => \N__6664\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__6669\,
            I => \N__6664\
        );

    \I__1157\ : Span4Mux_v
    port map (
            O => \N__6664\,
            I => \N__6661\
        );

    \I__1156\ : Odrv4
    port map (
            O => \N__6661\,
            I => \U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1\
        );

    \I__1155\ : InMux
    port map (
            O => \N__6658\,
            I => \N__6654\
        );

    \I__1154\ : InMux
    port map (
            O => \N__6657\,
            I => \N__6651\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__6654\,
            I => \N__6646\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__6651\,
            I => \N__6646\
        );

    \I__1151\ : Span4Mux_h
    port map (
            O => \N__6646\,
            I => \N__6642\
        );

    \I__1150\ : InMux
    port map (
            O => \N__6645\,
            I => \N__6639\
        );

    \I__1149\ : Odrv4
    port map (
            O => \N__6642\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__6639\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1147\ : IoInMux
    port map (
            O => \N__6634\,
            I => \N__6631\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__6631\,
            I => \N__6628\
        );

    \I__1145\ : IoSpan4Mux
    port map (
            O => \N__6628\,
            I => \N__6625\
        );

    \I__1144\ : Span4Mux_s2_v
    port map (
            O => \N__6625\,
            I => \N__6622\
        );

    \I__1143\ : Sp12to4
    port map (
            O => \N__6622\,
            I => \N__6619\
        );

    \I__1142\ : Span12Mux_s9_v
    port map (
            O => \N__6619\,
            I => \N__6616\
        );

    \I__1141\ : Odrv12
    port map (
            O => \N__6616\,
            I => \N_202_i\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6613\,
            I => \N__6610\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__6610\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1138\ : InMux
    port map (
            O => \N__6607\,
            I => \N__6604\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__6604\,
            I => \N__6599\
        );

    \I__1136\ : InMux
    port map (
            O => \N__6603\,
            I => \N__6596\
        );

    \I__1135\ : InMux
    port map (
            O => \N__6602\,
            I => \N__6593\
        );

    \I__1134\ : Odrv12
    port map (
            O => \N__6599\,
            I => \U712_CHIP_RAM.N_305\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__6596\,
            I => \U712_CHIP_RAM.N_305\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__6593\,
            I => \U712_CHIP_RAM.N_305\
        );

    \I__1131\ : CascadeMux
    port map (
            O => \N__6586\,
            I => \U712_CHIP_RAM.m123_i_2_cascade_\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6583\,
            I => \N__6580\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6580\,
            I => \N__6577\
        );

    \I__1128\ : Span4Mux_v
    port map (
            O => \N__6577\,
            I => \N__6574\
        );

    \I__1127\ : Span4Mux_v
    port map (
            O => \N__6574\,
            I => \N__6571\
        );

    \I__1126\ : Sp12to4
    port map (
            O => \N__6571\,
            I => \N__6568\
        );

    \I__1125\ : Span12Mux_h
    port map (
            O => \N__6568\,
            I => \N__6565\
        );

    \I__1124\ : Odrv12
    port map (
            O => \N__6565\,
            I => \A_c_15\
        );

    \I__1123\ : InMux
    port map (
            O => \N__6562\,
            I => \N__6559\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__6559\,
            I => \N__6556\
        );

    \I__1121\ : Odrv12
    port map (
            O => \N__6556\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\
        );

    \I__1120\ : CascadeMux
    port map (
            O => \N__6553\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\
        );

    \I__1119\ : InMux
    port map (
            O => \N__6550\,
            I => \N__6547\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__6547\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_2_0\
        );

    \I__1117\ : InMux
    port map (
            O => \N__6544\,
            I => \N__6541\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__6541\,
            I => \U712_CHIP_RAM.N_390\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6538\,
            I => \N__6535\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__6535\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_2_3\
        );

    \I__1113\ : IoInMux
    port map (
            O => \N__6532\,
            I => \N__6529\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__6529\,
            I => \N__6526\
        );

    \I__1111\ : IoSpan4Mux
    port map (
            O => \N__6526\,
            I => \N__6523\
        );

    \I__1110\ : Span4Mux_s2_v
    port map (
            O => \N__6523\,
            I => \N__6519\
        );

    \I__1109\ : InMux
    port map (
            O => \N__6522\,
            I => \N__6516\
        );

    \I__1108\ : Sp12to4
    port map (
            O => \N__6519\,
            I => \N__6513\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__6516\,
            I => \N__6510\
        );

    \I__1106\ : Span12Mux_s8_v
    port map (
            O => \N__6513\,
            I => \N__6507\
        );

    \I__1105\ : Span4Mux_v
    port map (
            O => \N__6510\,
            I => \N__6504\
        );

    \I__1104\ : Span12Mux_h
    port map (
            O => \N__6507\,
            I => \N__6501\
        );

    \I__1103\ : Sp12to4
    port map (
            O => \N__6504\,
            I => \N__6498\
        );

    \I__1102\ : Span12Mux_v
    port map (
            O => \N__6501\,
            I => \N__6495\
        );

    \I__1101\ : Span12Mux_h
    port map (
            O => \N__6498\,
            I => \N__6492\
        );

    \I__1100\ : Odrv12
    port map (
            O => \N__6495\,
            I => \A_c_11\
        );

    \I__1099\ : Odrv12
    port map (
            O => \N__6492\,
            I => \A_c_11\
        );

    \I__1098\ : InMux
    port map (
            O => \N__6487\,
            I => \N__6484\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__6484\,
            I => \N__6481\
        );

    \I__1096\ : Odrv12
    port map (
            O => \N__6481\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\
        );

    \I__1095\ : InMux
    port map (
            O => \N__6478\,
            I => \N__6475\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__6475\,
            I => \N__6472\
        );

    \I__1093\ : Span12Mux_v
    port map (
            O => \N__6472\,
            I => \N__6469\
        );

    \I__1092\ : Span12Mux_h
    port map (
            O => \N__6469\,
            I => \N__6466\
        );

    \I__1091\ : Odrv12
    port map (
            O => \N__6466\,
            I => \A_c_3\
        );

    \I__1090\ : InMux
    port map (
            O => \N__6463\,
            I => \N__6460\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__6460\,
            I => \N__6457\
        );

    \I__1088\ : Odrv4
    port map (
            O => \N__6457\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\
        );

    \I__1087\ : InMux
    port map (
            O => \N__6454\,
            I => \N__6451\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__6451\,
            I => \N__6448\
        );

    \I__1085\ : Span4Mux_v
    port map (
            O => \N__6448\,
            I => \N__6445\
        );

    \I__1084\ : Span4Mux_v
    port map (
            O => \N__6445\,
            I => \N__6442\
        );

    \I__1083\ : Sp12to4
    port map (
            O => \N__6442\,
            I => \N__6439\
        );

    \I__1082\ : Span12Mux_h
    port map (
            O => \N__6439\,
            I => \N__6436\
        );

    \I__1081\ : Odrv12
    port map (
            O => \N__6436\,
            I => \A_c_5\
        );

    \I__1080\ : InMux
    port map (
            O => \N__6433\,
            I => \N__6430\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__6430\,
            I => \N__6427\
        );

    \I__1078\ : Odrv4
    port map (
            O => \N__6427\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\
        );

    \I__1077\ : InMux
    port map (
            O => \N__6424\,
            I => \N__6421\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__6421\,
            I => \N__6418\
        );

    \I__1075\ : Span12Mux_v
    port map (
            O => \N__6418\,
            I => \N__6415\
        );

    \I__1074\ : Span12Mux_h
    port map (
            O => \N__6415\,
            I => \N__6412\
        );

    \I__1073\ : Odrv12
    port map (
            O => \N__6412\,
            I => \A_c_6\
        );

    \I__1072\ : CEMux
    port map (
            O => \N__6409\,
            I => \N__6404\
        );

    \I__1071\ : CEMux
    port map (
            O => \N__6408\,
            I => \N__6401\
        );

    \I__1070\ : CEMux
    port map (
            O => \N__6407\,
            I => \N__6398\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__6404\,
            I => \N__6395\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__6401\,
            I => \N__6392\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__6398\,
            I => \N__6389\
        );

    \I__1066\ : Span4Mux_h
    port map (
            O => \N__6395\,
            I => \N__6386\
        );

    \I__1065\ : Span4Mux_h
    port map (
            O => \N__6392\,
            I => \N__6383\
        );

    \I__1064\ : Span4Mux_h
    port map (
            O => \N__6389\,
            I => \N__6380\
        );

    \I__1063\ : Odrv4
    port map (
            O => \N__6386\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\
        );

    \I__1062\ : Odrv4
    port map (
            O => \N__6383\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\
        );

    \I__1061\ : Odrv4
    port map (
            O => \N__6380\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\
        );

    \I__1060\ : InMux
    port map (
            O => \N__6373\,
            I => \N__6370\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__6370\,
            I => \N__6366\
        );

    \I__1058\ : InMux
    port map (
            O => \N__6369\,
            I => \N__6363\
        );

    \I__1057\ : Span4Mux_h
    port map (
            O => \N__6366\,
            I => \N__6360\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__6363\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_4\
        );

    \I__1055\ : Odrv4
    port map (
            O => \N__6360\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_4\
        );

    \I__1054\ : InMux
    port map (
            O => \N__6355\,
            I => \U712_CHIP_RAM.un3_DBR_COUNT_cry_3\
        );

    \I__1053\ : InMux
    port map (
            O => \N__6352\,
            I => \N__6349\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__6349\,
            I => \N__6345\
        );

    \I__1051\ : InMux
    port map (
            O => \N__6348\,
            I => \N__6342\
        );

    \I__1050\ : Span4Mux_v
    port map (
            O => \N__6345\,
            I => \N__6339\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__6342\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_5\
        );

    \I__1048\ : Odrv4
    port map (
            O => \N__6339\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_5\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6334\,
            I => \U712_CHIP_RAM.un3_DBR_COUNT_cry_4\
        );

    \I__1046\ : InMux
    port map (
            O => \N__6331\,
            I => \N__6328\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__6328\,
            I => \N__6324\
        );

    \I__1044\ : InMux
    port map (
            O => \N__6327\,
            I => \N__6321\
        );

    \I__1043\ : Span4Mux_v
    port map (
            O => \N__6324\,
            I => \N__6318\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__6321\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_6\
        );

    \I__1041\ : Odrv4
    port map (
            O => \N__6318\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_6\
        );

    \I__1040\ : InMux
    port map (
            O => \N__6313\,
            I => \U712_CHIP_RAM.un3_DBR_COUNT_cry_5\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6310\,
            I => \U712_CHIP_RAM.un3_DBR_COUNT_cry_6\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6307\,
            I => \N__6304\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__6304\,
            I => \N__6301\
        );

    \I__1036\ : Span12Mux_v
    port map (
            O => \N__6301\,
            I => \N__6298\
        );

    \I__1035\ : Span12Mux_h
    port map (
            O => \N__6298\,
            I => \N__6295\
        );

    \I__1034\ : Odrv12
    port map (
            O => \N__6295\,
            I => \A_c_12\
        );

    \I__1033\ : IoInMux
    port map (
            O => \N__6292\,
            I => \N__6289\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__6289\,
            I => \N__6286\
        );

    \I__1031\ : Span4Mux_s0_v
    port map (
            O => \N__6286\,
            I => \N__6283\
        );

    \I__1030\ : Span4Mux_v
    port map (
            O => \N__6283\,
            I => \N__6280\
        );

    \I__1029\ : Span4Mux_v
    port map (
            O => \N__6280\,
            I => \N__6277\
        );

    \I__1028\ : Sp12to4
    port map (
            O => \N__6277\,
            I => \N__6273\
        );

    \I__1027\ : InMux
    port map (
            O => \N__6276\,
            I => \N__6270\
        );

    \I__1026\ : Span12Mux_h
    port map (
            O => \N__6273\,
            I => \N__6267\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__6270\,
            I => \N__6264\
        );

    \I__1024\ : Span12Mux_v
    port map (
            O => \N__6267\,
            I => \N__6259\
        );

    \I__1023\ : Span12Mux_h
    port map (
            O => \N__6264\,
            I => \N__6259\
        );

    \I__1022\ : Odrv12
    port map (
            O => \N__6259\,
            I => \A_c_10\
        );

    \I__1021\ : InMux
    port map (
            O => \N__6256\,
            I => \N__6252\
        );

    \I__1020\ : InMux
    port map (
            O => \N__6255\,
            I => \N__6249\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__6252\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_3\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__6249\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_3\
        );

    \I__1017\ : InMux
    port map (
            O => \N__6244\,
            I => \N__6240\
        );

    \I__1016\ : InMux
    port map (
            O => \N__6243\,
            I => \N__6237\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__6240\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_2\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__6237\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_2\
        );

    \I__1013\ : CascadeMux
    port map (
            O => \N__6232\,
            I => \N__6227\
        );

    \I__1012\ : InMux
    port map (
            O => \N__6231\,
            I => \N__6224\
        );

    \I__1011\ : InMux
    port map (
            O => \N__6230\,
            I => \N__6221\
        );

    \I__1010\ : InMux
    port map (
            O => \N__6227\,
            I => \N__6218\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__6224\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_1\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__6221\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_1\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__6218\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_1\
        );

    \I__1006\ : InMux
    port map (
            O => \N__6211\,
            I => \N__6207\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6210\,
            I => \N__6204\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__6207\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_7\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__6204\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_7\
        );

    \I__1002\ : InMux
    port map (
            O => \N__6199\,
            I => \N__6196\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__6196\,
            I => \N__6193\
        );

    \I__1000\ : Odrv4
    port map (
            O => \N__6193\,
            I => \U712_CHIP_RAM.m93_i_a2_5\
        );

    \I__999\ : SRMux
    port map (
            O => \N__6190\,
            I => \N__6187\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__6187\,
            I => \N__6183\
        );

    \I__997\ : InMux
    port map (
            O => \N__6186\,
            I => \N__6180\
        );

    \I__996\ : Span4Mux_v
    port map (
            O => \N__6183\,
            I => \N__6177\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__6180\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__994\ : Odrv4
    port map (
            O => \N__6177\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__993\ : InMux
    port map (
            O => \N__6172\,
            I => \N__6169\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__6169\,
            I => \N__6164\
        );

    \I__991\ : InMux
    port map (
            O => \N__6168\,
            I => \N__6161\
        );

    \I__990\ : InMux
    port map (
            O => \N__6167\,
            I => \N__6158\
        );

    \I__989\ : Odrv4
    port map (
            O => \N__6164\,
            I => \U712_CHIP_RAM.N_304\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__6161\,
            I => \U712_CHIP_RAM.N_304\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__6158\,
            I => \U712_CHIP_RAM.N_304\
        );

    \I__986\ : InMux
    port map (
            O => \N__6151\,
            I => \N__6148\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__6148\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__984\ : InMux
    port map (
            O => \N__6145\,
            I => \N__6142\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__6142\,
            I => \N__6137\
        );

    \I__982\ : InMux
    port map (
            O => \N__6141\,
            I => \N__6132\
        );

    \I__981\ : InMux
    port map (
            O => \N__6140\,
            I => \N__6132\
        );

    \I__980\ : Odrv4
    port map (
            O => \N__6137\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__6132\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__978\ : IoInMux
    port map (
            O => \N__6127\,
            I => \N__6124\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__6124\,
            I => \N__6120\
        );

    \I__976\ : IoInMux
    port map (
            O => \N__6123\,
            I => \N__6117\
        );

    \I__975\ : IoSpan4Mux
    port map (
            O => \N__6120\,
            I => \N__6114\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__6117\,
            I => \N__6110\
        );

    \I__973\ : Sp12to4
    port map (
            O => \N__6114\,
            I => \N__6107\
        );

    \I__972\ : IoInMux
    port map (
            O => \N__6113\,
            I => \N__6104\
        );

    \I__971\ : Span4Mux_s1_h
    port map (
            O => \N__6110\,
            I => \N__6101\
        );

    \I__970\ : Span12Mux_s7_v
    port map (
            O => \N__6107\,
            I => \N__6098\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__6104\,
            I => \N__6095\
        );

    \I__968\ : Span4Mux_h
    port map (
            O => \N__6101\,
            I => \N__6092\
        );

    \I__967\ : Span12Mux_h
    port map (
            O => \N__6098\,
            I => \N__6089\
        );

    \I__966\ : Span12Mux_s7_v
    port map (
            O => \N__6095\,
            I => \N__6086\
        );

    \I__965\ : Sp12to4
    port map (
            O => \N__6092\,
            I => \N__6083\
        );

    \I__964\ : Span12Mux_v
    port map (
            O => \N__6089\,
            I => \N__6075\
        );

    \I__963\ : Span12Mux_v
    port map (
            O => \N__6086\,
            I => \N__6075\
        );

    \I__962\ : Span12Mux_v
    port map (
            O => \N__6083\,
            I => \N__6075\
        );

    \I__961\ : InMux
    port map (
            O => \N__6082\,
            I => \N__6072\
        );

    \I__960\ : Odrv12
    port map (
            O => \N__6075\,
            I => \TACK_OUTn\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__6072\,
            I => \TACK_OUTn\
        );

    \I__958\ : InMux
    port map (
            O => \N__6067\,
            I => \N__6064\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__6064\,
            I => \N__6061\
        );

    \I__956\ : Odrv4
    port map (
            O => \N__6061\,
            I => \U712_REG_SM.N_404\
        );

    \I__955\ : IoInMux
    port map (
            O => \N__6058\,
            I => \N__6055\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__6055\,
            I => \N__6052\
        );

    \I__953\ : IoSpan4Mux
    port map (
            O => \N__6052\,
            I => \N__6049\
        );

    \I__952\ : Span4Mux_s0_v
    port map (
            O => \N__6049\,
            I => \N__6046\
        );

    \I__951\ : Sp12to4
    port map (
            O => \N__6046\,
            I => \N__6043\
        );

    \I__950\ : Span12Mux_v
    port map (
            O => \N__6043\,
            I => \N__6039\
        );

    \I__949\ : InMux
    port map (
            O => \N__6042\,
            I => \N__6036\
        );

    \I__948\ : Odrv12
    port map (
            O => \N__6039\,
            I => \LDSn_c\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__6036\,
            I => \LDSn_c\
        );

    \I__946\ : IoInMux
    port map (
            O => \N__6031\,
            I => \N__6028\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__6028\,
            I => \N__6025\
        );

    \I__944\ : IoSpan4Mux
    port map (
            O => \N__6025\,
            I => \N__6022\
        );

    \I__943\ : Span4Mux_s3_h
    port map (
            O => \N__6022\,
            I => \N__6019\
        );

    \I__942\ : Span4Mux_v
    port map (
            O => \N__6019\,
            I => \N__6015\
        );

    \I__941\ : InMux
    port map (
            O => \N__6018\,
            I => \N__6012\
        );

    \I__940\ : Span4Mux_h
    port map (
            O => \N__6015\,
            I => \N__6009\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__6012\,
            I => \N__6006\
        );

    \I__938\ : Sp12to4
    port map (
            O => \N__6009\,
            I => \N__6003\
        );

    \I__937\ : Span4Mux_v
    port map (
            O => \N__6006\,
            I => \N__6000\
        );

    \I__936\ : Span12Mux_h
    port map (
            O => \N__6003\,
            I => \N__5995\
        );

    \I__935\ : Sp12to4
    port map (
            O => \N__6000\,
            I => \N__5995\
        );

    \I__934\ : Span12Mux_h
    port map (
            O => \N__5995\,
            I => \N__5992\
        );

    \I__933\ : Odrv12
    port map (
            O => \N__5992\,
            I => \C3_c\
        );

    \I__932\ : InMux
    port map (
            O => \N__5989\,
            I => \N__5986\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__5986\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__930\ : InMux
    port map (
            O => \N__5983\,
            I => \N__5980\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__5980\,
            I => \U712_REG_SM.N_459\
        );

    \I__928\ : IoInMux
    port map (
            O => \N__5977\,
            I => \N__5974\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__5974\,
            I => \N__5971\
        );

    \I__926\ : IoSpan4Mux
    port map (
            O => \N__5971\,
            I => \N__5968\
        );

    \I__925\ : IoSpan4Mux
    port map (
            O => \N__5968\,
            I => \N__5965\
        );

    \I__924\ : Span4Mux_s3_v
    port map (
            O => \N__5965\,
            I => \N__5962\
        );

    \I__923\ : Sp12to4
    port map (
            O => \N__5962\,
            I => \N__5958\
        );

    \I__922\ : CascadeMux
    port map (
            O => \N__5961\,
            I => \N__5955\
        );

    \I__921\ : Span12Mux_s11_v
    port map (
            O => \N__5958\,
            I => \N__5952\
        );

    \I__920\ : InMux
    port map (
            O => \N__5955\,
            I => \N__5949\
        );

    \I__919\ : Odrv12
    port map (
            O => \N__5952\,
            I => \UDSn_c\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__5949\,
            I => \UDSn_c\
        );

    \I__917\ : InMux
    port map (
            O => \N__5944\,
            I => \N__5941\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__5941\,
            I => \N__5935\
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__5940\,
            I => \N__5932\
        );

    \I__914\ : InMux
    port map (
            O => \N__5939\,
            I => \N__5927\
        );

    \I__913\ : InMux
    port map (
            O => \N__5938\,
            I => \N__5927\
        );

    \I__912\ : Span4Mux_h
    port map (
            O => \N__5935\,
            I => \N__5924\
        );

    \I__911\ : InMux
    port map (
            O => \N__5932\,
            I => \N__5921\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__5927\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_0\
        );

    \I__909\ : Odrv4
    port map (
            O => \N__5924\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_0\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__5921\,
            I => \U712_CHIP_RAM.DBR_COUNTZ0Z_0\
        );

    \I__907\ : InMux
    port map (
            O => \N__5914\,
            I => \U712_CHIP_RAM.un3_DBR_COUNT_cry_1\
        );

    \I__906\ : InMux
    port map (
            O => \N__5911\,
            I => \U712_CHIP_RAM.un3_DBR_COUNT_cry_2\
        );

    \I__905\ : InMux
    port map (
            O => \N__5908\,
            I => \N__5902\
        );

    \I__904\ : InMux
    port map (
            O => \N__5907\,
            I => \N__5902\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5902\,
            I => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\
        );

    \I__902\ : CascadeMux
    port map (
            O => \N__5899\,
            I => \U712_REG_SM.N_410_cascade_\
        );

    \I__901\ : InMux
    port map (
            O => \N__5896\,
            I => \N__5893\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__5893\,
            I => \U712_REG_SM.N_331\
        );

    \I__899\ : InMux
    port map (
            O => \N__5890\,
            I => \N__5886\
        );

    \I__898\ : IoInMux
    port map (
            O => \N__5889\,
            I => \N__5883\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__5886\,
            I => \N__5880\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__5883\,
            I => \N__5877\
        );

    \I__895\ : Span4Mux_v
    port map (
            O => \N__5880\,
            I => \N__5874\
        );

    \I__894\ : IoSpan4Mux
    port map (
            O => \N__5877\,
            I => \N__5871\
        );

    \I__893\ : Sp12to4
    port map (
            O => \N__5874\,
            I => \N__5868\
        );

    \I__892\ : IoSpan4Mux
    port map (
            O => \N__5871\,
            I => \N__5865\
        );

    \I__891\ : Span12Mux_h
    port map (
            O => \N__5868\,
            I => \N__5862\
        );

    \I__890\ : IoSpan4Mux
    port map (
            O => \N__5865\,
            I => \N__5859\
        );

    \I__889\ : Odrv12
    port map (
            O => \N__5862\,
            I => \C1_c\
        );

    \I__888\ : Odrv4
    port map (
            O => \N__5859\,
            I => \C1_c\
        );

    \I__887\ : InMux
    port map (
            O => \N__5854\,
            I => \N__5848\
        );

    \I__886\ : InMux
    port map (
            O => \N__5853\,
            I => \N__5848\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5848\,
            I => \N__5845\
        );

    \I__884\ : Span4Mux_h
    port map (
            O => \N__5845\,
            I => \N__5842\
        );

    \I__883\ : Odrv4
    port map (
            O => \N__5842\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\
        );

    \I__882\ : InMux
    port map (
            O => \N__5839\,
            I => \N__5835\
        );

    \I__881\ : InMux
    port map (
            O => \N__5838\,
            I => \N__5832\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__5835\,
            I => \U712_CHIP_RAM.N_435\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__5832\,
            I => \U712_CHIP_RAM.N_435\
        );

    \I__878\ : InMux
    port map (
            O => \N__5827\,
            I => \N__5824\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__5824\,
            I => \N__5821\
        );

    \I__876\ : Odrv4
    port map (
            O => \N__5821\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__5818\,
            I => \U712_REG_SM.N_413_cascade_\
        );

    \I__874\ : IoInMux
    port map (
            O => \N__5815\,
            I => \N__5812\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__5812\,
            I => \N__5809\
        );

    \I__872\ : Span4Mux_s3_v
    port map (
            O => \N__5809\,
            I => \N__5806\
        );

    \I__871\ : Span4Mux_h
    port map (
            O => \N__5806\,
            I => \N__5803\
        );

    \I__870\ : Sp12to4
    port map (
            O => \N__5803\,
            I => \N__5797\
        );

    \I__869\ : InMux
    port map (
            O => \N__5802\,
            I => \N__5792\
        );

    \I__868\ : InMux
    port map (
            O => \N__5801\,
            I => \N__5792\
        );

    \I__867\ : InMux
    port map (
            O => \N__5800\,
            I => \N__5789\
        );

    \I__866\ : Odrv12
    port map (
            O => \N__5797\,
            I => \DBENn_c\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__5792\,
            I => \DBENn_c\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__5789\,
            I => \DBENn_c\
        );

    \I__863\ : InMux
    port map (
            O => \N__5782\,
            I => \N__5776\
        );

    \I__862\ : InMux
    port map (
            O => \N__5781\,
            I => \N__5776\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__5776\,
            I => \N__5773\
        );

    \I__860\ : Span4Mux_v
    port map (
            O => \N__5773\,
            I => \N__5768\
        );

    \I__859\ : InMux
    port map (
            O => \N__5772\,
            I => \N__5765\
        );

    \I__858\ : InMux
    port map (
            O => \N__5771\,
            I => \N__5762\
        );

    \I__857\ : Odrv4
    port map (
            O => \N__5768\,
            I => \DMA_CYCLEm\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__5765\,
            I => \DMA_CYCLEm\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__5762\,
            I => \DMA_CYCLEm\
        );

    \I__854\ : InMux
    port map (
            O => \N__5755\,
            I => \N__5752\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__5752\,
            I => \U712_REG_SM.N_308\
        );

    \I__852\ : CascadeMux
    port map (
            O => \N__5749\,
            I => \U712_REG_SM.N_308_cascade_\
        );

    \I__851\ : CascadeMux
    port map (
            O => \N__5746\,
            I => \N__5743\
        );

    \I__850\ : InMux
    port map (
            O => \N__5743\,
            I => \N__5740\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__5740\,
            I => \U712_CHIP_RAM.DBENn_7_0_0\
        );

    \I__848\ : InMux
    port map (
            O => \N__5737\,
            I => \N__5734\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__5734\,
            I => \N__5728\
        );

    \I__846\ : InMux
    port map (
            O => \N__5733\,
            I => \N__5724\
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__5732\,
            I => \N__5721\
        );

    \I__844\ : CascadeMux
    port map (
            O => \N__5731\,
            I => \N__5718\
        );

    \I__843\ : Span4Mux_v
    port map (
            O => \N__5728\,
            I => \N__5715\
        );

    \I__842\ : CascadeMux
    port map (
            O => \N__5727\,
            I => \N__5711\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__5724\,
            I => \N__5708\
        );

    \I__840\ : InMux
    port map (
            O => \N__5721\,
            I => \N__5703\
        );

    \I__839\ : InMux
    port map (
            O => \N__5718\,
            I => \N__5699\
        );

    \I__838\ : Span4Mux_h
    port map (
            O => \N__5715\,
            I => \N__5696\
        );

    \I__837\ : InMux
    port map (
            O => \N__5714\,
            I => \N__5691\
        );

    \I__836\ : InMux
    port map (
            O => \N__5711\,
            I => \N__5691\
        );

    \I__835\ : Span4Mux_h
    port map (
            O => \N__5708\,
            I => \N__5688\
        );

    \I__834\ : InMux
    port map (
            O => \N__5707\,
            I => \N__5683\
        );

    \I__833\ : InMux
    port map (
            O => \N__5706\,
            I => \N__5683\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__5703\,
            I => \N__5680\
        );

    \I__831\ : InMux
    port map (
            O => \N__5702\,
            I => \N__5677\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__5699\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__829\ : Odrv4
    port map (
            O => \N__5696\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__5691\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__827\ : Odrv4
    port map (
            O => \N__5688\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__5683\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__825\ : Odrv4
    port map (
            O => \N__5680\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__5677\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__823\ : InMux
    port map (
            O => \N__5662\,
            I => \N__5659\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__5659\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1\
        );

    \I__821\ : CascadeMux
    port map (
            O => \N__5656\,
            I => \U712_CHIP_RAM.N_344_cascade_\
        );

    \I__820\ : InMux
    port map (
            O => \N__5653\,
            I => \N__5648\
        );

    \I__819\ : InMux
    port map (
            O => \N__5652\,
            I => \N__5645\
        );

    \I__818\ : InMux
    port map (
            O => \N__5651\,
            I => \N__5642\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__5648\,
            I => \U712_CHIP_RAM.N_551\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__5645\,
            I => \U712_CHIP_RAM.N_551\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__5642\,
            I => \U712_CHIP_RAM.N_551\
        );

    \I__814\ : CascadeMux
    port map (
            O => \N__5635\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_2_0_cascade_\
        );

    \I__813\ : InMux
    port map (
            O => \N__5632\,
            I => \N__5629\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5629\,
            I => \U712_CHIP_RAM.LATCH_CLK_6\
        );

    \I__811\ : IoInMux
    port map (
            O => \N__5626\,
            I => \N__5623\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__5623\,
            I => \N__5620\
        );

    \I__809\ : IoSpan4Mux
    port map (
            O => \N__5620\,
            I => \N__5617\
        );

    \I__808\ : Span4Mux_s3_v
    port map (
            O => \N__5617\,
            I => \N__5614\
        );

    \I__807\ : Span4Mux_v
    port map (
            O => \N__5614\,
            I => \N__5611\
        );

    \I__806\ : Sp12to4
    port map (
            O => \N__5611\,
            I => \N__5608\
        );

    \I__805\ : Span12Mux_v
    port map (
            O => \N__5608\,
            I => \N__5604\
        );

    \I__804\ : InMux
    port map (
            O => \N__5607\,
            I => \N__5601\
        );

    \I__803\ : Odrv12
    port map (
            O => \N__5604\,
            I => \LATCH_CLK_c\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__5601\,
            I => \LATCH_CLK_c\
        );

    \I__801\ : InMux
    port map (
            O => \N__5596\,
            I => \N__5590\
        );

    \I__800\ : InMux
    port map (
            O => \N__5595\,
            I => \N__5590\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__5590\,
            I => \N__5586\
        );

    \I__798\ : InMux
    port map (
            O => \N__5589\,
            I => \N__5583\
        );

    \I__797\ : Span4Mux_h
    port map (
            O => \N__5586\,
            I => \N__5580\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__5583\,
            I => \N__5577\
        );

    \I__795\ : Span4Mux_v
    port map (
            O => \N__5580\,
            I => \N__5572\
        );

    \I__794\ : Span4Mux_v
    port map (
            O => \N__5577\,
            I => \N__5572\
        );

    \I__793\ : Span4Mux_h
    port map (
            O => \N__5572\,
            I => \N__5569\
        );

    \I__792\ : Sp12to4
    port map (
            O => \N__5569\,
            I => \N__5566\
        );

    \I__791\ : Odrv12
    port map (
            O => \N__5566\,
            I => \AWEn_c\
        );

    \I__790\ : InMux
    port map (
            O => \N__5563\,
            I => \N__5559\
        );

    \I__789\ : InMux
    port map (
            O => \N__5562\,
            I => \N__5556\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__5559\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5556\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\
        );

    \I__786\ : InMux
    port map (
            O => \N__5551\,
            I => \N__5548\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__5548\,
            I => \N__5545\
        );

    \I__784\ : Sp12to4
    port map (
            O => \N__5545\,
            I => \N__5542\
        );

    \I__783\ : Span12Mux_v
    port map (
            O => \N__5542\,
            I => \N__5539\
        );

    \I__782\ : Span12Mux_h
    port map (
            O => \N__5539\,
            I => \N__5536\
        );

    \I__781\ : Odrv12
    port map (
            O => \N__5536\,
            I => \A_c_20\
        );

    \I__780\ : InMux
    port map (
            O => \N__5533\,
            I => \N__5529\
        );

    \I__779\ : InMux
    port map (
            O => \N__5532\,
            I => \N__5526\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__5529\,
            I => \N__5523\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__5526\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\
        );

    \I__776\ : Odrv12
    port map (
            O => \N__5523\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\
        );

    \I__775\ : InMux
    port map (
            O => \N__5518\,
            I => \N__5515\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__5515\,
            I => \N__5510\
        );

    \I__773\ : InMux
    port map (
            O => \N__5514\,
            I => \N__5507\
        );

    \I__772\ : InMux
    port map (
            O => \N__5513\,
            I => \N__5504\
        );

    \I__771\ : Odrv4
    port map (
            O => \N__5510\,
            I => \U712_CHIP_RAM.N_194\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__5507\,
            I => \U712_CHIP_RAM.N_194\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__5504\,
            I => \U712_CHIP_RAM.N_194\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__5497\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_2_2_cascade_\
        );

    \I__767\ : InMux
    port map (
            O => \N__5494\,
            I => \N__5491\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__5491\,
            I => \U712_CHIP_RAM.N_449\
        );

    \I__765\ : InMux
    port map (
            O => \N__5488\,
            I => \N__5485\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__5485\,
            I => \N__5481\
        );

    \I__763\ : InMux
    port map (
            O => \N__5484\,
            I => \N__5478\
        );

    \I__762\ : Span4Mux_h
    port map (
            O => \N__5481\,
            I => \N__5475\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__5478\,
            I => \U712_CHIP_RAM.N_476\
        );

    \I__760\ : Odrv4
    port map (
            O => \N__5475\,
            I => \U712_CHIP_RAM.N_476\
        );

    \I__759\ : InMux
    port map (
            O => \N__5470\,
            I => \N__5467\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__5467\,
            I => \N__5464\
        );

    \I__757\ : Span4Mux_v
    port map (
            O => \N__5464\,
            I => \N__5460\
        );

    \I__756\ : InMux
    port map (
            O => \N__5463\,
            I => \N__5457\
        );

    \I__755\ : Odrv4
    port map (
            O => \N__5460\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__5457\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3\
        );

    \I__753\ : InMux
    port map (
            O => \N__5452\,
            I => \N__5449\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__5449\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__751\ : CascadeMux
    port map (
            O => \N__5446\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1_cascade_\
        );

    \I__750\ : CascadeMux
    port map (
            O => \N__5443\,
            I => \U712_CHIP_RAM.N_304_cascade_\
        );

    \I__749\ : CascadeMux
    port map (
            O => \N__5440\,
            I => \U712_CHIP_RAM.N_312_cascade_\
        );

    \I__748\ : CascadeMux
    port map (
            O => \N__5437\,
            I => \U712_CHIP_RAM.N_326_cascade_\
        );

    \I__747\ : InMux
    port map (
            O => \N__5434\,
            I => \N__5431\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__5431\,
            I => \N__5427\
        );

    \I__745\ : InMux
    port map (
            O => \N__5430\,
            I => \N__5424\
        );

    \I__744\ : Span4Mux_v
    port map (
            O => \N__5427\,
            I => \N__5417\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__5424\,
            I => \N__5414\
        );

    \I__742\ : InMux
    port map (
            O => \N__5423\,
            I => \N__5407\
        );

    \I__741\ : InMux
    port map (
            O => \N__5422\,
            I => \N__5407\
        );

    \I__740\ : InMux
    port map (
            O => \N__5421\,
            I => \N__5407\
        );

    \I__739\ : InMux
    port map (
            O => \N__5420\,
            I => \N__5404\
        );

    \I__738\ : Odrv4
    port map (
            O => \N__5417\,
            I => \U712_CHIP_RAM.N_467\
        );

    \I__737\ : Odrv4
    port map (
            O => \N__5414\,
            I => \U712_CHIP_RAM.N_467\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__5407\,
            I => \U712_CHIP_RAM.N_467\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__5404\,
            I => \U712_CHIP_RAM.N_467\
        );

    \I__734\ : InMux
    port map (
            O => \N__5395\,
            I => \N__5386\
        );

    \I__733\ : InMux
    port map (
            O => \N__5394\,
            I => \N__5386\
        );

    \I__732\ : InMux
    port map (
            O => \N__5393\,
            I => \N__5386\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__5386\,
            I => \N__5379\
        );

    \I__730\ : InMux
    port map (
            O => \N__5385\,
            I => \N__5376\
        );

    \I__729\ : InMux
    port map (
            O => \N__5384\,
            I => \N__5369\
        );

    \I__728\ : InMux
    port map (
            O => \N__5383\,
            I => \N__5369\
        );

    \I__727\ : InMux
    port map (
            O => \N__5382\,
            I => \N__5369\
        );

    \I__726\ : Odrv4
    port map (
            O => \N__5379\,
            I => \U712_CHIP_RAM.N_39\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__5376\,
            I => \U712_CHIP_RAM.N_39\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__5369\,
            I => \U712_CHIP_RAM.N_39\
        );

    \I__723\ : InMux
    port map (
            O => \N__5362\,
            I => \N__5359\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__5359\,
            I => \N__5356\
        );

    \I__721\ : Odrv4
    port map (
            O => \N__5356\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__720\ : InMux
    port map (
            O => \N__5353\,
            I => \N__5350\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__5350\,
            I => \N__5347\
        );

    \I__718\ : Odrv12
    port map (
            O => \N__5347\,
            I => \U712_CHIP_RAM.N_440\
        );

    \I__717\ : CascadeMux
    port map (
            O => \N__5344\,
            I => \U712_CHIP_RAM.N_39_cascade_\
        );

    \I__716\ : InMux
    port map (
            O => \N__5341\,
            I => \N__5338\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__5338\,
            I => \U712_CHIP_RAM.N_326\
        );

    \I__714\ : CEMux
    port map (
            O => \N__5335\,
            I => \N__5332\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__5332\,
            I => \N__5328\
        );

    \I__712\ : CEMux
    port map (
            O => \N__5331\,
            I => \N__5325\
        );

    \I__711\ : Span4Mux_h
    port map (
            O => \N__5328\,
            I => \N__5322\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__5325\,
            I => \N__5319\
        );

    \I__709\ : Odrv4
    port map (
            O => \N__5322\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__708\ : Odrv12
    port map (
            O => \N__5319\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__707\ : InMux
    port map (
            O => \N__5314\,
            I => \N__5311\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__5311\,
            I => \N__5308\
        );

    \I__705\ : Span4Mux_v
    port map (
            O => \N__5308\,
            I => \N__5305\
        );

    \I__704\ : Span4Mux_v
    port map (
            O => \N__5305\,
            I => \N__5302\
        );

    \I__703\ : Sp12to4
    port map (
            O => \N__5302\,
            I => \N__5299\
        );

    \I__702\ : Odrv12
    port map (
            O => \N__5299\,
            I => \A_c_17\
        );

    \I__701\ : CascadeMux
    port map (
            O => \N__5296\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_\
        );

    \I__700\ : InMux
    port map (
            O => \N__5293\,
            I => \N__5290\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__5290\,
            I => \N__5287\
        );

    \I__698\ : Sp12to4
    port map (
            O => \N__5287\,
            I => \N__5284\
        );

    \I__697\ : Span12Mux_v
    port map (
            O => \N__5284\,
            I => \N__5281\
        );

    \I__696\ : Span12Mux_h
    port map (
            O => \N__5281\,
            I => \N__5278\
        );

    \I__695\ : Odrv12
    port map (
            O => \N__5278\,
            I => \A_c_18\
        );

    \I__694\ : InMux
    port map (
            O => \N__5275\,
            I => \N__5272\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__5272\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\
        );

    \I__692\ : CascadeMux
    port map (
            O => \N__5269\,
            I => \N__5266\
        );

    \I__691\ : InMux
    port map (
            O => \N__5266\,
            I => \N__5263\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__5263\,
            I => \N__5260\
        );

    \I__689\ : Odrv4
    port map (
            O => \N__5260\,
            I => \U712_CHIP_RAM.N_555\
        );

    \I__688\ : CascadeMux
    port map (
            O => \N__5257\,
            I => \U712_CHIP_RAM.N_555_cascade_\
        );

    \I__687\ : InMux
    port map (
            O => \N__5254\,
            I => \N__5251\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__5251\,
            I => \U712_REG_SM.N_412\
        );

    \I__685\ : InMux
    port map (
            O => \N__5248\,
            I => \N__5245\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__5245\,
            I => \N__5242\
        );

    \I__683\ : Odrv12
    port map (
            O => \N__5242\,
            I => \U712_REG_SM.N_402\
        );

    \I__682\ : InMux
    port map (
            O => \N__5239\,
            I => \N__5235\
        );

    \I__681\ : InMux
    port map (
            O => \N__5238\,
            I => \N__5232\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__5235\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_0\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__5232\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_0\
        );

    \I__678\ : IoInMux
    port map (
            O => \N__5227\,
            I => \N__5224\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__5224\,
            I => \N__5221\
        );

    \I__676\ : Span4Mux_s3_v
    port map (
            O => \N__5221\,
            I => \N__5218\
        );

    \I__675\ : Sp12to4
    port map (
            O => \N__5218\,
            I => \N__5215\
        );

    \I__674\ : Span12Mux_s9_h
    port map (
            O => \N__5215\,
            I => \N__5210\
        );

    \I__673\ : CascadeMux
    port map (
            O => \N__5214\,
            I => \N__5207\
        );

    \I__672\ : InMux
    port map (
            O => \N__5213\,
            I => \N__5204\
        );

    \I__671\ : Span12Mux_v
    port map (
            O => \N__5210\,
            I => \N__5201\
        );

    \I__670\ : InMux
    port map (
            O => \N__5207\,
            I => \N__5198\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__5204\,
            I => \N__5195\
        );

    \I__668\ : Odrv12
    port map (
            O => \N__5201\,
            I => \REGENn_c\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__5198\,
            I => \REGENn_c\
        );

    \I__666\ : Odrv4
    port map (
            O => \N__5195\,
            I => \REGENn_c\
        );

    \I__665\ : CascadeMux
    port map (
            O => \N__5188\,
            I => \N__5184\
        );

    \I__664\ : InMux
    port map (
            O => \N__5187\,
            I => \N__5179\
        );

    \I__663\ : InMux
    port map (
            O => \N__5184\,
            I => \N__5172\
        );

    \I__662\ : InMux
    port map (
            O => \N__5183\,
            I => \N__5172\
        );

    \I__661\ : InMux
    port map (
            O => \N__5182\,
            I => \N__5172\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__5179\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__5172\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__658\ : InMux
    port map (
            O => \N__5167\,
            I => \N__5164\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__5164\,
            I => \N__5161\
        );

    \I__656\ : Odrv4
    port map (
            O => \N__5161\,
            I => \U712_REG_SM.REGENn_e_1\
        );

    \I__655\ : InMux
    port map (
            O => \N__5158\,
            I => \N__5155\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__5155\,
            I => \N__5152\
        );

    \I__653\ : Sp12to4
    port map (
            O => \N__5152\,
            I => \N__5149\
        );

    \I__652\ : Span12Mux_v
    port map (
            O => \N__5149\,
            I => \N__5146\
        );

    \I__651\ : Span12Mux_h
    port map (
            O => \N__5146\,
            I => \N__5143\
        );

    \I__650\ : Odrv12
    port map (
            O => \N__5143\,
            I => \A_c_16\
        );

    \I__649\ : CascadeMux
    port map (
            O => \N__5140\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa_cascade_\
        );

    \I__648\ : InMux
    port map (
            O => \N__5137\,
            I => \N__5134\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__5134\,
            I => \N__5131\
        );

    \I__646\ : Odrv12
    port map (
            O => \N__5131\,
            I => \U712_CHIP_RAM.N_378\
        );

    \I__645\ : CascadeMux
    port map (
            O => \N__5128\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_\
        );

    \I__644\ : CascadeMux
    port map (
            O => \N__5125\,
            I => \U712_CHIP_RAM.N_551_cascade_\
        );

    \I__643\ : InMux
    port map (
            O => \N__5122\,
            I => \N__5119\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__5119\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_0_a3_0_a2_0\
        );

    \I__641\ : IoInMux
    port map (
            O => \N__5116\,
            I => \N__5113\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__5113\,
            I => \N__5110\
        );

    \I__639\ : Span4Mux_s0_h
    port map (
            O => \N__5110\,
            I => \N__5107\
        );

    \I__638\ : Sp12to4
    port map (
            O => \N__5107\,
            I => \N__5104\
        );

    \I__637\ : Span12Mux_v
    port map (
            O => \N__5104\,
            I => \N__5101\
        );

    \I__636\ : Span12Mux_h
    port map (
            O => \N__5101\,
            I => \N__5097\
        );

    \I__635\ : InMux
    port map (
            O => \N__5100\,
            I => \N__5094\
        );

    \I__634\ : Odrv12
    port map (
            O => \N__5097\,
            I => \CLK_EN_c\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__5094\,
            I => \CLK_EN_c\
        );

    \I__632\ : InMux
    port map (
            O => \N__5089\,
            I => \N__5085\
        );

    \I__631\ : InMux
    port map (
            O => \N__5088\,
            I => \N__5082\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__5085\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__5082\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0\
        );

    \I__628\ : IoInMux
    port map (
            O => \N__5077\,
            I => \N__5074\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__5074\,
            I => \N__5071\
        );

    \I__626\ : Span4Mux_s3_v
    port map (
            O => \N__5071\,
            I => \N__5068\
        );

    \I__625\ : Span4Mux_v
    port map (
            O => \N__5068\,
            I => \N__5065\
        );

    \I__624\ : Span4Mux_v
    port map (
            O => \N__5065\,
            I => \N__5062\
        );

    \I__623\ : Span4Mux_v
    port map (
            O => \N__5062\,
            I => \N__5058\
        );

    \I__622\ : InMux
    port map (
            O => \N__5061\,
            I => \N__5055\
        );

    \I__621\ : Odrv4
    port map (
            O => \N__5058\,
            I => \DBDIR_c\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__5055\,
            I => \DBDIR_c\
        );

    \I__619\ : InMux
    port map (
            O => \N__5050\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__618\ : InMux
    port map (
            O => \N__5047\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__617\ : InMux
    port map (
            O => \N__5044\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__616\ : InMux
    port map (
            O => \N__5041\,
            I => \N__5034\
        );

    \I__615\ : InMux
    port map (
            O => \N__5040\,
            I => \N__5034\
        );

    \I__614\ : InMux
    port map (
            O => \N__5039\,
            I => \N__5029\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__5034\,
            I => \N__5026\
        );

    \I__612\ : InMux
    port map (
            O => \N__5033\,
            I => \N__5023\
        );

    \I__611\ : InMux
    port map (
            O => \N__5032\,
            I => \N__5020\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__5029\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__609\ : Odrv4
    port map (
            O => \N__5026\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__5023\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__5020\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__606\ : InMux
    port map (
            O => \N__5011\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__605\ : InMux
    port map (
            O => \N__5008\,
            I => \N__5003\
        );

    \I__604\ : CascadeMux
    port map (
            O => \N__5007\,
            I => \N__5000\
        );

    \I__603\ : InMux
    port map (
            O => \N__5006\,
            I => \N__4997\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__5003\,
            I => \N__4994\
        );

    \I__601\ : InMux
    port map (
            O => \N__5000\,
            I => \N__4991\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__4997\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__599\ : Odrv4
    port map (
            O => \N__4994\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__4991\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__597\ : InMux
    port map (
            O => \N__4984\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__596\ : CascadeMux
    port map (
            O => \N__4981\,
            I => \N__4978\
        );

    \I__595\ : InMux
    port map (
            O => \N__4978\,
            I => \N__4975\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__4975\,
            I => \N__4969\
        );

    \I__593\ : InMux
    port map (
            O => \N__4974\,
            I => \N__4966\
        );

    \I__592\ : InMux
    port map (
            O => \N__4973\,
            I => \N__4962\
        );

    \I__591\ : InMux
    port map (
            O => \N__4972\,
            I => \N__4959\
        );

    \I__590\ : Sp12to4
    port map (
            O => \N__4969\,
            I => \N__4954\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__4966\,
            I => \N__4954\
        );

    \I__588\ : InMux
    port map (
            O => \N__4965\,
            I => \N__4951\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__4962\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__4959\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__585\ : Odrv12
    port map (
            O => \N__4954\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__4951\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__583\ : InMux
    port map (
            O => \N__4942\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__582\ : InMux
    port map (
            O => \N__4939\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__581\ : InMux
    port map (
            O => \N__4936\,
            I => \N__4932\
        );

    \I__580\ : InMux
    port map (
            O => \N__4935\,
            I => \N__4929\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__4932\,
            I => \N__4925\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__4929\,
            I => \N__4922\
        );

    \I__577\ : InMux
    port map (
            O => \N__4928\,
            I => \N__4919\
        );

    \I__576\ : Odrv4
    port map (
            O => \N__4925\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__575\ : Odrv4
    port map (
            O => \N__4922\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__4919\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__573\ : InMux
    port map (
            O => \N__4912\,
            I => \N__4909\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__4909\,
            I => \N__4906\
        );

    \I__571\ : Odrv4
    port map (
            O => \N__4906\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_1\
        );

    \I__570\ : CascadeMux
    port map (
            O => \N__4903\,
            I => \U712_CHIP_RAM.N_305_cascade_\
        );

    \I__569\ : CascadeMux
    port map (
            O => \N__4900\,
            I => \N__4896\
        );

    \I__568\ : CascadeMux
    port map (
            O => \N__4899\,
            I => \N__4893\
        );

    \I__567\ : InMux
    port map (
            O => \N__4896\,
            I => \N__4887\
        );

    \I__566\ : InMux
    port map (
            O => \N__4893\,
            I => \N__4887\
        );

    \I__565\ : InMux
    port map (
            O => \N__4892\,
            I => \N__4884\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__4887\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__4884\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__562\ : CascadeMux
    port map (
            O => \N__4879\,
            I => \N__4876\
        );

    \I__561\ : InMux
    port map (
            O => \N__4876\,
            I => \N__4873\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__4873\,
            I => \N__4868\
        );

    \I__559\ : InMux
    port map (
            O => \N__4872\,
            I => \N__4865\
        );

    \I__558\ : InMux
    port map (
            O => \N__4871\,
            I => \N__4862\
        );

    \I__557\ : Odrv4
    port map (
            O => \N__4868\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__4865\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__4862\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__554\ : InMux
    port map (
            O => \N__4855\,
            I => \N__4850\
        );

    \I__553\ : InMux
    port map (
            O => \N__4854\,
            I => \N__4847\
        );

    \I__552\ : InMux
    port map (
            O => \N__4853\,
            I => \N__4844\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__4850\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__4847\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__4844\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\
        );

    \I__548\ : InMux
    port map (
            O => \N__4837\,
            I => \N__4834\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4834\,
            I => \U712_CHIP_RAM.N_325\
        );

    \I__546\ : CascadeMux
    port map (
            O => \N__4831\,
            I => \U712_CHIP_RAM.N_325_cascade_\
        );

    \I__545\ : CascadeMux
    port map (
            O => \N__4828\,
            I => \U712_CHIP_RAM.m101_i_0_cascade_\
        );

    \I__544\ : InMux
    port map (
            O => \N__4825\,
            I => \N__4822\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__4822\,
            I => \U712_CHIP_RAM.m101_i_1\
        );

    \I__542\ : InMux
    port map (
            O => \N__4819\,
            I => \N__4816\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__4816\,
            I => \U712_CHIP_RAM.N_376\
        );

    \I__540\ : CascadeMux
    port map (
            O => \N__4813\,
            I => \U712_CHIP_RAM.m101_i_2_cascade_\
        );

    \I__539\ : InMux
    port map (
            O => \N__4810\,
            I => \N__4807\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__4807\,
            I => \U712_CHIP_RAM.N_436\
        );

    \I__537\ : CascadeMux
    port map (
            O => \N__4804\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_5_cascade_\
        );

    \I__536\ : CascadeMux
    port map (
            O => \N__4801\,
            I => \N__4798\
        );

    \I__535\ : InMux
    port map (
            O => \N__4798\,
            I => \N__4789\
        );

    \I__534\ : InMux
    port map (
            O => \N__4797\,
            I => \N__4789\
        );

    \I__533\ : InMux
    port map (
            O => \N__4796\,
            I => \N__4789\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__4789\,
            I => \U712_CHIP_RAM.SDRAM_CMDs_0_4\
        );

    \I__531\ : CascadeMux
    port map (
            O => \N__4786\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_1_1_cascade_\
        );

    \I__530\ : CascadeMux
    port map (
            O => \N__4783\,
            I => \U712_CHIP_RAM.N_396_cascade_\
        );

    \I__529\ : InMux
    port map (
            O => \N__4780\,
            I => \N__4777\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__4777\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_0_2\
        );

    \I__527\ : InMux
    port map (
            O => \N__4774\,
            I => \N__4771\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__4771\,
            I => \U712_CHIP_RAM.N_397\
        );

    \I__525\ : InMux
    port map (
            O => \N__4768\,
            I => \N__4765\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__4765\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_1_3\
        );

    \I__523\ : InMux
    port map (
            O => \N__4762\,
            I => \N__4756\
        );

    \I__522\ : InMux
    port map (
            O => \N__4761\,
            I => \N__4756\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__4756\,
            I => \N__4753\
        );

    \I__520\ : Odrv4
    port map (
            O => \N__4753\,
            I => \U712_CHIP_RAM.SDRAM_CMDs_0_1\
        );

    \I__519\ : CEMux
    port map (
            O => \N__4750\,
            I => \N__4747\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__4747\,
            I => \N__4744\
        );

    \I__517\ : Span4Mux_v
    port map (
            O => \N__4744\,
            I => \N__4741\
        );

    \I__516\ : Span4Mux_h
    port map (
            O => \N__4741\,
            I => \N__4738\
        );

    \I__515\ : Odrv4
    port map (
            O => \N__4738\,
            I => \U712_CHIP_RAM.N_194_0\
        );

    \I__514\ : InMux
    port map (
            O => \N__4735\,
            I => \N__4729\
        );

    \I__513\ : InMux
    port map (
            O => \N__4734\,
            I => \N__4729\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__4729\,
            I => \N__4726\
        );

    \I__511\ : Odrv4
    port map (
            O => \N__4726\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_3\
        );

    \I__510\ : CEMux
    port map (
            O => \N__4723\,
            I => \N__4720\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__4720\,
            I => \N__4717\
        );

    \I__508\ : Odrv4
    port map (
            O => \N__4717\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_0\
        );

    \I__507\ : InMux
    port map (
            O => \N__4714\,
            I => \N__4710\
        );

    \I__506\ : InMux
    port map (
            O => \N__4713\,
            I => \N__4707\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4710\,
            I => \N__4704\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__4707\,
            I => \N__4701\
        );

    \I__503\ : Span4Mux_v
    port map (
            O => \N__4704\,
            I => \N__4698\
        );

    \I__502\ : Span4Mux_v
    port map (
            O => \N__4701\,
            I => \N__4695\
        );

    \I__501\ : Sp12to4
    port map (
            O => \N__4698\,
            I => \N__4692\
        );

    \I__500\ : Span4Mux_h
    port map (
            O => \N__4695\,
            I => \N__4689\
        );

    \I__499\ : Span12Mux_h
    port map (
            O => \N__4692\,
            I => \N__4684\
        );

    \I__498\ : Sp12to4
    port map (
            O => \N__4689\,
            I => \N__4684\
        );

    \I__497\ : Span12Mux_v
    port map (
            O => \N__4684\,
            I => \N__4681\
        );

    \I__496\ : Odrv12
    port map (
            O => \N__4681\,
            I => \DBRn_c\
        );

    \I__495\ : InMux
    port map (
            O => \N__4678\,
            I => \N__4675\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__4675\,
            I => \N__4671\
        );

    \I__493\ : InMux
    port map (
            O => \N__4674\,
            I => \N__4668\
        );

    \I__492\ : Span4Mux_v
    port map (
            O => \N__4671\,
            I => \N__4663\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__4668\,
            I => \N__4663\
        );

    \I__490\ : Span4Mux_v
    port map (
            O => \N__4663\,
            I => \N__4660\
        );

    \I__489\ : Span4Mux_v
    port map (
            O => \N__4660\,
            I => \N__4657\
        );

    \I__488\ : Span4Mux_h
    port map (
            O => \N__4657\,
            I => \N__4654\
        );

    \I__487\ : Odrv4
    port map (
            O => \N__4654\,
            I => \TSn_c\
        );

    \I__486\ : InMux
    port map (
            O => \N__4651\,
            I => \N__4648\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__4648\,
            I => \N__4645\
        );

    \I__484\ : Span12Mux_v
    port map (
            O => \N__4645\,
            I => \N__4642\
        );

    \I__483\ : Odrv12
    port map (
            O => \N__4642\,
            I => \RAMSPACEn_c\
        );

    \I__482\ : InMux
    port map (
            O => \N__4639\,
            I => \N__4636\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__4636\,
            I => \N__4633\
        );

    \I__480\ : Span12Mux_v
    port map (
            O => \N__4633\,
            I => \N__4630\
        );

    \I__479\ : Odrv12
    port map (
            O => \N__4630\,
            I => \U712_CHIP_RAM.N_419\
        );

    \I__478\ : IoInMux
    port map (
            O => \N__4627\,
            I => \N__4624\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__4624\,
            I => \N__4621\
        );

    \I__476\ : Odrv12
    port map (
            O => \N__4621\,
            I => \VBENn_c\
        );

    \I__475\ : InMux
    port map (
            O => \N__4618\,
            I => \N__4615\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__4615\,
            I => \U712_CHIP_RAM.N_428\
        );

    \I__473\ : CascadeMux
    port map (
            O => \N__4612\,
            I => \U712_CHIP_RAM.N_307_cascade_\
        );

    \I__472\ : CascadeMux
    port map (
            O => \N__4609\,
            I => \U712_CHIP_RAM.N_467_cascade_\
        );

    \I__471\ : CascadeMux
    port map (
            O => \N__4606\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_\
        );

    \I__470\ : InMux
    port map (
            O => \N__4603\,
            I => \N__4599\
        );

    \I__469\ : InMux
    port map (
            O => \N__4602\,
            I => \N__4596\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__4599\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__4596\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__466\ : InMux
    port map (
            O => \N__4591\,
            I => \N__4587\
        );

    \I__465\ : InMux
    port map (
            O => \N__4590\,
            I => \N__4584\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__4587\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__4584\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__462\ : InMux
    port map (
            O => \N__4579\,
            I => \N__4575\
        );

    \I__461\ : InMux
    port map (
            O => \N__4578\,
            I => \N__4572\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__4575\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__4572\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__458\ : CascadeMux
    port map (
            O => \N__4567\,
            I => \U712_CHIP_RAM.REFRESH5lto7_0_cascade_\
        );

    \I__457\ : InMux
    port map (
            O => \N__4564\,
            I => \N__4560\
        );

    \I__456\ : InMux
    port map (
            O => \N__4563\,
            I => \N__4557\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__4560\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__4557\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__453\ : InMux
    port map (
            O => \N__4552\,
            I => \N__4548\
        );

    \I__452\ : InMux
    port map (
            O => \N__4551\,
            I => \N__4545\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__4548\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__4545\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__449\ : CascadeMux
    port map (
            O => \N__4540\,
            I => \N__4536\
        );

    \I__448\ : InMux
    port map (
            O => \N__4539\,
            I => \N__4533\
        );

    \I__447\ : InMux
    port map (
            O => \N__4536\,
            I => \N__4530\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__4533\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__4530\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__444\ : InMux
    port map (
            O => \N__4525\,
            I => \N__4521\
        );

    \I__443\ : InMux
    port map (
            O => \N__4524\,
            I => \N__4518\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__4521\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__4518\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__440\ : InMux
    port map (
            O => \N__4513\,
            I => \N__4510\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__4510\,
            I => \U712_CHIP_RAM.REFRESH5lt7\
        );

    \I__438\ : CascadeMux
    port map (
            O => \N__4507\,
            I => \U712_CHIP_RAM.N_430_cascade_\
        );

    \I__437\ : InMux
    port map (
            O => \N__4504\,
            I => \N__4501\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__4501\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\
        );

    \I__435\ : InMux
    port map (
            O => \N__4498\,
            I => \N__4495\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__4495\,
            I => \N__4492\
        );

    \I__433\ : Span4Mux_h
    port map (
            O => \N__4492\,
            I => \N__4489\
        );

    \I__432\ : Sp12to4
    port map (
            O => \N__4489\,
            I => \N__4486\
        );

    \I__431\ : Span12Mux_v
    port map (
            O => \N__4486\,
            I => \N__4483\
        );

    \I__430\ : Odrv12
    port map (
            O => \N__4483\,
            I => \A_c_2\
        );

    \I__429\ : InMux
    port map (
            O => \N__4480\,
            I => \N__4477\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__4477\,
            I => \N__4474\
        );

    \I__427\ : Span12Mux_v
    port map (
            O => \N__4474\,
            I => \N__4471\
        );

    \I__426\ : Odrv12
    port map (
            O => \N__4471\,
            I => \A_c_4\
        );

    \I__425\ : InMux
    port map (
            O => \N__4468\,
            I => \N__4465\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__4465\,
            I => \N__4462\
        );

    \I__423\ : Span4Mux_v
    port map (
            O => \N__4462\,
            I => \N__4459\
        );

    \I__422\ : Span4Mux_v
    port map (
            O => \N__4459\,
            I => \N__4456\
        );

    \I__421\ : Sp12to4
    port map (
            O => \N__4456\,
            I => \N__4453\
        );

    \I__420\ : Odrv12
    port map (
            O => \N__4453\,
            I => \A_c_7\
        );

    \I__419\ : InMux
    port map (
            O => \N__4450\,
            I => \N__4447\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__4447\,
            I => \N__4444\
        );

    \I__417\ : Span12Mux_v
    port map (
            O => \N__4444\,
            I => \N__4441\
        );

    \I__416\ : Odrv12
    port map (
            O => \N__4441\,
            I => \A_c_8\
        );

    \I__415\ : InMux
    port map (
            O => \N__4438\,
            I => \N__4435\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__4435\,
            I => \N__4432\
        );

    \I__413\ : Span12Mux_h
    port map (
            O => \N__4432\,
            I => \N__4429\
        );

    \I__412\ : Span12Mux_v
    port map (
            O => \N__4429\,
            I => \N__4426\
        );

    \I__411\ : Odrv12
    port map (
            O => \N__4426\,
            I => \REGSPACEn_c\
        );

    \I__410\ : CascadeMux
    port map (
            O => \N__4423\,
            I => \U712_CHIP_RAM.m93_i_a2_4_cascade_\
        );

    \I__409\ : IoInMux
    port map (
            O => \N__4420\,
            I => \N__4417\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__4417\,
            I => \N__4414\
        );

    \I__407\ : Span4Mux_s2_v
    port map (
            O => \N__4414\,
            I => \N__4411\
        );

    \I__406\ : Span4Mux_v
    port map (
            O => \N__4411\,
            I => \N__4408\
        );

    \I__405\ : Span4Mux_h
    port map (
            O => \N__4408\,
            I => \N__4405\
        );

    \I__404\ : Odrv4
    port map (
            O => \N__4405\,
            I => \CLK80_PLL_i_i\
        );

    \I__403\ : InMux
    port map (
            O => \N__4402\,
            I => \N__4399\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__4399\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__401\ : InMux
    port map (
            O => \N__4396\,
            I => \bfn_6_6_0_\
        );

    \I__400\ : InMux
    port map (
            O => \N__4393\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__399\ : InMux
    port map (
            O => \N__4390\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__398\ : InMux
    port map (
            O => \N__4387\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__397\ : InMux
    port map (
            O => \N__4384\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__396\ : InMux
    port map (
            O => \N__4381\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__395\ : InMux
    port map (
            O => \N__4378\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__394\ : InMux
    port map (
            O => \N__4375\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__393\ : ClkMux
    port map (
            O => \N__4372\,
            I => \N__4348\
        );

    \I__392\ : ClkMux
    port map (
            O => \N__4371\,
            I => \N__4348\
        );

    \I__391\ : ClkMux
    port map (
            O => \N__4370\,
            I => \N__4348\
        );

    \I__390\ : ClkMux
    port map (
            O => \N__4369\,
            I => \N__4348\
        );

    \I__389\ : ClkMux
    port map (
            O => \N__4368\,
            I => \N__4348\
        );

    \I__388\ : ClkMux
    port map (
            O => \N__4367\,
            I => \N__4348\
        );

    \I__387\ : ClkMux
    port map (
            O => \N__4366\,
            I => \N__4348\
        );

    \I__386\ : ClkMux
    port map (
            O => \N__4365\,
            I => \N__4348\
        );

    \I__385\ : GlobalMux
    port map (
            O => \N__4348\,
            I => \N__4345\
        );

    \I__384\ : gio2CtrlBuf
    port map (
            O => \N__4345\,
            I => \C1_c_g\
        );

    \I__383\ : IoInMux
    port map (
            O => \N__4342\,
            I => \N__4339\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__4339\,
            I => \N__4336\
        );

    \I__381\ : Span12Mux_s4_h
    port map (
            O => \N__4336\,
            I => \N__4333\
        );

    \I__380\ : Odrv12
    port map (
            O => \N__4333\,
            I => \DBRn_c_i_0\
        );

    \I__379\ : IoInMux
    port map (
            O => \N__4330\,
            I => \N__4327\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__4327\,
            I => \N__4324\
        );

    \I__377\ : Span4Mux_s0_v
    port map (
            O => \N__4324\,
            I => \N__4321\
        );

    \I__376\ : Span4Mux_v
    port map (
            O => \N__4321\,
            I => \N__4318\
        );

    \I__375\ : Sp12to4
    port map (
            O => \N__4318\,
            I => \N__4315\
        );

    \I__374\ : Span12Mux_h
    port map (
            O => \N__4315\,
            I => \N__4312\
        );

    \I__373\ : Span12Mux_v
    port map (
            O => \N__4312\,
            I => \N__4309\
        );

    \I__372\ : Odrv12
    port map (
            O => \N__4309\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            I => \N__4371\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__4365\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            I => \N__4366\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            I => \N__4369\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__4368\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\,
            I => \N__4367\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            I => \N__4370\
        );

    \IN_MUX_bfv_10_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_5_0_\
        );

    \IN_MUX_bfv_6_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_6_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_8_0_\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5889\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__9592\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4342\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6031\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__8220\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10567\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9973\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4402\,
            in2 => \_gnd_net_\,
            in3 => \N__4396\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_6_6_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__4372\,
            ce => 'H',
            sr => \N__6190\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4525\,
            in2 => \_gnd_net_\,
            in3 => \N__4393\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__4372\,
            ce => 'H',
            sr => \N__6190\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4552\,
            in2 => \_gnd_net_\,
            in3 => \N__4390\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__4372\,
            ce => 'H',
            sr => \N__6190\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4564\,
            in2 => \_gnd_net_\,
            in3 => \N__4387\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__4372\,
            ce => 'H',
            sr => \N__6190\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4539\,
            in2 => \_gnd_net_\,
            in3 => \N__4384\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__4372\,
            ce => 'H',
            sr => \N__6190\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4591\,
            in2 => \_gnd_net_\,
            in3 => \N__4381\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__4372\,
            ce => 'H',
            sr => \N__6190\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4603\,
            in2 => \_gnd_net_\,
            in3 => \N__4378\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__4372\,
            ce => 'H',
            sr => \N__6190\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4578\,
            in2 => \_gnd_net_\,
            in3 => \N__4375\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4372\,
            ce => 'H',
            sr => \N__6190\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4498\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9948\,
            ce => \N__6407\,
            sr => \N__10539\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4480\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9948\,
            ce => \N__6407\,
            sr => \N__10539\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4468\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9948\,
            ce => \N__6407\,
            sr => \N__10539\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4450\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9948\,
            ce => \N__6407\,
            sr => \N__10539\
        );

    \DBRn_ibuf_RNIBAB_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4713\,
            lcout => \DBRn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__4438\,
            in1 => \N__4678\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.N_402\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__6885\,
            in1 => \N__7194\,
            in2 => \N__7344\,
            in3 => \N__7033\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDs_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4855\,
            in1 => \N__6352\,
            in2 => \_gnd_net_\,
            in3 => \N__6373\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m93_i_a2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6331\,
            in1 => \N__6199\,
            in2 => \N__4423\,
            in3 => \N__5944\,
            lcout => \U712_CHIP_RAM.N_428\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4602\,
            in2 => \_gnd_net_\,
            in3 => \N__4590\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.REFRESH5lto7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001010"
        )
    port map (
            in0 => \N__10207\,
            in1 => \N__4579\,
            in2 => \N__4567\,
            in3 => \N__4513\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9943\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__4563\,
            in1 => \N__4551\,
            in2 => \N__4540\,
            in3 => \N__4524\,
            lcout => \U712_CHIP_RAM.REFRESH5lt7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6ORT_7_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4935\,
            in2 => \_gnd_net_\,
            in3 => \N__5008\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDs_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIJNSTA_0_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10566\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5513\,
            lcout => \U712_CHIP_RAM.N_194_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6657\,
            in1 => \N__4734\,
            in2 => \_gnd_net_\,
            in3 => \N__4504\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_430_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__5707\,
            in1 => \N__10199\,
            in2 => \N__4507\,
            in3 => \N__5772\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9945\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011001000"
        )
    port map (
            in0 => \N__4639\,
            in1 => \N__10193\,
            in2 => \N__4900\,
            in3 => \N__11675\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9945\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_4_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4735\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10200\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9945\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__4872\,
            in1 => \N__4854\,
            in2 => \N__4899\,
            in3 => \N__5706\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6658\,
            in1 => \N__7645\,
            in2 => \N__10206\,
            in3 => \N__4618\,
            lcout => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9945\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI3M1M2_1_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__7159\,
            in1 => \N__6856\,
            in2 => \_gnd_net_\,
            in3 => \N__7221\,
            lcout => \U712_CHIP_RAM.m101_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__4837\,
            in1 => \N__10202\,
            in2 => \N__5727\,
            in3 => \N__5484\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4965\,
            in1 => \N__5032\,
            in2 => \N__5007\,
            in3 => \N__4928\,
            lcout => \U712_CHIP_RAM.N_307\,
            ltout => \U712_CHIP_RAM.N_307_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6777\,
            in1 => \N__6859\,
            in2 => \N__4612\,
            in3 => \N__7307\,
            lcout => \U712_CHIP_RAM.N_467\,
            ltout => \U712_CHIP_RAM.N_467_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7023\,
            in2 => \N__4609\,
            in3 => \N__7129\,
            lcout => \U712_CHIP_RAM.N_476\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU7TF5_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7024\,
            in1 => \N__5463\,
            in2 => \N__7170\,
            in3 => \N__5421\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKHPV5_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10565\,
            in1 => \_gnd_net_\,
            in2 => \N__4606\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__7025\,
            in1 => \_gnd_net_\,
            in2 => \N__7171\,
            in3 => \N__5422\,
            lcout => \U712_CHIP_RAM.N_440\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5423\,
            in1 => \N__7026\,
            in2 => \N__7195\,
            in3 => \N__5714\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9949\,
            ce => \N__4723\,
            sr => \N__10529\
        );

    \U712_CHIP_RAM.RAS_SYNC_3_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10201\,
            in2 => \_gnd_net_\,
            in3 => \N__9982\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9954\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10564\,
            in2 => \_gnd_net_\,
            in3 => \N__5088\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBR_SYNC_0_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4714\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9959\,
            ce => 'H',
            sr => \N__10515\
        );

    \U712_REG_SM.WRITE_CYCLE_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__10380\,
            in1 => \N__7455\,
            in2 => \_gnd_net_\,
            in3 => \N__8522\,
            lcout => \U712_REG_SM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9968\,
            ce => 'H',
            sr => \N__10500\
        );

    \U712_REG_SM.LDSn_RNO_0_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__11208\,
            in1 => \N__11332\,
            in2 => \N__11100\,
            in3 => \N__10384\,
            lcout => \U712_REG_SM.N_404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4674\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4651\,
            lcout => \U712_CHIP_RAM.N_419\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_0_a2_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__11676\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7441\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__6172\,
            in1 => \N__7187\,
            in2 => \N__4801\,
            in3 => \N__4912\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMDsr_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101111001000"
        )
    port map (
            in0 => \N__6691\,
            in1 => \N__5518\,
            in2 => \N__4804\,
            in3 => \N__8138\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9936\,
            ce => 'H',
            sr => \N__10540\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_1_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4796\,
            in1 => \N__5041\,
            in2 => \N__4981\,
            in3 => \N__5137\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_2_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011110"
        )
    port map (
            in0 => \N__7032\,
            in1 => \N__4974\,
            in2 => \N__6793\,
            in3 => \N__5040\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMDsr_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_2_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__7335\,
            in1 => \N__4797\,
            in2 => \N__4786\,
            in3 => \N__6791\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_1_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100000000"
        )
    port map (
            in0 => \N__6886\,
            in1 => \N__7031\,
            in2 => \N__4879\,
            in3 => \N__7186\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_396_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_1_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4774\,
            in1 => \N__4761\,
            in2 => \N__4783\,
            in3 => \N__4780\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9939\,
            ce => \N__4750\,
            sr => \N__10535\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_1_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001000"
        )
    port map (
            in0 => \N__7336\,
            in1 => \N__7185\,
            in2 => \N__5731\,
            in3 => \N__7030\,
            lcout => \U712_CHIP_RAM.N_397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_2_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4768\,
            in1 => \N__5494\,
            in2 => \N__5269\,
            in3 => \N__4762\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9939\,
            ce => \N__4750\,
            sr => \N__10535\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__6784\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7833\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__7304\,
            in1 => \N__4972\,
            in2 => \_gnd_net_\,
            in3 => \N__5033\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6855\,
            in2 => \_gnd_net_\,
            in3 => \N__6752\,
            lcout => \U712_CHIP_RAM.N_305\,
            ltout => \U712_CHIP_RAM.N_305_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNI7MCB2_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110100001"
        )
    port map (
            in0 => \N__7302\,
            in1 => \N__5702\,
            in2 => \N__4903\,
            in3 => \N__6977\,
            lcout => \U712_CHIP_RAM.N_376\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__4892\,
            in1 => \N__4871\,
            in2 => \_gnd_net_\,
            in3 => \N__4853\,
            lcout => \U712_CHIP_RAM.N_325\,
            ltout => \U712_CHIP_RAM.N_325_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNICN5A2_2_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6978\,
            in2 => \N__4831\,
            in3 => \N__6602\,
            lcout => \U712_CHIP_RAM.N_436\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIGB4P1_3_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010101010101"
        )
    port map (
            in0 => \N__10198\,
            in1 => \N__7160\,
            in2 => \N__7021\,
            in3 => \N__7303\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m101_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI7AC23_0_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110101"
        )
    port map (
            in0 => \N__7161\,
            in1 => \N__6758\,
            in2 => \N__4828\,
            in3 => \N__6982\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m101_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITD0EA_0_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__4825\,
            in1 => \N__4819\,
            in2 => \N__4813\,
            in3 => \N__4810\,
            lcout => \U712_CHIP_RAM.N_194\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6773\,
            in2 => \_gnd_net_\,
            in3 => \N__5771\,
            lcout => \U712_CHIP_RAM.LATCH_CLK_6\,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5393\,
            in1 => \N__6873\,
            in2 => \_gnd_net_\,
            in3 => \N__5050\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__9946\,
            ce => \N__5331\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7018\,
            in2 => \_gnd_net_\,
            in3 => \N__5047\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5394\,
            in1 => \N__7325\,
            in2 => \_gnd_net_\,
            in3 => \N__5044\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__9946\,
            ce => \N__5331\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5382\,
            in1 => \N__5039\,
            in2 => \_gnd_net_\,
            in3 => \N__5011\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__9946\,
            ce => \N__5331\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5395\,
            in1 => \N__5006\,
            in2 => \_gnd_net_\,
            in3 => \N__4984\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__9946\,
            ce => \N__5331\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5383\,
            in1 => \N__4973\,
            in2 => \_gnd_net_\,
            in3 => \N__4942\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__9946\,
            ce => \N__5331\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__4936\,
            in1 => \N__5384\,
            in2 => \_gnd_net_\,
            in3 => \N__4939\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9946\,
            ce => \N__5331\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__7126\,
            in1 => \N__7306\,
            in2 => \N__6792\,
            in3 => \N__6986\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_0_a3_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6764\,
            in1 => \N__5652\,
            in2 => \N__7022\,
            in3 => \N__7127\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__7128\,
            in1 => \_gnd_net_\,
            in2 => \N__5140\,
            in3 => \N__10172\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9950\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_3_1_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011010011"
        )
    port map (
            in0 => \N__6985\,
            in1 => \N__6858\,
            in2 => \N__6778\,
            in3 => \N__7125\,
            lcout => \U712_CHIP_RAM.N_378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__7124\,
            in1 => \N__6984\,
            in2 => \N__5732\,
            in3 => \N__5420\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI41RO8_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5128\,
            in3 => \N__5838\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI8UIP2_3_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__6857\,
            in1 => \N__7305\,
            in2 => \_gnd_net_\,
            in3 => \N__7222\,
            lcout => \U712_CHIP_RAM.N_551\,
            ltout => \U712_CHIP_RAM.N_551_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOBA64_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6983\,
            in1 => \N__7123\,
            in2 => \N__5125\,
            in3 => \N__6167\,
            lcout => \U712_CHIP_RAM.N_435\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111011100000010"
        )
    port map (
            in0 => \N__5122\,
            in1 => \N__7357\,
            in2 => \N__7246\,
            in3 => \N__5100\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9955\,
            ce => 'H',
            sr => \N__10509\
        );

    \U712_CHIP_RAM.DBENn_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101111111001100"
        )
    port map (
            in0 => \N__5434\,
            in1 => \N__5800\,
            in2 => \N__5746\,
            in3 => \N__5089\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9955\,
            ce => 'H',
            sr => \N__10509\
        );

    \U712_CHIP_RAM.DBDIR_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__5589\,
            in1 => \N__5061\,
            in2 => \_gnd_net_\,
            in3 => \N__5562\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9955\,
            ce => 'H',
            sr => \N__10509\
        );

    \U712_REG_SM.REGENn_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011010010110000"
        )
    port map (
            in0 => \N__7958\,
            in1 => \N__5167\,
            in2 => \N__5214\,
            in3 => \N__5239\,
            lcout => \REGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9960\,
            ce => 'H',
            sr => \N__10504\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001101"
        )
    port map (
            in0 => \N__5755\,
            in1 => \N__5254\,
            in2 => \N__7680\,
            in3 => \N__8035\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9963\,
            ce => 'H',
            sr => \N__10501\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7570\,
            in1 => \N__8038\,
            in2 => \N__7681\,
            in3 => \N__5183\,
            lcout => \U712_REG_SM.N_412\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010101000"
        )
    port map (
            in0 => \N__10166\,
            in1 => \N__5248\,
            in2 => \N__5188\,
            in3 => \N__8467\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9965\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5182\,
            in1 => \N__5238\,
            in2 => \N__7535\,
            in3 => \N__7940\,
            lcout => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_RNO_0_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100001011000"
        )
    port map (
            in0 => \N__5213\,
            in1 => \N__8495\,
            in2 => \N__7537\,
            in3 => \N__5187\,
            lcout => \U712_REG_SM.REGENn_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDSn_RNO_0_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__11342\,
            in1 => \N__11087\,
            in2 => \N__11263\,
            in3 => \N__10385\,
            lcout => \U712_REG_SM.N_459\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBR_COUNT_1_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__5939\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6231\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9934\,
            ce => 'H',
            sr => \N__6676\
        );

    \U712_CHIP_RAM.DBR_COUNT_0_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5938\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9934\,
            ce => 'H',
            sr => \N__6676\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5158\,
            in1 => \N__5275\,
            in2 => \_gnd_net_\,
            in3 => \N__8857\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8858\,
            in1 => \N__5314\,
            in2 => \_gnd_net_\,
            in3 => \N__5533\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__11610\,
            in1 => \N__8859\,
            in2 => \N__5296\,
            in3 => \N__8203\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5293\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9937\,
            ce => \N__6409\,
            sr => \N__10530\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__8131\,
            in1 => \N__8888\,
            in2 => \_gnd_net_\,
            in3 => \N__8159\,
            lcout => \U712_CHIP_RAM.CMA_5_i_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIUI4B1_0_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8158\,
            in1 => \N__8130\,
            in2 => \N__9572\,
            in3 => \N__8856\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_3_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110100001010"
        )
    port map (
            in0 => \N__6760\,
            in1 => \N__7308\,
            in2 => \N__7188\,
            in3 => \N__7002\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIMT791_1_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7162\,
            in1 => \N__6863\,
            in2 => \_gnd_net_\,
            in3 => \N__6759\,
            lcout => \U712_CHIP_RAM.N_555\,
            ltout => \U712_CHIP_RAM.N_555_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6603\,
            in2 => \N__5257\,
            in3 => \N__7309\,
            lcout => \U712_CHIP_RAM.N_390\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__7004\,
            in1 => \N__7167\,
            in2 => \_gnd_net_\,
            in3 => \N__6865\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMDsr_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101111001000"
        )
    port map (
            in0 => \N__6538\,
            in1 => \N__5514\,
            in2 => \N__5497\,
            in3 => \N__9566\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9940\,
            ce => 'H',
            sr => \N__10522\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_2_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__7003\,
            in1 => \N__7166\,
            in2 => \_gnd_net_\,
            in3 => \N__6864\,
            lcout => \U712_CHIP_RAM.N_449\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIB0JV5_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__5488\,
            in1 => \N__5470\,
            in2 => \_gnd_net_\,
            in3 => \N__5733\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__10173\,
            in1 => \N__5452\,
            in2 => \N__5446\,
            in3 => \N__5385\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9944\,
            ce => \N__5335\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7384\,
            in2 => \_gnd_net_\,
            in3 => \N__6753\,
            lcout => \U712_CHIP_RAM.N_304\,
            ltout => \U712_CHIP_RAM.N_304_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNID3LR1_0_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010001000"
        )
    port map (
            in0 => \N__6754\,
            in1 => \N__6999\,
            in2 => \N__5443\,
            in3 => \N__7168\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_312_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIBB455_0_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10174\,
            in2 => \N__5440\,
            in3 => \N__5651\,
            lcout => \U712_CHIP_RAM.N_326\,
            ltout => \U712_CHIP_RAM.N_326_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIA8V79_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111110000"
        )
    port map (
            in0 => \N__7169\,
            in1 => \N__7000\,
            in2 => \N__5437\,
            in3 => \N__5430\,
            lcout => \U712_CHIP_RAM.N_39\,
            ltout => \U712_CHIP_RAM.N_39_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000111010"
        )
    port map (
            in0 => \N__5362\,
            in1 => \N__5353\,
            in2 => \N__5344\,
            in3 => \N__5341\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9944\,
            ce => \N__5335\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7019\,
            in2 => \_gnd_net_\,
            in3 => \N__9754\,
            lcout => \U712_CHIP_RAM.DBENn_7_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__5737\,
            in1 => \N__10389\,
            in2 => \_gnd_net_\,
            in3 => \N__5596\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_344_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__10171\,
            in1 => \N__5662\,
            in2 => \N__5656\,
            in3 => \N__7386\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9947\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7020\,
            in1 => \N__7366\,
            in2 => \N__7190\,
            in3 => \N__5653\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER41_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__10170\,
            in1 => \N__5607\,
            in2 => \N__5635\,
            in3 => \N__5632\,
            lcout => \LATCH_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9947\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIDTSL_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__7385\,
            in1 => \N__6866\,
            in2 => \_gnd_net_\,
            in3 => \N__11568\,
            lcout => \U712_CHIP_RAM.N_20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011000000"
        )
    port map (
            in0 => \N__5595\,
            in1 => \N__11738\,
            in2 => \N__10197\,
            in3 => \N__5563\,
            lcout => \DMA_WRITE_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9947\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__5854\,
            in1 => \N__5551\,
            in2 => \N__10867\,
            in3 => \N__5532\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9951\,
            ce => 'H',
            sr => \N__10505\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__11606\,
            in1 => \N__5853\,
            in2 => \_gnd_net_\,
            in3 => \N__5839\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9951\,
            ce => 'H',
            sr => \N__10505\
        );

    \DBR_SYNC_1_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5827\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9951\,
            ce => 'H',
            sr => \N__10505\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5801\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5781\,
            lcout => \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__8030\,
            in1 => \N__7600\,
            in2 => \N__7543\,
            in3 => \N__7632\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_413_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000010"
        )
    port map (
            in0 => \N__10183\,
            in1 => \N__7542\,
            in2 => \N__5818\,
            in3 => \N__7959\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9956\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNIFFA4_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__5802\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5782\,
            lcout => \U712_CHIP_RAM.m50_i_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__7568\,
            in1 => \N__7536\,
            in2 => \_gnd_net_\,
            in3 => \N__7957\,
            lcout => \U712_REG_SM.N_308\,
            ltout => \U712_REG_SM.N_308_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__10163\,
            in1 => \N__8034\,
            in2 => \N__5749\,
            in3 => \N__7569\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9961\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__10160\,
            in1 => \N__9210\,
            in2 => \_gnd_net_\,
            in3 => \N__8611\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9961\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5908\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10161\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9961\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10162\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6141\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9961\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6140\,
            in2 => \_gnd_net_\,
            in3 => \N__5907\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__10165\,
            in1 => \N__5896\,
            in2 => \N__8524\,
            in3 => \N__8494\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9964\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNINRSB_2_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7594\,
            in2 => \_gnd_net_\,
            in3 => \N__8492\,
            lcout => \U712_REG_SM.N_328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_0_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7595\,
            in1 => \N__7641\,
            in2 => \N__7534\,
            in3 => \N__7936\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_410_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011100100"
        )
    port map (
            in0 => \N__10164\,
            in1 => \N__7422\,
            in2 => \N__5899\,
            in3 => \N__7462\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9964\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIVCF31_4_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011011111"
        )
    port map (
            in0 => \N__7566\,
            in1 => \N__7506\,
            in2 => \N__7956\,
            in3 => \N__8493\,
            lcout => \U712_REG_SM.un1_REGENn_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7533\,
            in3 => \N__7935\,
            lcout => \U712_REG_SM.N_331\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_0_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5890\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9966\,
            ce => 'H',
            sr => \N__10493\
        );

    \U712_REG_SM.C1_SYNC_1_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6151\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9966\,
            ce => 'H',
            sr => \N__10493\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110110011101110"
        )
    port map (
            in0 => \N__6082\,
            in1 => \N__6145\,
            in2 => \N__9211\,
            in3 => \N__8610\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9966\,
            ce => 'H',
            sr => \N__10493\
        );

    \U712_REG_SM.LDSn_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011101110111000"
        )
    port map (
            in0 => \N__6042\,
            in1 => \N__7989\,
            in2 => \N__7960\,
            in3 => \N__6067\,
            lcout => \LDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9966\,
            ce => 'H',
            sr => \N__10493\
        );

    \U712_REG_SM.C3_SYNC_0_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6018\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9966\,
            ce => 'H',
            sr => \N__10493\
        );

    \U712_REG_SM.C3_SYNC_1_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5989\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9966\,
            ce => 'H',
            sr => \N__10493\
        );

    \U712_REG_SM.UDSn_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111001111100010"
        )
    port map (
            in0 => \N__5983\,
            in1 => \N__7990\,
            in2 => \N__5961\,
            in3 => \N__7951\,
            lcout => \UDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9969\,
            ce => 'H',
            sr => \N__10488\
        );

    \U712_CHIP_RAM.un3_DBR_COUNT_cry_1_c_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6230\,
            in2 => \N__5940\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_5_0_\,
            carryout => \U712_CHIP_RAM.un3_DBR_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBR_COUNT_2_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6244\,
            in2 => \_gnd_net_\,
            in3 => \N__5914\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un3_DBR_COUNT_cry_1\,
            carryout => \U712_CHIP_RAM.un3_DBR_COUNT_cry_2\,
            clk => \N__9929\,
            ce => 'H',
            sr => \N__6675\
        );

    \U712_CHIP_RAM.DBR_COUNT_3_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6256\,
            in2 => \_gnd_net_\,
            in3 => \N__5911\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un3_DBR_COUNT_cry_2\,
            carryout => \U712_CHIP_RAM.un3_DBR_COUNT_cry_3\,
            clk => \N__9929\,
            ce => 'H',
            sr => \N__6675\
        );

    \U712_CHIP_RAM.DBR_COUNT_4_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6369\,
            in2 => \_gnd_net_\,
            in3 => \N__6355\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un3_DBR_COUNT_cry_3\,
            carryout => \U712_CHIP_RAM.un3_DBR_COUNT_cry_4\,
            clk => \N__9929\,
            ce => 'H',
            sr => \N__6675\
        );

    \U712_CHIP_RAM.DBR_COUNT_5_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6348\,
            in2 => \_gnd_net_\,
            in3 => \N__6334\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un3_DBR_COUNT_cry_4\,
            carryout => \U712_CHIP_RAM.un3_DBR_COUNT_cry_5\,
            clk => \N__9929\,
            ce => 'H',
            sr => \N__6675\
        );

    \U712_CHIP_RAM.DBR_COUNT_6_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6327\,
            in2 => \_gnd_net_\,
            in3 => \N__6313\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un3_DBR_COUNT_cry_5\,
            carryout => \U712_CHIP_RAM.un3_DBR_COUNT_cry_6\,
            clk => \N__9929\,
            ce => 'H',
            sr => \N__6675\
        );

    \U712_CHIP_RAM.DBR_COUNT_7_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6211\,
            in2 => \_gnd_net_\,
            in3 => \N__6310\,
            lcout => \U712_CHIP_RAM.DBR_COUNTZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9929\,
            ce => 'H',
            sr => \N__6675\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6307\,
            in1 => \N__6433\,
            in2 => \_gnd_net_\,
            in3 => \N__8890\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6276\,
            in1 => \N__6463\,
            in2 => \_gnd_net_\,
            in3 => \N__8891\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_2_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6255\,
            in1 => \N__6243\,
            in2 => \N__6232\,
            in3 => \N__6210\,
            lcout => \U712_CHIP_RAM.m93_i_a2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIB72G2_3_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__8889\,
            in1 => \N__9565\,
            in2 => \N__8177\,
            in3 => \N__6186\,
            lcout => \U712_CHIP_RAM.un1_CMA25_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011110100111"
        )
    port map (
            in0 => \N__7017\,
            in1 => \N__6891\,
            in2 => \N__7345\,
            in3 => \N__6168\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m123_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__7189\,
            in1 => \N__6607\,
            in2 => \N__6586\,
            in3 => \N__7244\,
            lcout => \U712_CHIP_RAM.N_190\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6583\,
            in1 => \N__6562\,
            in2 => \_gnd_net_\,
            in3 => \N__8960\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8961\,
            in1 => \N__11611\,
            in2 => \N__6553\,
            in3 => \N__9292\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__7243\,
            in1 => \N__6550\,
            in2 => \_gnd_net_\,
            in3 => \N__6544\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6522\,
            in1 => \N__6487\,
            in2 => \_gnd_net_\,
            in3 => \N__8959\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6478\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9941\,
            ce => \N__6408\,
            sr => \N__10510\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6454\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9941\,
            ce => \N__6408\,
            sr => \N__10510\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6424\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9941\,
            ce => \N__6408\,
            sr => \N__10510\
        );

    \U712_BUFFERS.N_167_i_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101010"
        )
    port map (
            in0 => \N__11573\,
            in1 => \N__11845\,
            in2 => \N__10318\,
            in3 => \N__7434\,
            lcout => \N_167_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_0_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7387\,
            in2 => \_gnd_net_\,
            in3 => \N__6772\,
            lcout => \U712_CHIP_RAM.N_321\,
            ltout => \U712_CHIP_RAM.N_321_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__11572\,
            in1 => \N__7016\,
            in2 => \N__7360\,
            in3 => \N__6890\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.m77_0_a2_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__7356\,
            in1 => \N__7340\,
            in2 => \N__7249\,
            in3 => \N__7245\,
            lcout => \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101101110"
        )
    port map (
            in0 => \N__7172\,
            in1 => \N__7001\,
            in2 => \N__6892\,
            in3 => \N__6771\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_RNIEU0T_1_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__10152\,
            in1 => \N__6645\,
            in2 => \_gnd_net_\,
            in3 => \N__7636\,
            lcout => \U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10056\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6613\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9952\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNIVU9S_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000111"
        )
    port map (
            in0 => \N__11580\,
            in1 => \N__7969\,
            in2 => \N__9255\,
            in3 => \N__10314\,
            lcout => \N_202_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__11835\,
            in1 => \N__10055\,
            in2 => \_gnd_net_\,
            in3 => \N__10313\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9952\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000111000001100"
        )
    port map (
            in0 => \N__7765\,
            in1 => \N__7759\,
            in2 => \N__8609\,
            in3 => \N__8530\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9957\,
            ce => 'H',
            sr => \N__10495\
        );

    \U712_CYCLE_TERM.TACK_EN_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011111111"
        )
    port map (
            in0 => \N__7758\,
            in1 => \N__7696\,
            in2 => \_gnd_net_\,
            in3 => \N__8185\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9957\,
            ce => 'H',
            sr => \N__10495\
        );

    \U712_REG_SM.REG_TACK_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__8575\,
            in1 => \N__7673\,
            in2 => \N__7654\,
            in3 => \N__7996\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9957\,
            ce => 'H',
            sr => \N__10495\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__7942\,
            in1 => \N__8037\,
            in2 => \_gnd_net_\,
            in3 => \N__7526\,
            lcout => \U712_REG_SM.N_406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7527\,
            in2 => \_gnd_net_\,
            in3 => \N__7640\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_330_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000100010"
        )
    port map (
            in0 => \N__10159\,
            in1 => \N__7576\,
            in2 => \N__7603\,
            in3 => \N__7944\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9962\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111011"
        )
    port map (
            in0 => \N__7943\,
            in1 => \N__8496\,
            in2 => \N__7538\,
            in3 => \N__7596\,
            lcout => \U712_REG_SM.STATE_COUNTc_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__7567\,
            in1 => \N__7522\,
            in2 => \_gnd_net_\,
            in3 => \N__7941\,
            lcout => \U712_REG_SM.N_373\,
            ltout => \U712_REG_SM.N_373_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111001001110"
        )
    port map (
            in0 => \N__7456\,
            in1 => \N__8036\,
            in2 => \N__7999\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.N_130\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_ess_RNO_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10562\,
            in2 => \_gnd_net_\,
            in3 => \N__7985\,
            lcout => \U712_REG_SM.un1_REGENn_0_sqmuxa_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m37_i_o2_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010001111"
        )
    port map (
            in0 => \N__11447\,
            in1 => \N__11349\,
            in2 => \N__11149\,
            in3 => \N__11207\,
            lcout => \U712_CHIP_RAM.N_335\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_ess_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7955\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9967\,
            ce => \N__7864\,
            sr => \N__10487\
        );

    \U712_BUFFERS.N_165_i_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__11831\,
            in1 => \N__10299\,
            in2 => \_gnd_net_\,
            in3 => \N__11757\,
            lcout => \N_165_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RASn_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8179\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9925\,
            ce => 'H',
            sr => \N__10531\
        );

    \U712_CHIP_RAM.WEn_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8143\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9925\,
            ce => 'H',
            sr => \N__10531\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000001111"
        )
    port map (
            in0 => \N__11655\,
            in1 => \N__9271\,
            in2 => \N__8966\,
            in3 => \N__8737\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIE8IL_0_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8178\,
            in2 => \_gnd_net_\,
            in3 => \N__8139\,
            lcout => \U712_CHIP_RAM.N_314\,
            ltout => \U712_CHIP_RAM.N_314_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__11654\,
            in1 => \N__9270\,
            in2 => \N__8110\,
            in3 => \N__8949\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8107\,
            in1 => \N__11656\,
            in2 => \_gnd_net_\,
            in3 => \N__9604\,
            lcout => \U712_CHIP_RAM.N_361\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8942\,
            in1 => \N__11658\,
            in2 => \N__8086\,
            in3 => \N__9394\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI1HUV2_3_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10563\,
            in2 => \_gnd_net_\,
            in3 => \N__8077\,
            lcout => \U712_CHIP_RAM.un1_CMA25_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__11659\,
            in1 => \N__8071\,
            in2 => \N__8965\,
            in3 => \N__9370\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNII0RI_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11657\,
            in2 => \_gnd_net_\,
            in3 => \N__8938\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11660\,
            in1 => \N__8065\,
            in2 => \_gnd_net_\,
            in3 => \N__9382\,
            lcout => \U712_CHIP_RAM.N_367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__8053\,
            in1 => \N__11661\,
            in2 => \N__8964\,
            in3 => \N__8230\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__8817\,
            in1 => \N__10921\,
            in2 => \N__8783\,
            in3 => \N__8044\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9935\,
            ce => \N__9451\,
            sr => \N__10511\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__9358\,
            in1 => \N__8818\,
            in2 => \N__8785\,
            in3 => \N__8236\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9935\,
            ce => \N__9451\,
            sr => \N__10511\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__8819\,
            in1 => \N__10645\,
            in2 => \N__8784\,
            in3 => \N__8308\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9935\,
            ce => \N__9451\,
            sr => \N__10511\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__8551\,
            in1 => \N__10153\,
            in2 => \N__8278\,
            in3 => \N__8269\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8263\,
            in1 => \N__8245\,
            in2 => \_gnd_net_\,
            in3 => \N__8962\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8963\,
            in1 => \N__11646\,
            in2 => \N__8239\,
            in3 => \N__9658\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8673\,
            in1 => \N__10862\,
            in2 => \_gnd_net_\,
            in3 => \N__9332\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__10598\,
            sr => \N__10502\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__10861\,
            in1 => \N__8672\,
            in2 => \N__8221\,
            in3 => \N__8199\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\,
            ce => 'H',
            sr => \N__10497\
        );

    \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__8572\,
            in1 => \N__8553\,
            in2 => \_gnd_net_\,
            in3 => \N__8624\,
            lcout => \U712_CYCLE_TERM.N_332\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110111"
        )
    port map (
            in0 => \N__8574\,
            in1 => \N__8625\,
            in2 => \N__8557\,
            in3 => \N__8605\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_455_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__8626\,
            in1 => \N__10141\,
            in2 => \N__8614\,
            in3 => \N__9208\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9953\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__8573\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8552\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.START_RST_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__8463\,
            in1 => \N__8523\,
            in2 => \_gnd_net_\,
            in3 => \N__8500\,
            lcout => \U712_REG_SM.START_RSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9958\,
            ce => 'H',
            sr => \N__10489\
        );

    \U712_CHIP_RAM.CASn_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8958\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9923\,
            ce => 'H',
            sr => \N__10528\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__8752\,
            in1 => \N__8437\,
            in2 => \N__8971\,
            in3 => \N__8431\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9924\,
            ce => \N__9460\,
            sr => \N__10514\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__8751\,
            in1 => \N__9579\,
            in2 => \_gnd_net_\,
            in3 => \N__8970\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9924\,
            ce => \N__9460\,
            sr => \N__10514\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8383\,
            in1 => \N__8377\,
            in2 => \_gnd_net_\,
            in3 => \N__8371\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9924\,
            ce => \N__9460\,
            sr => \N__10514\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__8820\,
            in1 => \N__8689\,
            in2 => \N__8771\,
            in3 => \N__9103\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9926\,
            ce => \N__9459\,
            sr => \N__10508\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__8815\,
            in1 => \N__9280\,
            in2 => \N__8781\,
            in3 => \N__8986\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9926\,
            ce => \N__9459\,
            sr => \N__10508\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__8816\,
            in1 => \N__9352\,
            in2 => \N__8782\,
            in3 => \N__9052\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9926\,
            ce => \N__9459\,
            sr => \N__10508\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9021\,
            in1 => \N__8998\,
            in2 => \_gnd_net_\,
            in3 => \N__8950\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8951\,
            in1 => \N__11647\,
            in2 => \N__8989\,
            in3 => \N__9343\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__11648\,
            in1 => \N__8980\,
            in2 => \N__9403\,
            in3 => \N__8952\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__8821\,
            in1 => \N__9667\,
            in2 => \N__8788\,
            in3 => \N__8770\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9928\,
            ce => \N__9458\,
            sr => \N__10503\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__9334\,
            in1 => \_gnd_net_\,
            in2 => \N__10863\,
            in3 => \N__8679\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10633\,
            ce => \N__10602\,
            sr => \N__10499\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10857\,
            in1 => \N__10230\,
            in2 => \_gnd_net_\,
            in3 => \N__8680\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10633\,
            ce => \N__10602\,
            sr => \N__10499\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11010\,
            in1 => \N__10852\,
            in2 => \_gnd_net_\,
            in3 => \N__9649\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10633\,
            ce => \N__10602\,
            sr => \N__10499\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10690\,
            in1 => \N__9333\,
            in2 => \_gnd_net_\,
            in3 => \N__10853\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10633\,
            ce => \N__10602\,
            sr => \N__10499\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10848\,
            in1 => \N__9714\,
            in2 => \_gnd_net_\,
            in3 => \N__9821\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__10600\,
            sr => \N__10496\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10851\,
            in1 => \N__9331\,
            in2 => \_gnd_net_\,
            in3 => \N__10689\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__10600\,
            sr => \N__10496\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10846\,
            in1 => \N__9828\,
            in2 => \_gnd_net_\,
            in3 => \N__9775\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10630\,
            ce => \N__10599\,
            sr => \N__10494\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9829\,
            in1 => \N__10847\,
            in2 => \_gnd_net_\,
            in3 => \N__9707\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10630\,
            ce => \N__10599\,
            sr => \N__10494\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNI8LI41_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000111110011"
        )
    port map (
            in0 => \N__9220\,
            in1 => \N__9256\,
            in2 => \N__11841\,
            in3 => \N__11649\,
            lcout => \N_200_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.m34_i_o2_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111000111011"
        )
    port map (
            in0 => \N__11430\,
            in1 => \N__11265\,
            in2 => \N__11362\,
            in3 => \N__11096\,
            lcout => \U712_CHIP_RAM.N_337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_RNI8MQ3_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9209\,
            lcout => \CLK40_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10088\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CRCSn_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9583\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9927\,
            ce => 'H',
            sr => \N__10523\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__9520\,
            in1 => \N__9511\,
            in2 => \N__11677\,
            in3 => \N__9490\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9930\,
            ce => \N__9444\,
            sr => \N__10516\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10838\,
            in1 => \N__11011\,
            in2 => \_gnd_net_\,
            in3 => \N__10957\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__10605\,
            sr => \N__10512\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10956\,
            in1 => \N__10837\,
            in2 => \_gnd_net_\,
            in3 => \N__9715\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__10605\,
            sr => \N__10512\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10904\,
            in1 => \N__10850\,
            in2 => \_gnd_net_\,
            in3 => \N__10688\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__10603\,
            sr => \N__10506\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9645\,
            in1 => \N__10849\,
            in2 => \_gnd_net_\,
            in3 => \N__11006\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__10603\,
            sr => \N__10506\
        );

    \U712_CHIP_RAM.RAS_SYNC_1_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10102\,
            in2 => \_gnd_net_\,
            in3 => \N__10213\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_0_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__10101\,
            in1 => \N__10249\,
            in2 => \_gnd_net_\,
            in3 => \N__10237\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_2_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10103\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9988\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__9822\,
            in1 => \N__9774\,
            in2 => \_gnd_net_\,
            in3 => \N__10795\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10601\,
            sr => \N__10498\
        );

    \U712_CHIP_RAM.m40_i_o2_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010001011111"
        )
    port map (
            in0 => \N__11449\,
            in1 => \N__11363\,
            in2 => \N__11269\,
            in3 => \N__11147\,
            lcout => OPEN,
            ltout => \N_334_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_177_i_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100010011"
        )
    port map (
            in0 => \N__11653\,
            in1 => \N__11703\,
            in2 => \N__9739\,
            in3 => \N__10298\,
            lcout => \N_177_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10950\,
            in1 => \N__10774\,
            in2 => \_gnd_net_\,
            in3 => \N__9697\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10632\,
            ce => \N__10607\,
            sr => \N__10517\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10912\,
            in1 => \N__10772\,
            in2 => \_gnd_net_\,
            in3 => \N__9638\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__10606\,
            sr => \N__10513\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10895\,
            in1 => \N__10771\,
            in2 => \_gnd_net_\,
            in3 => \N__9637\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10628\,
            ce => \N__10604\,
            sr => \N__10507\
        );

    \U712_CHIP_RAM.m58_i_o2_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100011111"
        )
    port map (
            in0 => \N__11448\,
            in1 => \N__11364\,
            in2 => \N__11262\,
            in3 => \N__11148\,
            lcout => OPEN,
            ltout => \N_336_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_175_i_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__11836\,
            in1 => \N__11707\,
            in2 => \N__11680\,
            in3 => \N__11671\,
            lcout => \N_175_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.N_337_i_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110110000"
        )
    port map (
            in0 => \N__11368\,
            in1 => \N__11437\,
            in2 => \N__11140\,
            in3 => \N__11255\,
            lcout => \N_337_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.N_336_i_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011100000"
        )
    port map (
            in0 => \N__11367\,
            in1 => \N__11436\,
            in2 => \N__11139\,
            in3 => \N__11254\,
            lcout => \N_336_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.N_335_i_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001101110000"
        )
    port map (
            in0 => \N__11366\,
            in1 => \N__11435\,
            in2 => \N__11138\,
            in3 => \N__11253\,
            lcout => \N_335_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.N_334_i_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110100000"
        )
    port map (
            in0 => \N__11434\,
            in1 => \N__11365\,
            in2 => \N__11264\,
            in3 => \N__11119\,
            lcout => \N_334_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10773\,
            in1 => \N__10996\,
            in2 => \_gnd_net_\,
            in3 => \N__10949\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10631\,
            ce => \N__10609\,
            sr => \N__10524\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10911\,
            in1 => \N__10839\,
            in2 => \_gnd_net_\,
            in3 => \N__10687\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10629\,
            ce => \N__10608\,
            sr => \N__10518\
        );

    \U712_BUFFERS.DRDDIR_i_m2_LC_24_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001111111"
        )
    port map (
            in0 => \N__10390\,
            in1 => \N__10274\,
            in2 => \N__11840\,
            in3 => \N__11764\,
            lcout => \N_379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 10 2025 20:32:12

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U400_TOP" view "INTERFACE"

module U400_TOP (
    SIZ,
    MA,
    A,
    LBENn,
    CS0n,
    UUBEn,
    TAn,
    CLK40,
    RnW,
    BANK1,
    UMBEn,
    WEn,
    LLBEn,
    TSn,
    LMBEn,
    RASn,
    CS1n,
    RESETn,
    CLK_EN,
    CASn,
    BANK0);

    input [1:0] SIZ;
    output [12:0] MA;
    input [31:0] A;
    output LBENn;
    output CS0n;
    output UUBEn;
    output TAn;
    input CLK40;
    input RnW;
    output BANK1;
    output UMBEn;
    output WEn;
    output LLBEn;
    input TSn;
    output LMBEn;
    output RASn;
    output CS1n;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;

    wire N__7251;
    wire N__7250;
    wire N__7249;
    wire N__7242;
    wire N__7241;
    wire N__7240;
    wire N__7233;
    wire N__7232;
    wire N__7231;
    wire N__7224;
    wire N__7223;
    wire N__7222;
    wire N__7215;
    wire N__7214;
    wire N__7213;
    wire N__7206;
    wire N__7205;
    wire N__7204;
    wire N__7197;
    wire N__7196;
    wire N__7195;
    wire N__7188;
    wire N__7187;
    wire N__7186;
    wire N__7179;
    wire N__7178;
    wire N__7177;
    wire N__7170;
    wire N__7169;
    wire N__7168;
    wire N__7161;
    wire N__7160;
    wire N__7159;
    wire N__7152;
    wire N__7151;
    wire N__7150;
    wire N__7143;
    wire N__7142;
    wire N__7141;
    wire N__7134;
    wire N__7133;
    wire N__7132;
    wire N__7125;
    wire N__7124;
    wire N__7123;
    wire N__7116;
    wire N__7115;
    wire N__7114;
    wire N__7107;
    wire N__7106;
    wire N__7105;
    wire N__7098;
    wire N__7097;
    wire N__7096;
    wire N__7089;
    wire N__7088;
    wire N__7087;
    wire N__7080;
    wire N__7079;
    wire N__7078;
    wire N__7071;
    wire N__7070;
    wire N__7069;
    wire N__7062;
    wire N__7061;
    wire N__7060;
    wire N__7053;
    wire N__7052;
    wire N__7051;
    wire N__7044;
    wire N__7043;
    wire N__7042;
    wire N__7035;
    wire N__7034;
    wire N__7033;
    wire N__7026;
    wire N__7025;
    wire N__7024;
    wire N__7017;
    wire N__7016;
    wire N__7015;
    wire N__7008;
    wire N__7007;
    wire N__7006;
    wire N__6999;
    wire N__6998;
    wire N__6997;
    wire N__6990;
    wire N__6989;
    wire N__6988;
    wire N__6981;
    wire N__6980;
    wire N__6979;
    wire N__6972;
    wire N__6971;
    wire N__6970;
    wire N__6963;
    wire N__6962;
    wire N__6961;
    wire N__6954;
    wire N__6953;
    wire N__6952;
    wire N__6945;
    wire N__6944;
    wire N__6943;
    wire N__6936;
    wire N__6935;
    wire N__6934;
    wire N__6927;
    wire N__6926;
    wire N__6925;
    wire N__6918;
    wire N__6917;
    wire N__6916;
    wire N__6909;
    wire N__6908;
    wire N__6907;
    wire N__6900;
    wire N__6899;
    wire N__6898;
    wire N__6891;
    wire N__6890;
    wire N__6889;
    wire N__6882;
    wire N__6881;
    wire N__6880;
    wire N__6873;
    wire N__6872;
    wire N__6871;
    wire N__6864;
    wire N__6863;
    wire N__6862;
    wire N__6855;
    wire N__6854;
    wire N__6853;
    wire N__6846;
    wire N__6845;
    wire N__6844;
    wire N__6837;
    wire N__6836;
    wire N__6835;
    wire N__6828;
    wire N__6827;
    wire N__6826;
    wire N__6819;
    wire N__6818;
    wire N__6817;
    wire N__6810;
    wire N__6809;
    wire N__6808;
    wire N__6801;
    wire N__6800;
    wire N__6799;
    wire N__6792;
    wire N__6791;
    wire N__6790;
    wire N__6783;
    wire N__6782;
    wire N__6781;
    wire N__6774;
    wire N__6773;
    wire N__6772;
    wire N__6765;
    wire N__6764;
    wire N__6763;
    wire N__6756;
    wire N__6755;
    wire N__6754;
    wire N__6747;
    wire N__6746;
    wire N__6745;
    wire N__6738;
    wire N__6737;
    wire N__6736;
    wire N__6729;
    wire N__6728;
    wire N__6727;
    wire N__6720;
    wire N__6719;
    wire N__6718;
    wire N__6711;
    wire N__6710;
    wire N__6709;
    wire N__6702;
    wire N__6701;
    wire N__6700;
    wire N__6693;
    wire N__6692;
    wire N__6691;
    wire N__6684;
    wire N__6683;
    wire N__6682;
    wire N__6675;
    wire N__6674;
    wire N__6673;
    wire N__6656;
    wire N__6653;
    wire N__6650;
    wire N__6647;
    wire N__6644;
    wire N__6641;
    wire N__6638;
    wire N__6635;
    wire N__6632;
    wire N__6629;
    wire N__6626;
    wire N__6623;
    wire N__6620;
    wire N__6617;
    wire N__6616;
    wire N__6615;
    wire N__6614;
    wire N__6613;
    wire N__6612;
    wire N__6609;
    wire N__6604;
    wire N__6597;
    wire N__6596;
    wire N__6595;
    wire N__6594;
    wire N__6593;
    wire N__6592;
    wire N__6591;
    wire N__6590;
    wire N__6585;
    wire N__6582;
    wire N__6579;
    wire N__6578;
    wire N__6577;
    wire N__6576;
    wire N__6571;
    wire N__6568;
    wire N__6565;
    wire N__6560;
    wire N__6553;
    wire N__6550;
    wire N__6549;
    wire N__6544;
    wire N__6539;
    wire N__6538;
    wire N__6533;
    wire N__6530;
    wire N__6529;
    wire N__6524;
    wire N__6521;
    wire N__6518;
    wire N__6515;
    wire N__6510;
    wire N__6507;
    wire N__6502;
    wire N__6491;
    wire N__6488;
    wire N__6485;
    wire N__6482;
    wire N__6481;
    wire N__6480;
    wire N__6479;
    wire N__6476;
    wire N__6473;
    wire N__6468;
    wire N__6463;
    wire N__6462;
    wire N__6461;
    wire N__6460;
    wire N__6457;
    wire N__6456;
    wire N__6455;
    wire N__6452;
    wire N__6445;
    wire N__6442;
    wire N__6437;
    wire N__6428;
    wire N__6425;
    wire N__6422;
    wire N__6421;
    wire N__6420;
    wire N__6419;
    wire N__6418;
    wire N__6415;
    wire N__6412;
    wire N__6409;
    wire N__6406;
    wire N__6403;
    wire N__6400;
    wire N__6397;
    wire N__6392;
    wire N__6389;
    wire N__6386;
    wire N__6383;
    wire N__6378;
    wire N__6371;
    wire N__6368;
    wire N__6365;
    wire N__6364;
    wire N__6363;
    wire N__6362;
    wire N__6359;
    wire N__6358;
    wire N__6357;
    wire N__6356;
    wire N__6355;
    wire N__6354;
    wire N__6353;
    wire N__6352;
    wire N__6351;
    wire N__6350;
    wire N__6349;
    wire N__6348;
    wire N__6347;
    wire N__6346;
    wire N__6345;
    wire N__6344;
    wire N__6305;
    wire N__6302;
    wire N__6299;
    wire N__6296;
    wire N__6293;
    wire N__6290;
    wire N__6287;
    wire N__6284;
    wire N__6281;
    wire N__6278;
    wire N__6275;
    wire N__6272;
    wire N__6269;
    wire N__6266;
    wire N__6263;
    wire N__6260;
    wire N__6257;
    wire N__6254;
    wire N__6251;
    wire N__6248;
    wire N__6245;
    wire N__6242;
    wire N__6239;
    wire N__6236;
    wire N__6233;
    wire N__6230;
    wire N__6227;
    wire N__6224;
    wire N__6223;
    wire N__6220;
    wire N__6217;
    wire N__6212;
    wire N__6209;
    wire N__6206;
    wire N__6203;
    wire N__6200;
    wire N__6199;
    wire N__6194;
    wire N__6191;
    wire N__6190;
    wire N__6187;
    wire N__6186;
    wire N__6185;
    wire N__6182;
    wire N__6179;
    wire N__6174;
    wire N__6173;
    wire N__6172;
    wire N__6171;
    wire N__6170;
    wire N__6167;
    wire N__6162;
    wire N__6159;
    wire N__6156;
    wire N__6153;
    wire N__6150;
    wire N__6147;
    wire N__6140;
    wire N__6137;
    wire N__6134;
    wire N__6129;
    wire N__6126;
    wire N__6119;
    wire N__6118;
    wire N__6115;
    wire N__6114;
    wire N__6113;
    wire N__6112;
    wire N__6109;
    wire N__6106;
    wire N__6103;
    wire N__6100;
    wire N__6097;
    wire N__6094;
    wire N__6089;
    wire N__6084;
    wire N__6083;
    wire N__6082;
    wire N__6077;
    wire N__6074;
    wire N__6071;
    wire N__6068;
    wire N__6061;
    wire N__6058;
    wire N__6057;
    wire N__6052;
    wire N__6049;
    wire N__6044;
    wire N__6041;
    wire N__6038;
    wire N__6035;
    wire N__6032;
    wire N__6029;
    wire N__6026;
    wire N__6025;
    wire N__6022;
    wire N__6021;
    wire N__6018;
    wire N__6015;
    wire N__6012;
    wire N__6009;
    wire N__6004;
    wire N__6001;
    wire N__5998;
    wire N__5995;
    wire N__5992;
    wire N__5989;
    wire N__5984;
    wire N__5981;
    wire N__5980;
    wire N__5979;
    wire N__5978;
    wire N__5975;
    wire N__5972;
    wire N__5969;
    wire N__5966;
    wire N__5963;
    wire N__5960;
    wire N__5957;
    wire N__5954;
    wire N__5945;
    wire N__5942;
    wire N__5939;
    wire N__5936;
    wire N__5933;
    wire N__5932;
    wire N__5927;
    wire N__5926;
    wire N__5923;
    wire N__5920;
    wire N__5919;
    wire N__5914;
    wire N__5911;
    wire N__5908;
    wire N__5905;
    wire N__5902;
    wire N__5899;
    wire N__5894;
    wire N__5891;
    wire N__5888;
    wire N__5885;
    wire N__5882;
    wire N__5879;
    wire N__5878;
    wire N__5875;
    wire N__5874;
    wire N__5873;
    wire N__5872;
    wire N__5869;
    wire N__5868;
    wire N__5867;
    wire N__5866;
    wire N__5863;
    wire N__5862;
    wire N__5861;
    wire N__5858;
    wire N__5853;
    wire N__5850;
    wire N__5847;
    wire N__5844;
    wire N__5843;
    wire N__5840;
    wire N__5837;
    wire N__5832;
    wire N__5831;
    wire N__5828;
    wire N__5825;
    wire N__5818;
    wire N__5815;
    wire N__5808;
    wire N__5805;
    wire N__5802;
    wire N__5799;
    wire N__5796;
    wire N__5791;
    wire N__5780;
    wire N__5777;
    wire N__5774;
    wire N__5771;
    wire N__5768;
    wire N__5765;
    wire N__5764;
    wire N__5763;
    wire N__5760;
    wire N__5755;
    wire N__5754;
    wire N__5753;
    wire N__5752;
    wire N__5751;
    wire N__5748;
    wire N__5745;
    wire N__5742;
    wire N__5739;
    wire N__5736;
    wire N__5733;
    wire N__5726;
    wire N__5725;
    wire N__5724;
    wire N__5723;
    wire N__5722;
    wire N__5717;
    wire N__5714;
    wire N__5713;
    wire N__5710;
    wire N__5707;
    wire N__5702;
    wire N__5699;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5687;
    wire N__5682;
    wire N__5669;
    wire N__5668;
    wire N__5667;
    wire N__5664;
    wire N__5661;
    wire N__5658;
    wire N__5655;
    wire N__5648;
    wire N__5645;
    wire N__5642;
    wire N__5639;
    wire N__5636;
    wire N__5633;
    wire N__5630;
    wire N__5627;
    wire N__5624;
    wire N__5621;
    wire N__5618;
    wire N__5615;
    wire N__5612;
    wire N__5609;
    wire N__5606;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5594;
    wire N__5591;
    wire N__5588;
    wire N__5585;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5570;
    wire N__5567;
    wire N__5564;
    wire N__5561;
    wire N__5558;
    wire N__5555;
    wire N__5552;
    wire N__5551;
    wire N__5550;
    wire N__5547;
    wire N__5544;
    wire N__5541;
    wire N__5538;
    wire N__5531;
    wire N__5528;
    wire N__5525;
    wire N__5524;
    wire N__5523;
    wire N__5520;
    wire N__5515;
    wire N__5510;
    wire N__5509;
    wire N__5506;
    wire N__5503;
    wire N__5498;
    wire N__5497;
    wire N__5496;
    wire N__5495;
    wire N__5494;
    wire N__5493;
    wire N__5492;
    wire N__5491;
    wire N__5490;
    wire N__5489;
    wire N__5488;
    wire N__5487;
    wire N__5486;
    wire N__5485;
    wire N__5484;
    wire N__5483;
    wire N__5482;
    wire N__5481;
    wire N__5480;
    wire N__5479;
    wire N__5478;
    wire N__5477;
    wire N__5476;
    wire N__5475;
    wire N__5474;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5416;
    wire N__5413;
    wire N__5410;
    wire N__5407;
    wire N__5406;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5396;
    wire N__5393;
    wire N__5384;
    wire N__5383;
    wire N__5382;
    wire N__5381;
    wire N__5378;
    wire N__5375;
    wire N__5372;
    wire N__5369;
    wire N__5360;
    wire N__5357;
    wire N__5354;
    wire N__5351;
    wire N__5348;
    wire N__5347;
    wire N__5346;
    wire N__5343;
    wire N__5340;
    wire N__5339;
    wire N__5338;
    wire N__5337;
    wire N__5336;
    wire N__5335;
    wire N__5332;
    wire N__5327;
    wire N__5324;
    wire N__5323;
    wire N__5322;
    wire N__5319;
    wire N__5316;
    wire N__5313;
    wire N__5310;
    wire N__5309;
    wire N__5308;
    wire N__5305;
    wire N__5300;
    wire N__5297;
    wire N__5296;
    wire N__5293;
    wire N__5292;
    wire N__5289;
    wire N__5286;
    wire N__5283;
    wire N__5280;
    wire N__5277;
    wire N__5274;
    wire N__5273;
    wire N__5266;
    wire N__5263;
    wire N__5258;
    wire N__5255;
    wire N__5246;
    wire N__5241;
    wire N__5234;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5222;
    wire N__5219;
    wire N__5214;
    wire N__5211;
    wire N__5204;
    wire N__5203;
    wire N__5202;
    wire N__5199;
    wire N__5196;
    wire N__5193;
    wire N__5190;
    wire N__5183;
    wire N__5180;
    wire N__5179;
    wire N__5178;
    wire N__5175;
    wire N__5174;
    wire N__5169;
    wire N__5166;
    wire N__5165;
    wire N__5162;
    wire N__5159;
    wire N__5156;
    wire N__5153;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5137;
    wire N__5134;
    wire N__5131;
    wire N__5128;
    wire N__5123;
    wire N__5122;
    wire N__5119;
    wire N__5116;
    wire N__5111;
    wire N__5110;
    wire N__5107;
    wire N__5104;
    wire N__5101;
    wire N__5098;
    wire N__5093;
    wire N__5090;
    wire N__5087;
    wire N__5084;
    wire N__5083;
    wire N__5082;
    wire N__5081;
    wire N__5078;
    wire N__5077;
    wire N__5074;
    wire N__5069;
    wire N__5068;
    wire N__5067;
    wire N__5066;
    wire N__5063;
    wire N__5060;
    wire N__5055;
    wire N__5054;
    wire N__5053;
    wire N__5052;
    wire N__5051;
    wire N__5050;
    wire N__5049;
    wire N__5048;
    wire N__5047;
    wire N__5044;
    wire N__5039;
    wire N__5032;
    wire N__5027;
    wire N__5020;
    wire N__5017;
    wire N__5014;
    wire N__5011;
    wire N__4994;
    wire N__4991;
    wire N__4988;
    wire N__4985;
    wire N__4982;
    wire N__4979;
    wire N__4978;
    wire N__4973;
    wire N__4972;
    wire N__4971;
    wire N__4970;
    wire N__4969;
    wire N__4968;
    wire N__4965;
    wire N__4958;
    wire N__4957;
    wire N__4956;
    wire N__4953;
    wire N__4950;
    wire N__4947;
    wire N__4944;
    wire N__4939;
    wire N__4934;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4918;
    wire N__4917;
    wire N__4916;
    wire N__4915;
    wire N__4914;
    wire N__4913;
    wire N__4912;
    wire N__4909;
    wire N__4904;
    wire N__4901;
    wire N__4900;
    wire N__4897;
    wire N__4890;
    wire N__4889;
    wire N__4888;
    wire N__4881;
    wire N__4878;
    wire N__4873;
    wire N__4870;
    wire N__4867;
    wire N__4856;
    wire N__4855;
    wire N__4852;
    wire N__4847;
    wire N__4844;
    wire N__4841;
    wire N__4838;
    wire N__4835;
    wire N__4832;
    wire N__4829;
    wire N__4826;
    wire N__4823;
    wire N__4820;
    wire N__4817;
    wire N__4814;
    wire N__4813;
    wire N__4812;
    wire N__4809;
    wire N__4806;
    wire N__4805;
    wire N__4802;
    wire N__4799;
    wire N__4796;
    wire N__4793;
    wire N__4784;
    wire N__4781;
    wire N__4778;
    wire N__4777;
    wire N__4774;
    wire N__4773;
    wire N__4770;
    wire N__4767;
    wire N__4762;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4750;
    wire N__4749;
    wire N__4748;
    wire N__4745;
    wire N__4744;
    wire N__4743;
    wire N__4742;
    wire N__4741;
    wire N__4740;
    wire N__4739;
    wire N__4738;
    wire N__4737;
    wire N__4732;
    wire N__4729;
    wire N__4728;
    wire N__4727;
    wire N__4726;
    wire N__4725;
    wire N__4724;
    wire N__4721;
    wire N__4714;
    wire N__4711;
    wire N__4708;
    wire N__4703;
    wire N__4700;
    wire N__4695;
    wire N__4688;
    wire N__4685;
    wire N__4682;
    wire N__4677;
    wire N__4674;
    wire N__4655;
    wire N__4654;
    wire N__4653;
    wire N__4652;
    wire N__4651;
    wire N__4650;
    wire N__4649;
    wire N__4648;
    wire N__4647;
    wire N__4646;
    wire N__4645;
    wire N__4644;
    wire N__4643;
    wire N__4642;
    wire N__4641;
    wire N__4638;
    wire N__4635;
    wire N__4630;
    wire N__4627;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4611;
    wire N__4606;
    wire N__4605;
    wire N__4604;
    wire N__4603;
    wire N__4602;
    wire N__4601;
    wire N__4600;
    wire N__4599;
    wire N__4594;
    wire N__4589;
    wire N__4578;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4564;
    wire N__4557;
    wire N__4554;
    wire N__4553;
    wire N__4552;
    wire N__4549;
    wire N__4544;
    wire N__4541;
    wire N__4538;
    wire N__4535;
    wire N__4528;
    wire N__4523;
    wire N__4508;
    wire N__4507;
    wire N__4504;
    wire N__4503;
    wire N__4502;
    wire N__4501;
    wire N__4500;
    wire N__4497;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4484;
    wire N__4479;
    wire N__4478;
    wire N__4477;
    wire N__4476;
    wire N__4475;
    wire N__4472;
    wire N__4471;
    wire N__4470;
    wire N__4469;
    wire N__4468;
    wire N__4467;
    wire N__4464;
    wire N__4459;
    wire N__4454;
    wire N__4451;
    wire N__4446;
    wire N__4443;
    wire N__4440;
    wire N__4437;
    wire N__4434;
    wire N__4427;
    wire N__4406;
    wire N__4405;
    wire N__4404;
    wire N__4403;
    wire N__4402;
    wire N__4401;
    wire N__4400;
    wire N__4397;
    wire N__4392;
    wire N__4389;
    wire N__4388;
    wire N__4387;
    wire N__4386;
    wire N__4385;
    wire N__4384;
    wire N__4379;
    wire N__4378;
    wire N__4377;
    wire N__4374;
    wire N__4369;
    wire N__4366;
    wire N__4363;
    wire N__4360;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4348;
    wire N__4347;
    wire N__4346;
    wire N__4345;
    wire N__4344;
    wire N__4341;
    wire N__4338;
    wire N__4335;
    wire N__4328;
    wire N__4323;
    wire N__4318;
    wire N__4311;
    wire N__4306;
    wire N__4289;
    wire N__4286;
    wire N__4283;
    wire N__4280;
    wire N__4277;
    wire N__4274;
    wire N__4271;
    wire N__4268;
    wire N__4265;
    wire N__4264;
    wire N__4261;
    wire N__4258;
    wire N__4253;
    wire N__4250;
    wire N__4249;
    wire N__4248;
    wire N__4245;
    wire N__4242;
    wire N__4239;
    wire N__4232;
    wire N__4229;
    wire N__4228;
    wire N__4227;
    wire N__4224;
    wire N__4221;
    wire N__4218;
    wire N__4211;
    wire N__4208;
    wire N__4205;
    wire N__4204;
    wire N__4203;
    wire N__4202;
    wire N__4201;
    wire N__4200;
    wire N__4199;
    wire N__4198;
    wire N__4195;
    wire N__4192;
    wire N__4183;
    wire N__4178;
    wire N__4169;
    wire N__4166;
    wire N__4165;
    wire N__4162;
    wire N__4159;
    wire N__4156;
    wire N__4151;
    wire N__4150;
    wire N__4149;
    wire N__4146;
    wire N__4143;
    wire N__4140;
    wire N__4137;
    wire N__4134;
    wire N__4131;
    wire N__4124;
    wire N__4121;
    wire N__4120;
    wire N__4117;
    wire N__4114;
    wire N__4109;
    wire N__4106;
    wire N__4103;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4088;
    wire N__4085;
    wire N__4082;
    wire N__4079;
    wire N__4076;
    wire N__4073;
    wire N__4070;
    wire N__4067;
    wire N__4064;
    wire N__4061;
    wire N__4058;
    wire N__4055;
    wire N__4052;
    wire N__4051;
    wire N__4050;
    wire N__4047;
    wire N__4044;
    wire N__4041;
    wire N__4034;
    wire N__4031;
    wire N__4028;
    wire N__4025;
    wire N__4022;
    wire N__4019;
    wire N__4016;
    wire N__4015;
    wire N__4014;
    wire N__4009;
    wire N__4006;
    wire N__4001;
    wire N__3998;
    wire N__3995;
    wire N__3992;
    wire N__3989;
    wire N__3986;
    wire N__3983;
    wire N__3980;
    wire N__3977;
    wire N__3974;
    wire N__3971;
    wire N__3968;
    wire N__3965;
    wire N__3962;
    wire N__3959;
    wire N__3956;
    wire N__3953;
    wire N__3950;
    wire N__3947;
    wire N__3944;
    wire N__3941;
    wire N__3938;
    wire N__3935;
    wire N__3932;
    wire N__3929;
    wire N__3926;
    wire N__3923;
    wire N__3920;
    wire N__3917;
    wire N__3914;
    wire N__3911;
    wire N__3908;
    wire N__3905;
    wire N__3902;
    wire N__3899;
    wire N__3896;
    wire N__3893;
    wire N__3890;
    wire N__3887;
    wire N__3884;
    wire N__3881;
    wire N__3878;
    wire N__3875;
    wire N__3872;
    wire N__3869;
    wire N__3866;
    wire N__3863;
    wire N__3860;
    wire N__3857;
    wire N__3856;
    wire N__3853;
    wire N__3850;
    wire N__3845;
    wire N__3842;
    wire N__3839;
    wire N__3836;
    wire N__3833;
    wire N__3830;
    wire N__3827;
    wire N__3824;
    wire N__3823;
    wire N__3820;
    wire N__3817;
    wire N__3816;
    wire N__3813;
    wire N__3810;
    wire N__3807;
    wire N__3800;
    wire N__3797;
    wire N__3794;
    wire N__3791;
    wire N__3790;
    wire N__3789;
    wire N__3784;
    wire N__3781;
    wire N__3780;
    wire N__3777;
    wire N__3776;
    wire N__3773;
    wire N__3770;
    wire N__3767;
    wire N__3764;
    wire N__3755;
    wire N__3752;
    wire N__3749;
    wire N__3746;
    wire N__3745;
    wire N__3742;
    wire N__3739;
    wire N__3734;
    wire N__3733;
    wire N__3732;
    wire N__3727;
    wire N__3724;
    wire N__3721;
    wire N__3716;
    wire N__3713;
    wire N__3710;
    wire N__3707;
    wire N__3704;
    wire N__3701;
    wire N__3698;
    wire N__3695;
    wire N__3692;
    wire N__3689;
    wire N__3688;
    wire N__3687;
    wire N__3684;
    wire N__3681;
    wire N__3678;
    wire N__3671;
    wire N__3668;
    wire N__3667;
    wire N__3664;
    wire N__3661;
    wire N__3656;
    wire N__3655;
    wire N__3652;
    wire N__3649;
    wire N__3644;
    wire N__3641;
    wire N__3638;
    wire N__3635;
    wire N__3632;
    wire N__3631;
    wire N__3628;
    wire N__3627;
    wire N__3626;
    wire N__3625;
    wire N__3622;
    wire N__3619;
    wire N__3614;
    wire N__3613;
    wire N__3612;
    wire N__3611;
    wire N__3610;
    wire N__3607;
    wire N__3600;
    wire N__3591;
    wire N__3584;
    wire N__3581;
    wire N__3578;
    wire N__3575;
    wire N__3572;
    wire N__3569;
    wire N__3566;
    wire N__3563;
    wire N__3560;
    wire N__3559;
    wire N__3558;
    wire N__3557;
    wire N__3554;
    wire N__3549;
    wire N__3546;
    wire N__3539;
    wire N__3536;
    wire N__3533;
    wire N__3530;
    wire N__3527;
    wire N__3524;
    wire N__3521;
    wire N__3518;
    wire N__3517;
    wire N__3514;
    wire N__3511;
    wire N__3506;
    wire N__3503;
    wire N__3500;
    wire N__3497;
    wire N__3494;
    wire N__3491;
    wire N__3488;
    wire N__3485;
    wire N__3482;
    wire N__3479;
    wire N__3476;
    wire N__3473;
    wire N__3470;
    wire N__3467;
    wire N__3464;
    wire N__3461;
    wire N__3458;
    wire N__3455;
    wire N__3452;
    wire N__3449;
    wire N__3446;
    wire N__3443;
    wire N__3440;
    wire N__3437;
    wire N__3434;
    wire N__3431;
    wire N__3428;
    wire N__3425;
    wire N__3422;
    wire N__3419;
    wire N__3416;
    wire N__3413;
    wire N__3410;
    wire N__3407;
    wire N__3404;
    wire N__3401;
    wire N__3398;
    wire N__3395;
    wire N__3392;
    wire N__3389;
    wire N__3386;
    wire N__3383;
    wire N__3380;
    wire N__3377;
    wire N__3374;
    wire N__3371;
    wire N__3368;
    wire N__3365;
    wire N__3362;
    wire N__3359;
    wire N__3356;
    wire N__3353;
    wire N__3350;
    wire N__3347;
    wire N__3344;
    wire N__3341;
    wire N__3338;
    wire N__3335;
    wire N__3332;
    wire N__3331;
    wire N__3326;
    wire N__3325;
    wire N__3324;
    wire N__3321;
    wire N__3318;
    wire N__3317;
    wire N__3314;
    wire N__3311;
    wire N__3306;
    wire N__3299;
    wire N__3296;
    wire N__3293;
    wire N__3290;
    wire N__3287;
    wire N__3284;
    wire N__3283;
    wire N__3280;
    wire N__3277;
    wire N__3272;
    wire N__3269;
    wire N__3266;
    wire N__3263;
    wire N__3260;
    wire N__3257;
    wire N__3254;
    wire N__3251;
    wire N__3248;
    wire N__3245;
    wire N__3242;
    wire N__3239;
    wire N__3236;
    wire N__3233;
    wire N__3230;
    wire N__3227;
    wire N__3224;
    wire N__3221;
    wire N__3218;
    wire N__3215;
    wire N__3212;
    wire N__3209;
    wire N__3206;
    wire N__3203;
    wire N__3200;
    wire N__3197;
    wire N__3196;
    wire N__3193;
    wire N__3190;
    wire N__3185;
    wire N__3182;
    wire N__3181;
    wire N__3178;
    wire N__3173;
    wire N__3170;
    wire N__3167;
    wire N__3164;
    wire N__3161;
    wire N__3160;
    wire N__3155;
    wire N__3152;
    wire N__3149;
    wire N__3146;
    wire N__3143;
    wire N__3140;
    wire N__3137;
    wire N__3136;
    wire N__3131;
    wire N__3128;
    wire N__3125;
    wire N__3122;
    wire N__3119;
    wire N__3116;
    wire N__3113;
    wire N__3110;
    wire N__3109;
    wire N__3108;
    wire N__3105;
    wire N__3102;
    wire N__3097;
    wire N__3092;
    wire N__3089;
    wire N__3088;
    wire N__3085;
    wire N__3082;
    wire N__3077;
    wire N__3074;
    wire N__3071;
    wire N__3070;
    wire N__3067;
    wire N__3064;
    wire N__3061;
    wire N__3058;
    wire N__3053;
    wire N__3050;
    wire N__3047;
    wire N__3044;
    wire N__3041;
    wire N__3038;
    wire N__3035;
    wire N__3032;
    wire N__3029;
    wire N__3026;
    wire N__3023;
    wire N__3020;
    wire N__3017;
    wire N__3014;
    wire N__3013;
    wire N__3010;
    wire N__3007;
    wire N__3004;
    wire N__3001;
    wire N__2996;
    wire N__2993;
    wire N__2992;
    wire N__2989;
    wire N__2986;
    wire N__2981;
    wire N__2980;
    wire N__2977;
    wire N__2974;
    wire N__2969;
    wire N__2968;
    wire N__2965;
    wire N__2962;
    wire N__2957;
    wire N__2956;
    wire N__2953;
    wire N__2950;
    wire N__2945;
    wire N__2944;
    wire N__2941;
    wire N__2938;
    wire N__2933;
    wire N__2930;
    wire N__2929;
    wire N__2926;
    wire N__2923;
    wire N__2918;
    wire N__2915;
    wire N__2912;
    wire N__2909;
    wire N__2906;
    wire N__2905;
    wire N__2904;
    wire N__2901;
    wire N__2898;
    wire N__2895;
    wire N__2892;
    wire N__2885;
    wire N__2882;
    wire N__2879;
    wire N__2878;
    wire N__2875;
    wire N__2872;
    wire N__2867;
    wire N__2866;
    wire N__2865;
    wire N__2862;
    wire N__2857;
    wire N__2854;
    wire N__2849;
    wire N__2846;
    wire N__2843;
    wire N__2840;
    wire N__2837;
    wire N__2834;
    wire N__2831;
    wire N__2828;
    wire N__2825;
    wire N__2822;
    wire N__2819;
    wire N__2816;
    wire N__2813;
    wire N__2810;
    wire N__2807;
    wire N__2804;
    wire N__2803;
    wire N__2800;
    wire N__2797;
    wire N__2792;
    wire N__2789;
    wire N__2786;
    wire N__2783;
    wire N__2782;
    wire N__2779;
    wire N__2776;
    wire N__2771;
    wire N__2768;
    wire N__2765;
    wire N__2762;
    wire N__2759;
    wire N__2756;
    wire N__2753;
    wire N__2750;
    wire N__2747;
    wire N__2744;
    wire N__2743;
    wire N__2740;
    wire N__2737;
    wire N__2732;
    wire N__2731;
    wire N__2726;
    wire N__2723;
    wire N__2720;
    wire N__2717;
    wire N__2714;
    wire N__2711;
    wire N__2708;
    wire N__2705;
    wire N__2702;
    wire N__2699;
    wire CLK40_ibuf_gb_io_gb_input;
    wire GNDG0;
    wire VCCG0;
    wire \INVU400_SDRAM.REFRESH_COUNTER_1C_net ;
    wire A_c_21;
    wire BANK0_c;
    wire CONSTANT_ONE_NET;
    wire A_c_22;
    wire BANK1_c;
    wire \INVU400_SDRAM.BANK0C_net ;
    wire \INVU400_SDRAM.CS1_ENC_net ;
    wire \U400_SDRAM.un1_SDRAM_COUNTER59_0 ;
    wire \U400_SDRAM.SDRAM_CMD_5_sqmuxa ;
    wire \INVU400_SDRAM.RAM_CYCLEC_net ;
    wire RESETn_c_i;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_0 ;
    wire bfn_2_4_0_;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_2 ;
    wire \U400_SDRAM.un3_REFRESH_COUNTER_cry_1 ;
    wire \U400_SDRAM.un3_REFRESH_COUNTER_cry_2 ;
    wire \U400_SDRAM.un3_REFRESH_COUNTER_cry_3 ;
    wire \U400_SDRAM.un3_REFRESH_COUNTER_cry_4 ;
    wire \U400_SDRAM.un3_REFRESH_COUNTER_cry_5 ;
    wire \U400_SDRAM.un3_REFRESH_COUNTER_cry_6 ;
    wire \U400_SDRAM.un3_REFRESH_COUNTER_cry_7 ;
    wire \INVU400_SDRAM.REFRESH_COUNTER_2C_net ;
    wire \U400_SDRAM.SDRAM_COUNTER_RNIV59H2Z0Z_1 ;
    wire \INVU400_SDRAM.CS0_ENC_net ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_8 ;
    wire \U400_SDRAM.un1_REFRESH_COUNTERlt7_0_cascade_ ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U400_SDRAM.N_337_1_cascade_ ;
    wire \U400_SDRAM.N_64_cascade_ ;
    wire \U400_SDRAM.CS1_EN_0 ;
    wire \U400_SDRAM.N_64 ;
    wire \U400_SDRAM.N_72_cascade_ ;
    wire \U400_SDRAM.N_40 ;
    wire A_c_23;
    wire \U400_SDRAM.N_40_cascade_ ;
    wire \U400_SDRAM.CS0_EN_0 ;
    wire \U400_SDRAM.N_115 ;
    wire \U400_SDRAM.RAM_CYCLEZ0 ;
    wire \U400_SDRAM.CS1_ENZ0 ;
    wire CS1n_c;
    wire CASn_c;
    wire WEn_c;
    wire \INVU400_SDRAM.CS1nC_net ;
    wire RASn_c;
    wire \U400_SDRAM.CS0_ENZ0 ;
    wire CS0n_c;
    wire \INVU400_SDRAM.RASnC_net ;
    wire A_c_31;
    wire A_c_30;
    wire A_c_29;
    wire A_c_28;
    wire TSn_c;
    wire \U400_SDRAM.N_101 ;
    wire U400_ADDRESS_DECODE_RAM_SPACE_i_o3_2;
    wire A_c_27;
    wire U400_ADDRESS_DECODE_RAM_SPACE_i_o3_1;
    wire \INVU400_SDRAM.SDRAM_COUNTER_1C_net ;
    wire \INVU400_SDRAM.SDRAM_CONFIGUREDC_net ;
    wire \U400_SDRAM.N_113_cascade_ ;
    wire \U400_SDRAM.N_39_cascade_ ;
    wire \U400_SDRAM.SDRAM_COUNTER_1_sqmuxa_i_0_1 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_a2_1_0_0 ;
    wire \U400_SDRAM.N_78_cascade_ ;
    wire \U400_SDRAM.N_337_1 ;
    wire \U400_SDRAM.N_12_cascade_ ;
    wire \U400_SDRAM.N_91_cascade_ ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_0_0_103_i_i_a3_0_0 ;
    wire \U400_SDRAM.N_89 ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_0_0_103_i_i_0_cascade_ ;
    wire \INVU400_SDRAM.SDRAM_CMD_1C_net ;
    wire A_c_8;
    wire A_c_19;
    wire MA_c_6;
    wire A_c_6;
    wire A_c_17;
    wire MA_c_4;
    wire A_c_20;
    wire A_c_9;
    wire MA_c_7;
    wire \INVU400_SDRAM.MA_nesr_6C_net ;
    wire \U400_SDRAM.RAM_CYCLE_STARTZ0 ;
    wire \U400_SDRAM.SDRAM_COUNTER_4_sqmuxa_0_a3_0 ;
    wire RnW_c;
    wire \INVU400_SDRAM.TACKC_net ;
    wire \U400_SDRAM.N_113 ;
    wire \U400_SDRAM.N_63 ;
    wire \U400_SDRAM.N_20_cascade_ ;
    wire \U400_SDRAM.N_35 ;
    wire \U400_SDRAM.N_39 ;
    wire \U400_SDRAM.N_35_cascade_ ;
    wire \U400_SDRAM.N_44_cascade_ ;
    wire \U400_SDRAM.N_108 ;
    wire \U400_SDRAM.N_108_cascade_ ;
    wire \U400_SDRAM.N_109 ;
    wire \U400_SDRAM.N_52 ;
    wire \U400_SDRAM.SDRAM_COUNTER_s_0 ;
    wire \U400_SDRAM.N_86 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_1_0_cascade_ ;
    wire \U400_SDRAM.SDRAM_CMD_3_sqmuxa ;
    wire \U400_SDRAM.N_118 ;
    wire \U400_SDRAM.SDRAM_COUNTER_3_sqmuxa_0_a3_0_a2_0 ;
    wire \INVU400_SDRAM.SDRAM_COUNTER_0C_net ;
    wire \U400_SDRAM.N_46_cascade_ ;
    wire \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_a2_0_0_cascade_ ;
    wire \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_1_cascade_ ;
    wire \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_3 ;
    wire \U400_SDRAM.N_60 ;
    wire \U400_SDRAM.N_97_cascade_ ;
    wire \U400_SDRAM.N_20 ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_0_1_66_i_0_2_cascade_ ;
    wire A_c_18;
    wire \U400_SDRAM.N_11 ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_1 ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_3_cascade_ ;
    wire \U400_SDRAM.N_38 ;
    wire \INVU400_SDRAM.SDRAM_CMD_0C_net ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_a2_2_0_cascade_ ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_2 ;
    wire A_c_5;
    wire A_c_16;
    wire MA_c_3;
    wire A_c_26;
    wire MA_c_12;
    wire A_c_7;
    wire \U400_SDRAM.MA_5_iv_0_5 ;
    wire MA_c_5;
    wire \INVU400_SDRAM.MA_nesr_3C_net ;
    wire \U400_SDRAM.N_8_cascade_ ;
    wire \U400_SDRAM.un1_SDRAM_COUNTER59_4_i_1 ;
    wire \U400_SDRAM.N_15_cascade_ ;
    wire \U400_SDRAM.N_87 ;
    wire \U400_SDRAM.N_25 ;
    wire \U400_SDRAM.N_84 ;
    wire \U400_SDRAM.N_88 ;
    wire \U400_SDRAM.N_48 ;
    wire bfn_6_6_0_;
    wire \U400_SDRAM.SDRAM_COUNTER_s_1 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_0 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_1 ;
    wire \U400_SDRAM.SDRAM_COUNTER_s_3 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_2 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_3 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_4 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_5 ;
    wire \U400_SDRAM.N_29 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_6 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_7 ;
    wire \INVU400_SDRAM.SDRAM_COUNTER_2C_net ;
    wire \U400_SDRAM.SDRAM_COUNTERe_0_i ;
    wire \U400_SDRAM.N_336_1 ;
    wire \U400_SDRAM.N_56_cascade_ ;
    wire \U400_SDRAM.TACK_7_iv_i_0 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U400_SDRAM.N_28 ;
    wire \U400_SDRAM.N_110 ;
    wire \U400_SDRAM.WRITE_CYCLEZ0 ;
    wire \U400_SDRAM.N_13 ;
    wire \U400_SDRAM.N_44 ;
    wire \U400_SDRAM.N_8 ;
    wire \U400_SDRAM.N_13_cascade_ ;
    wire \U400_SDRAM.N_76 ;
    wire \U400_SDRAM.un1_SDRAM_COUNTER59_1_1_0 ;
    wire \U400_SDRAM.N_46 ;
    wire \U400_SDRAM.N_33_cascade_ ;
    wire \U400_SDRAM.N_67 ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_0_1_66_i_0_1 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U400_SDRAM.SDRAM_CONFIGUREDZ0 ;
    wire \U400_SDRAM.N_30 ;
    wire \U400_SDRAM.TA_COUNTER_srsts_0_a4_0_0 ;
    wire \U400_SDRAM.N_243_0 ;
    wire RESETn_c;
    wire \U400_SDRAM.TA_COUNTERZ0Z_0 ;
    wire \U400_SDRAM.N_243_0_cascade_ ;
    wire \U400_SDRAM.TACKZ0 ;
    wire \U400_SDRAM.N_241_0_en ;
    wire \U400_SDRAM.un1_TA_COUNTER_6_0_0 ;
    wire \U400_SDRAM.N_244_0 ;
    wire TA_OUT;
    wire N_53;
    wire \U400_SDRAM.TA_COUNTERZ0Z_1 ;
    wire \U400_SDRAM.TA_OUT_5_0 ;
    wire A_c_24;
    wire MA_c_11;
    wire A_c_11;
    wire MA_c_9;
    wire A_c_25;
    wire A_c_10;
    wire MA_c_8;
    wire \INVU400_SDRAM.MA_nesr_11C_net ;
    wire \U400_SDRAM.TA_COUNTERZ0Z_4 ;
    wire \U400_SDRAM.TA_COUNTERZ0Z_5 ;
    wire \U400_SDRAM.TA_COUNTERZ0Z_2 ;
    wire \U400_SDRAM.TA_COUNTERZ0Z_3 ;
    wire CLK40_c_g;
    wire \U400_SDRAM.SDRAM_CMD_1_sqmuxa_1 ;
    wire \U400_SDRAM.BURSTZ0 ;
    wire \INVU400_SDRAM.BURSTC_net ;
    wire A_c_12;
    wire MA_c_10;
    wire A_c_2;
    wire A_c_13;
    wire MA_c_0;
    wire \INVU400_SDRAM.MA_nesr_10C_net ;
    wire N_51;
    wire N_47;
    wire TA_EN_i;
    wire N_542_i;
    wire \U400_BYTE_ENABLE.N_71 ;
    wire SIZ_c_1;
    wire SIZ_c_0;
    wire \U400_BYTE_ENABLE.N_54_i ;
    wire A_c_0;
    wire RAM_SPACE_i_o3dup;
    wire \U400_BYTE_ENABLE.N_54_i_cascade_ ;
    wire A_c_1;
    wire N_49;
    wire \U400_SDRAM.SDRAM_CMDZ0Z_1 ;
    wire A_c_14;
    wire \U400_SDRAM.SDRAM_CMDZ0Z_0 ;
    wire A_c_3;
    wire \U400_SDRAM.MA_5_iv_0_1 ;
    wire MA_c_1;
    wire A_c_4;
    wire \U400_SDRAM.SDRAM_CMDZ0Z_2 ;
    wire A_c_15;
    wire \U400_SDRAM.MA20 ;
    wire MA_c_2;
    wire _gnd_net_;
    wire \INVU400_SDRAM.MA_nesr_1C_net ;
    wire \U400_SDRAM.un1_MA21_0_i_0 ;
    wire RESETn_c_i_g;

    IO_PAD MA_obuf_7_iopad (
            .OE(N__7251),
            .DIN(N__7250),
            .DOUT(N__7249),
            .PACKAGEPIN(MA[7]));
    defparam MA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_7_preio (
            .PADOEN(N__7251),
            .PADOUT(N__7250),
            .PADIN(N__7249),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3371),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__7242),
            .DIN(N__7241),
            .DOUT(N__7240),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__7242),
            .PADOUT(N__7241),
            .PADIN(N__7240),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__7233),
            .DIN(N__7232),
            .DOUT(N__7231),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__7233),
            .PADOUT(N__7232),
            .PADIN(N__7231),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3038),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__7224),
            .DIN(N__7223),
            .DOUT(N__7222),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__7224),
            .PADOUT(N__7223),
            .PADIN(N__7222),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2753),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_8_iopad (
            .OE(N__7215),
            .DIN(N__7214),
            .DOUT(N__7213),
            .PACKAGEPIN(MA[8]));
    defparam MA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_8_preio (
            .PADOEN(N__7215),
            .PADOUT(N__7214),
            .PADIN(N__7213),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5564),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_10_iopad (
            .OE(N__7206),
            .DIN(N__7205),
            .DOUT(N__7204),
            .PACKAGEPIN(MA[10]));
    defparam MA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_10_preio (
            .PADOEN(N__7206),
            .PADOUT(N__7205),
            .PADIN(N__7204),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6284),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_23_iopad (
            .OE(N__7197),
            .DIN(N__7196),
            .DOUT(N__7195),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__7197),
            .PADOUT(N__7196),
            .PADIN(N__7195),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_2_iopad (
            .OE(N__7188),
            .DIN(N__7187),
            .DOUT(N__7186),
            .PACKAGEPIN(MA[2]));
    defparam MA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_2_preio (
            .PADOEN(N__7188),
            .PADOUT(N__7187),
            .PADIN(N__7186),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6428),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__7179),
            .DIN(N__7178),
            .DOUT(N__7177),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__7179),
            .PADOUT(N__7178),
            .PADIN(N__7177),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__7170),
            .DIN(N__7169),
            .DOUT(N__7168),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__7170),
            .PADOUT(N__7169),
            .PADIN(N__7168),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__7161),
            .DIN(N__7160),
            .DOUT(N__7159),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__7161),
            .PADOUT(N__7160),
            .PADIN(N__7159),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5093),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_24_iopad (
            .OE(N__7152),
            .DIN(N__7151),
            .DOUT(N__7150),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__7152),
            .PADOUT(N__7151),
            .PADIN(N__7150),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_31_iopad (
            .OE(N__7143),
            .DIN(N__7142),
            .DOUT(N__7141),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__7143),
            .PADOUT(N__7142),
            .PADIN(N__7141),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__7134),
            .DIN(N__7133),
            .DOUT(N__7132),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__7134),
            .PADOUT(N__7133),
            .PADIN(N__7132),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_12_iopad (
            .OE(N__7125),
            .DIN(N__7124),
            .DOUT(N__7123),
            .PACKAGEPIN(MA[12]));
    defparam MA_obuf_12_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_12_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_12_preio (
            .PADOEN(N__7125),
            .PADOUT(N__7124),
            .PADIN(N__7123),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3932),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_1_iopad (
            .OE(N__7116),
            .DIN(N__7115),
            .DOUT(N__7114),
            .PACKAGEPIN(MA[1]));
    defparam MA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_1_preio (
            .PADOEN(N__7116),
            .PADOUT(N__7115),
            .PADIN(N__7114),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6638),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__7107),
            .DIN(N__7106),
            .DOUT(N__7105),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__7107),
            .PADOUT(N__7106),
            .PADIN(N__7105),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__7098),
            .DIN(N__7097),
            .DOUT(N__7096),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__7098),
            .PADOUT(N__7097),
            .PADIN(N__7096),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_21_iopad (
            .OE(N__7089),
            .DIN(N__7088),
            .DOUT(N__7087),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__7089),
            .PADOUT(N__7088),
            .PADIN(N__7087),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_4_iopad (
            .OE(N__7080),
            .DIN(N__7079),
            .DOUT(N__7078),
            .PACKAGEPIN(MA[4]));
    defparam MA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_4_preio (
            .PADOEN(N__7080),
            .PADOUT(N__7079),
            .PADIN(N__7078),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3416),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__7071),
            .DIN(N__7070),
            .DOUT(N__7069),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__7071),
            .PADOUT(N__7070),
            .PADIN(N__7069),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__7062),
            .DIN(N__7061),
            .DOUT(N__7060),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__7062),
            .PADOUT(N__7061),
            .PADIN(N__7060),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__7053),
            .DIN(N__7052),
            .DOUT(N__7051),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__7053),
            .PADOUT(N__7052),
            .PADIN(N__7051),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6236),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__7044),
            .DIN(N__7043),
            .DOUT(N__7042),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__7044),
            .PADOUT(N__7043),
            .PADIN(N__7042),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_9_iopad (
            .OE(N__7035),
            .DIN(N__7034),
            .DOUT(N__7033),
            .PACKAGEPIN(MA[9]));
    defparam MA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_9_preio (
            .PADOEN(N__7035),
            .PADOUT(N__7034),
            .PADIN(N__7033),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5600),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__7026),
            .DIN(N__7025),
            .DOUT(N__7024),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__7026),
            .PADOUT(N__7025),
            .PADIN(N__7024),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6245),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__7017),
            .DIN(N__7016),
            .DOUT(N__7015),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__7017),
            .PADOUT(N__7016),
            .PADIN(N__7015),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_29_iopad (
            .OE(N__7008),
            .DIN(N__7007),
            .DOUT(N__7006),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__7008),
            .PADOUT(N__7007),
            .PADIN(N__7006),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__6999),
            .DIN(N__6998),
            .DOUT(N__6997),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__6999),
            .PADOUT(N__6998),
            .PADIN(N__6997),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2792),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__6990),
            .DIN(N__6989),
            .DOUT(N__6988),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__6990),
            .PADOUT(N__6989),
            .PADIN(N__6988),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_22_iopad (
            .OE(N__6981),
            .DIN(N__6980),
            .DOUT(N__6979),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__6981),
            .PADOUT(N__6980),
            .PADIN(N__6979),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_3_iopad (
            .OE(N__6972),
            .DIN(N__6971),
            .DOUT(N__6970),
            .PACKAGEPIN(MA[3]));
    defparam MA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_3_preio (
            .PADOEN(N__6972),
            .PADOUT(N__6971),
            .PADIN(N__6970),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3965),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__6963),
            .DIN(N__6962),
            .DOUT(N__6961),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__6963),
            .PADOUT(N__6962),
            .PADIN(N__6961),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__6954),
            .DIN(N__6953),
            .DOUT(N__6952),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__6954),
            .PADOUT(N__6953),
            .PADIN(N__6952),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_27_iopad (
            .OE(N__6945),
            .DIN(N__6944),
            .DOUT(N__6943),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__6945),
            .PADOUT(N__6944),
            .PADIN(N__6943),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_6_iopad (
            .OE(N__6936),
            .DIN(N__6935),
            .DOUT(N__6934),
            .PACKAGEPIN(MA[6]));
    defparam MA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_6_preio (
            .PADOEN(N__6936),
            .PADOUT(N__6935),
            .PADIN(N__6934),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3449),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__6927),
            .DIN(N__6926),
            .DOUT(N__6925),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__6927),
            .PADOUT(N__6926),
            .PADIN(N__6925),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__6918),
            .DIN(N__6917),
            .DOUT(N__6916),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__6918),
            .PADOUT(N__6917),
            .PADIN(N__6916),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__6909),
            .DIN(N__6908),
            .DOUT(N__6907),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__6909),
            .PADOUT(N__6908),
            .PADIN(N__6907),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__6900),
            .DIN(N__6899),
            .DOUT(N__6898),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__6900),
            .PADOUT(N__6899),
            .PADIN(N__6898),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3299),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__6891),
            .DIN(N__6890),
            .DOUT(N__6889),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__6891),
            .PADOUT(N__6890),
            .PADIN(N__6889),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__6882),
            .DIN(N__6881),
            .DOUT(N__6880),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__6882),
            .PADOUT(N__6881),
            .PADIN(N__6880),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2816),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_11_iopad (
            .OE(N__6873),
            .DIN(N__6872),
            .DOUT(N__6871),
            .PACKAGEPIN(MA[11]));
    defparam MA_obuf_11_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_11_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_11_preio (
            .PADOEN(N__6873),
            .PADOUT(N__6872),
            .PADIN(N__6871),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5618),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TAn_obuft_iopad (
            .OE(N__6864),
            .DIN(N__6863),
            .DOUT(N__6862),
            .PACKAGEPIN(TAn));
    defparam TAn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TAn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TAn_obuft_preio (
            .PADOEN(N__6864),
            .PADOUT(N__6863),
            .PADIN(N__6862),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6212),
            .DIN0(),
            .DOUT0(N__5111),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__6855),
            .DIN(N__6854),
            .DOUT(N__6853),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__6855),
            .PADOUT(N__6854),
            .PADIN(N__6853),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_5_iopad (
            .OE(N__6846),
            .DIN(N__6845),
            .DOUT(N__6844),
            .PACKAGEPIN(MA[5]));
    defparam MA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_5_preio (
            .PADOEN(N__6846),
            .PADOUT(N__6845),
            .PADIN(N__6844),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3896),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__6837),
            .DIN(N__6836),
            .DOUT(N__6835),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__6837),
            .PADOUT(N__6836),
            .PADIN(N__6835),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__6828),
            .DIN(N__6827),
            .DOUT(N__6826),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__6828),
            .PADOUT(N__6827),
            .PADIN(N__6826),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam LBENn_obuf_iopad.PULLUP=1'b1;
    IO_PAD LBENn_obuf_iopad (
            .OE(N__6819),
            .DIN(N__6818),
            .DOUT(N__6817),
            .PACKAGEPIN(LBENn));
    defparam LBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LBENn_obuf_preio (
            .PADOEN(N__6819),
            .PADOUT(N__6818),
            .PADIN(N__6817),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5984),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_25_iopad (
            .OE(N__6810),
            .DIN(N__6809),
            .DOUT(N__6808),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__6810),
            .PADOUT(N__6809),
            .PADIN(N__6808),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CS1n_obuf_iopad (
            .OE(N__6801),
            .DIN(N__6800),
            .DOUT(N__6799),
            .PACKAGEPIN(CS1n));
    defparam CS1n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CS1n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CS1n_obuf_preio (
            .PADOEN(N__6801),
            .PADOUT(N__6800),
            .PADIN(N__6799),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3053),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__6792),
            .DIN(N__6791),
            .DOUT(N__6790),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__6792),
            .PADOUT(N__6791),
            .PADIN(N__6790),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_28_iopad (
            .OE(N__6783),
            .DIN(N__6782),
            .DOUT(N__6781),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__6783),
            .PADOUT(N__6782),
            .PADIN(N__6781),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_30_iopad (
            .OE(N__6774),
            .DIN(N__6773),
            .DOUT(N__6772),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__6774),
            .PADOUT(N__6773),
            .PADIN(N__6772),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__6765),
            .DIN(N__6764),
            .DOUT(N__6763),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__6765),
            .PADOUT(N__6764),
            .PADIN(N__6763),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__6756),
            .DIN(N__6755),
            .DOUT(N__6754),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__6756),
            .PADOUT(N__6755),
            .PADIN(N__6754),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3029),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_0_iopad (
            .OE(N__6747),
            .DIN(N__6746),
            .DOUT(N__6745),
            .PACKAGEPIN(MA[0]));
    defparam MA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_0_preio (
            .PADOEN(N__6747),
            .PADOUT(N__6746),
            .PADIN(N__6745),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6251),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__6738),
            .DIN(N__6737),
            .DOUT(N__6736),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__6738),
            .PADOUT(N__6737),
            .PADIN(N__6736),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__6729),
            .DIN(N__6728),
            .DOUT(N__6727),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__6729),
            .PADOUT(N__6728),
            .PADIN(N__6727),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__6720),
            .DIN(N__6719),
            .DOUT(N__6718),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__6720),
            .PADOUT(N__6719),
            .PADIN(N__6718),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CS0n_obuf_iopad (
            .OE(N__6711),
            .DIN(N__6710),
            .DOUT(N__6709),
            .PACKAGEPIN(CS0n));
    defparam CS0n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CS0n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CS0n_obuf_preio (
            .PADOEN(N__6711),
            .PADOUT(N__6710),
            .PADIN(N__6709),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3272),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_26_iopad (
            .OE(N__6702),
            .DIN(N__6701),
            .DOUT(N__6700),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__6702),
            .PADOUT(N__6701),
            .PADIN(N__6700),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__6693),
            .DIN(N__6692),
            .DOUT(N__6691),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__6693),
            .PADOUT(N__6692),
            .PADIN(N__6691),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5891),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__6684),
            .DIN(N__6683),
            .DOUT(N__6682),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__6684),
            .PADOUT(N__6683),
            .PADIN(N__6682),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_ibuf_gb_io_iopad (
            .OE(N__6675),
            .DIN(N__6674),
            .DOUT(N__6673),
            .PACKAGEPIN(CLK40));
    defparam CLK40_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_ibuf_gb_io_preio (
            .PADOEN(N__6675),
            .PADOUT(N__6674),
            .PADIN(N__6673),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1565 (
            .O(N__6656),
            .I(N__6653));
    LocalMux I__1564 (
            .O(N__6653),
            .I(N__6650));
    Span4Mux_h I__1563 (
            .O(N__6650),
            .I(N__6647));
    Odrv4 I__1562 (
            .O(N__6647),
            .I(A_c_3));
    InMux I__1561 (
            .O(N__6644),
            .I(N__6641));
    LocalMux I__1560 (
            .O(N__6641),
            .I(\U400_SDRAM.MA_5_iv_0_1 ));
    IoInMux I__1559 (
            .O(N__6638),
            .I(N__6635));
    LocalMux I__1558 (
            .O(N__6635),
            .I(MA_c_1));
    InMux I__1557 (
            .O(N__6632),
            .I(N__6629));
    LocalMux I__1556 (
            .O(N__6629),
            .I(N__6626));
    Span4Mux_s2_v I__1555 (
            .O(N__6626),
            .I(N__6623));
    IoSpan4Mux I__1554 (
            .O(N__6623),
            .I(N__6620));
    Odrv4 I__1553 (
            .O(N__6620),
            .I(A_c_4));
    InMux I__1552 (
            .O(N__6617),
            .I(N__6609));
    InMux I__1551 (
            .O(N__6616),
            .I(N__6604));
    InMux I__1550 (
            .O(N__6615),
            .I(N__6604));
    InMux I__1549 (
            .O(N__6614),
            .I(N__6597));
    InMux I__1548 (
            .O(N__6613),
            .I(N__6597));
    InMux I__1547 (
            .O(N__6612),
            .I(N__6597));
    LocalMux I__1546 (
            .O(N__6609),
            .I(N__6585));
    LocalMux I__1545 (
            .O(N__6604),
            .I(N__6585));
    LocalMux I__1544 (
            .O(N__6597),
            .I(N__6582));
    InMux I__1543 (
            .O(N__6596),
            .I(N__6579));
    InMux I__1542 (
            .O(N__6595),
            .I(N__6571));
    InMux I__1541 (
            .O(N__6594),
            .I(N__6571));
    InMux I__1540 (
            .O(N__6593),
            .I(N__6568));
    InMux I__1539 (
            .O(N__6592),
            .I(N__6565));
    InMux I__1538 (
            .O(N__6591),
            .I(N__6560));
    InMux I__1537 (
            .O(N__6590),
            .I(N__6560));
    Span4Mux_s1_v I__1536 (
            .O(N__6585),
            .I(N__6553));
    Span4Mux_h I__1535 (
            .O(N__6582),
            .I(N__6553));
    LocalMux I__1534 (
            .O(N__6579),
            .I(N__6553));
    CascadeMux I__1533 (
            .O(N__6578),
            .I(N__6550));
    InMux I__1532 (
            .O(N__6577),
            .I(N__6544));
    InMux I__1531 (
            .O(N__6576),
            .I(N__6544));
    LocalMux I__1530 (
            .O(N__6571),
            .I(N__6539));
    LocalMux I__1529 (
            .O(N__6568),
            .I(N__6539));
    LocalMux I__1528 (
            .O(N__6565),
            .I(N__6533));
    LocalMux I__1527 (
            .O(N__6560),
            .I(N__6533));
    Span4Mux_v I__1526 (
            .O(N__6553),
            .I(N__6530));
    InMux I__1525 (
            .O(N__6550),
            .I(N__6524));
    InMux I__1524 (
            .O(N__6549),
            .I(N__6524));
    LocalMux I__1523 (
            .O(N__6544),
            .I(N__6521));
    Span4Mux_v I__1522 (
            .O(N__6539),
            .I(N__6518));
    InMux I__1521 (
            .O(N__6538),
            .I(N__6515));
    Span4Mux_v I__1520 (
            .O(N__6533),
            .I(N__6510));
    Span4Mux_h I__1519 (
            .O(N__6530),
            .I(N__6510));
    InMux I__1518 (
            .O(N__6529),
            .I(N__6507));
    LocalMux I__1517 (
            .O(N__6524),
            .I(N__6502));
    Span12Mux_s3_v I__1516 (
            .O(N__6521),
            .I(N__6502));
    Odrv4 I__1515 (
            .O(N__6518),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1514 (
            .O(N__6515),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1513 (
            .O(N__6510),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1512 (
            .O(N__6507),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_2 ));
    Odrv12 I__1511 (
            .O(N__6502),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_2 ));
    CascadeMux I__1510 (
            .O(N__6491),
            .I(N__6488));
    InMux I__1509 (
            .O(N__6488),
            .I(N__6485));
    LocalMux I__1508 (
            .O(N__6485),
            .I(A_c_15));
    InMux I__1507 (
            .O(N__6482),
            .I(N__6476));
    InMux I__1506 (
            .O(N__6481),
            .I(N__6473));
    InMux I__1505 (
            .O(N__6480),
            .I(N__6468));
    InMux I__1504 (
            .O(N__6479),
            .I(N__6468));
    LocalMux I__1503 (
            .O(N__6476),
            .I(N__6463));
    LocalMux I__1502 (
            .O(N__6473),
            .I(N__6463));
    LocalMux I__1501 (
            .O(N__6468),
            .I(N__6457));
    Span4Mux_s2_v I__1500 (
            .O(N__6463),
            .I(N__6452));
    InMux I__1499 (
            .O(N__6462),
            .I(N__6445));
    InMux I__1498 (
            .O(N__6461),
            .I(N__6445));
    InMux I__1497 (
            .O(N__6460),
            .I(N__6445));
    Span4Mux_s2_v I__1496 (
            .O(N__6457),
            .I(N__6442));
    InMux I__1495 (
            .O(N__6456),
            .I(N__6437));
    InMux I__1494 (
            .O(N__6455),
            .I(N__6437));
    Odrv4 I__1493 (
            .O(N__6452),
            .I(\U400_SDRAM.MA20 ));
    LocalMux I__1492 (
            .O(N__6445),
            .I(\U400_SDRAM.MA20 ));
    Odrv4 I__1491 (
            .O(N__6442),
            .I(\U400_SDRAM.MA20 ));
    LocalMux I__1490 (
            .O(N__6437),
            .I(\U400_SDRAM.MA20 ));
    IoInMux I__1489 (
            .O(N__6428),
            .I(N__6425));
    LocalMux I__1488 (
            .O(N__6425),
            .I(MA_c_2));
    CEMux I__1487 (
            .O(N__6422),
            .I(N__6415));
    CEMux I__1486 (
            .O(N__6421),
            .I(N__6412));
    CEMux I__1485 (
            .O(N__6420),
            .I(N__6409));
    CEMux I__1484 (
            .O(N__6419),
            .I(N__6406));
    CEMux I__1483 (
            .O(N__6418),
            .I(N__6403));
    LocalMux I__1482 (
            .O(N__6415),
            .I(N__6400));
    LocalMux I__1481 (
            .O(N__6412),
            .I(N__6397));
    LocalMux I__1480 (
            .O(N__6409),
            .I(N__6392));
    LocalMux I__1479 (
            .O(N__6406),
            .I(N__6392));
    LocalMux I__1478 (
            .O(N__6403),
            .I(N__6389));
    Span4Mux_h I__1477 (
            .O(N__6400),
            .I(N__6386));
    Span4Mux_v I__1476 (
            .O(N__6397),
            .I(N__6383));
    Span4Mux_s2_v I__1475 (
            .O(N__6392),
            .I(N__6378));
    Span4Mux_v I__1474 (
            .O(N__6389),
            .I(N__6378));
    Odrv4 I__1473 (
            .O(N__6386),
            .I(\U400_SDRAM.un1_MA21_0_i_0 ));
    Odrv4 I__1472 (
            .O(N__6383),
            .I(\U400_SDRAM.un1_MA21_0_i_0 ));
    Odrv4 I__1471 (
            .O(N__6378),
            .I(\U400_SDRAM.un1_MA21_0_i_0 ));
    CascadeMux I__1470 (
            .O(N__6371),
            .I(N__6368));
    InMux I__1469 (
            .O(N__6368),
            .I(N__6365));
    LocalMux I__1468 (
            .O(N__6365),
            .I(N__6359));
    SRMux I__1467 (
            .O(N__6364),
            .I(N__6305));
    SRMux I__1466 (
            .O(N__6363),
            .I(N__6305));
    SRMux I__1465 (
            .O(N__6362),
            .I(N__6305));
    Glb2LocalMux I__1464 (
            .O(N__6359),
            .I(N__6305));
    SRMux I__1463 (
            .O(N__6358),
            .I(N__6305));
    SRMux I__1462 (
            .O(N__6357),
            .I(N__6305));
    SRMux I__1461 (
            .O(N__6356),
            .I(N__6305));
    SRMux I__1460 (
            .O(N__6355),
            .I(N__6305));
    SRMux I__1459 (
            .O(N__6354),
            .I(N__6305));
    SRMux I__1458 (
            .O(N__6353),
            .I(N__6305));
    SRMux I__1457 (
            .O(N__6352),
            .I(N__6305));
    SRMux I__1456 (
            .O(N__6351),
            .I(N__6305));
    SRMux I__1455 (
            .O(N__6350),
            .I(N__6305));
    SRMux I__1454 (
            .O(N__6349),
            .I(N__6305));
    SRMux I__1453 (
            .O(N__6348),
            .I(N__6305));
    SRMux I__1452 (
            .O(N__6347),
            .I(N__6305));
    SRMux I__1451 (
            .O(N__6346),
            .I(N__6305));
    SRMux I__1450 (
            .O(N__6345),
            .I(N__6305));
    SRMux I__1449 (
            .O(N__6344),
            .I(N__6305));
    GlobalMux I__1448 (
            .O(N__6305),
            .I(N__6302));
    gio2CtrlBuf I__1447 (
            .O(N__6302),
            .I(RESETn_c_i_g));
    CascadeMux I__1446 (
            .O(N__6299),
            .I(N__6296));
    InMux I__1445 (
            .O(N__6296),
            .I(N__6293));
    LocalMux I__1444 (
            .O(N__6293),
            .I(N__6290));
    Span4Mux_h I__1443 (
            .O(N__6290),
            .I(N__6287));
    Odrv4 I__1442 (
            .O(N__6287),
            .I(A_c_12));
    IoInMux I__1441 (
            .O(N__6284),
            .I(N__6281));
    LocalMux I__1440 (
            .O(N__6281),
            .I(MA_c_10));
    InMux I__1439 (
            .O(N__6278),
            .I(N__6275));
    LocalMux I__1438 (
            .O(N__6275),
            .I(N__6272));
    Span4Mux_h I__1437 (
            .O(N__6272),
            .I(N__6269));
    Odrv4 I__1436 (
            .O(N__6269),
            .I(A_c_2));
    CascadeMux I__1435 (
            .O(N__6266),
            .I(N__6263));
    InMux I__1434 (
            .O(N__6263),
            .I(N__6260));
    LocalMux I__1433 (
            .O(N__6260),
            .I(N__6257));
    Span12Mux_s5_v I__1432 (
            .O(N__6257),
            .I(N__6254));
    Odrv12 I__1431 (
            .O(N__6254),
            .I(A_c_13));
    IoInMux I__1430 (
            .O(N__6251),
            .I(N__6248));
    LocalMux I__1429 (
            .O(N__6248),
            .I(MA_c_0));
    IoInMux I__1428 (
            .O(N__6245),
            .I(N__6242));
    LocalMux I__1427 (
            .O(N__6242),
            .I(N__6239));
    Odrv4 I__1426 (
            .O(N__6239),
            .I(N_51));
    IoInMux I__1425 (
            .O(N__6236),
            .I(N__6233));
    LocalMux I__1424 (
            .O(N__6233),
            .I(N__6230));
    Odrv4 I__1423 (
            .O(N__6230),
            .I(N_47));
    InMux I__1422 (
            .O(N__6227),
            .I(N__6224));
    LocalMux I__1421 (
            .O(N__6224),
            .I(N__6220));
    InMux I__1420 (
            .O(N__6223),
            .I(N__6217));
    Odrv4 I__1419 (
            .O(N__6220),
            .I(TA_EN_i));
    LocalMux I__1418 (
            .O(N__6217),
            .I(TA_EN_i));
    IoInMux I__1417 (
            .O(N__6212),
            .I(N__6209));
    LocalMux I__1416 (
            .O(N__6209),
            .I(N__6206));
    IoSpan4Mux I__1415 (
            .O(N__6206),
            .I(N__6203));
    Odrv4 I__1414 (
            .O(N__6203),
            .I(N_542_i));
    InMux I__1413 (
            .O(N__6200),
            .I(N__6194));
    InMux I__1412 (
            .O(N__6199),
            .I(N__6194));
    LocalMux I__1411 (
            .O(N__6194),
            .I(\U400_BYTE_ENABLE.N_71 ));
    InMux I__1410 (
            .O(N__6191),
            .I(N__6187));
    InMux I__1409 (
            .O(N__6190),
            .I(N__6182));
    LocalMux I__1408 (
            .O(N__6187),
            .I(N__6179));
    InMux I__1407 (
            .O(N__6186),
            .I(N__6174));
    InMux I__1406 (
            .O(N__6185),
            .I(N__6174));
    LocalMux I__1405 (
            .O(N__6182),
            .I(N__6167));
    Span4Mux_h I__1404 (
            .O(N__6179),
            .I(N__6162));
    LocalMux I__1403 (
            .O(N__6174),
            .I(N__6162));
    InMux I__1402 (
            .O(N__6173),
            .I(N__6159));
    InMux I__1401 (
            .O(N__6172),
            .I(N__6156));
    InMux I__1400 (
            .O(N__6171),
            .I(N__6153));
    InMux I__1399 (
            .O(N__6170),
            .I(N__6150));
    Span4Mux_v I__1398 (
            .O(N__6167),
            .I(N__6147));
    Span4Mux_s3_h I__1397 (
            .O(N__6162),
            .I(N__6140));
    LocalMux I__1396 (
            .O(N__6159),
            .I(N__6140));
    LocalMux I__1395 (
            .O(N__6156),
            .I(N__6140));
    LocalMux I__1394 (
            .O(N__6153),
            .I(N__6137));
    LocalMux I__1393 (
            .O(N__6150),
            .I(N__6134));
    Span4Mux_h I__1392 (
            .O(N__6147),
            .I(N__6129));
    Span4Mux_v I__1391 (
            .O(N__6140),
            .I(N__6129));
    Span4Mux_v I__1390 (
            .O(N__6137),
            .I(N__6126));
    Odrv12 I__1389 (
            .O(N__6134),
            .I(SIZ_c_1));
    Odrv4 I__1388 (
            .O(N__6129),
            .I(SIZ_c_1));
    Odrv4 I__1387 (
            .O(N__6126),
            .I(SIZ_c_1));
    CascadeMux I__1386 (
            .O(N__6119),
            .I(N__6115));
    InMux I__1385 (
            .O(N__6118),
            .I(N__6109));
    InMux I__1384 (
            .O(N__6115),
            .I(N__6106));
    InMux I__1383 (
            .O(N__6114),
            .I(N__6103));
    CascadeMux I__1382 (
            .O(N__6113),
            .I(N__6100));
    CascadeMux I__1381 (
            .O(N__6112),
            .I(N__6097));
    LocalMux I__1380 (
            .O(N__6109),
            .I(N__6094));
    LocalMux I__1379 (
            .O(N__6106),
            .I(N__6089));
    LocalMux I__1378 (
            .O(N__6103),
            .I(N__6089));
    InMux I__1377 (
            .O(N__6100),
            .I(N__6084));
    InMux I__1376 (
            .O(N__6097),
            .I(N__6084));
    Span4Mux_s3_v I__1375 (
            .O(N__6094),
            .I(N__6077));
    Span4Mux_v I__1374 (
            .O(N__6089),
            .I(N__6077));
    LocalMux I__1373 (
            .O(N__6084),
            .I(N__6074));
    InMux I__1372 (
            .O(N__6083),
            .I(N__6071));
    CascadeMux I__1371 (
            .O(N__6082),
            .I(N__6068));
    Span4Mux_h I__1370 (
            .O(N__6077),
            .I(N__6061));
    Span4Mux_s3_v I__1369 (
            .O(N__6074),
            .I(N__6061));
    LocalMux I__1368 (
            .O(N__6071),
            .I(N__6061));
    InMux I__1367 (
            .O(N__6068),
            .I(N__6058));
    Span4Mux_s3_h I__1366 (
            .O(N__6061),
            .I(N__6052));
    LocalMux I__1365 (
            .O(N__6058),
            .I(N__6052));
    InMux I__1364 (
            .O(N__6057),
            .I(N__6049));
    Span4Mux_v I__1363 (
            .O(N__6052),
            .I(N__6044));
    LocalMux I__1362 (
            .O(N__6049),
            .I(N__6044));
    Odrv4 I__1361 (
            .O(N__6044),
            .I(SIZ_c_0));
    CascadeMux I__1360 (
            .O(N__6041),
            .I(N__6038));
    InMux I__1359 (
            .O(N__6038),
            .I(N__6035));
    LocalMux I__1358 (
            .O(N__6035),
            .I(N__6032));
    Span4Mux_v I__1357 (
            .O(N__6032),
            .I(N__6029));
    Odrv4 I__1356 (
            .O(N__6029),
            .I(\U400_BYTE_ENABLE.N_54_i ));
    InMux I__1355 (
            .O(N__6026),
            .I(N__6022));
    InMux I__1354 (
            .O(N__6025),
            .I(N__6018));
    LocalMux I__1353 (
            .O(N__6022),
            .I(N__6015));
    InMux I__1352 (
            .O(N__6021),
            .I(N__6012));
    LocalMux I__1351 (
            .O(N__6018),
            .I(N__6009));
    Span4Mux_v I__1350 (
            .O(N__6015),
            .I(N__6004));
    LocalMux I__1349 (
            .O(N__6012),
            .I(N__6004));
    Span4Mux_v I__1348 (
            .O(N__6009),
            .I(N__6001));
    Sp12to4 I__1347 (
            .O(N__6004),
            .I(N__5998));
    Span4Mux_v I__1346 (
            .O(N__6001),
            .I(N__5995));
    Span12Mux_v I__1345 (
            .O(N__5998),
            .I(N__5992));
    Span4Mux_h I__1344 (
            .O(N__5995),
            .I(N__5989));
    Odrv12 I__1343 (
            .O(N__5992),
            .I(A_c_0));
    Odrv4 I__1342 (
            .O(N__5989),
            .I(A_c_0));
    IoInMux I__1341 (
            .O(N__5984),
            .I(N__5981));
    LocalMux I__1340 (
            .O(N__5981),
            .I(N__5975));
    InMux I__1339 (
            .O(N__5980),
            .I(N__5972));
    InMux I__1338 (
            .O(N__5979),
            .I(N__5969));
    CascadeMux I__1337 (
            .O(N__5978),
            .I(N__5966));
    IoSpan4Mux I__1336 (
            .O(N__5975),
            .I(N__5963));
    LocalMux I__1335 (
            .O(N__5972),
            .I(N__5960));
    LocalMux I__1334 (
            .O(N__5969),
            .I(N__5957));
    InMux I__1333 (
            .O(N__5966),
            .I(N__5954));
    Span4Mux_s2_h I__1332 (
            .O(N__5963),
            .I(N__5945));
    Span4Mux_v I__1331 (
            .O(N__5960),
            .I(N__5945));
    Span4Mux_h I__1330 (
            .O(N__5957),
            .I(N__5945));
    LocalMux I__1329 (
            .O(N__5954),
            .I(N__5945));
    Span4Mux_v I__1328 (
            .O(N__5945),
            .I(N__5942));
    Span4Mux_h I__1327 (
            .O(N__5942),
            .I(N__5939));
    Odrv4 I__1326 (
            .O(N__5939),
            .I(RAM_SPACE_i_o3dup));
    CascadeMux I__1325 (
            .O(N__5936),
            .I(\U400_BYTE_ENABLE.N_54_i_cascade_ ));
    InMux I__1324 (
            .O(N__5933),
            .I(N__5927));
    InMux I__1323 (
            .O(N__5932),
            .I(N__5927));
    LocalMux I__1322 (
            .O(N__5927),
            .I(N__5923));
    InMux I__1321 (
            .O(N__5926),
            .I(N__5920));
    Span4Mux_v I__1320 (
            .O(N__5923),
            .I(N__5914));
    LocalMux I__1319 (
            .O(N__5920),
            .I(N__5914));
    InMux I__1318 (
            .O(N__5919),
            .I(N__5911));
    Span4Mux_v I__1317 (
            .O(N__5914),
            .I(N__5908));
    LocalMux I__1316 (
            .O(N__5911),
            .I(N__5905));
    Span4Mux_v I__1315 (
            .O(N__5908),
            .I(N__5902));
    Sp12to4 I__1314 (
            .O(N__5905),
            .I(N__5899));
    Sp12to4 I__1313 (
            .O(N__5902),
            .I(N__5894));
    Span12Mux_v I__1312 (
            .O(N__5899),
            .I(N__5894));
    Odrv12 I__1311 (
            .O(N__5894),
            .I(A_c_1));
    IoInMux I__1310 (
            .O(N__5891),
            .I(N__5888));
    LocalMux I__1309 (
            .O(N__5888),
            .I(N__5885));
    Span12Mux_s7_v I__1308 (
            .O(N__5885),
            .I(N__5882));
    Odrv12 I__1307 (
            .O(N__5882),
            .I(N_49));
    InMux I__1306 (
            .O(N__5879),
            .I(N__5875));
    CascadeMux I__1305 (
            .O(N__5878),
            .I(N__5869));
    LocalMux I__1304 (
            .O(N__5875),
            .I(N__5863));
    InMux I__1303 (
            .O(N__5874),
            .I(N__5858));
    InMux I__1302 (
            .O(N__5873),
            .I(N__5853));
    InMux I__1301 (
            .O(N__5872),
            .I(N__5853));
    InMux I__1300 (
            .O(N__5869),
            .I(N__5850));
    InMux I__1299 (
            .O(N__5868),
            .I(N__5847));
    InMux I__1298 (
            .O(N__5867),
            .I(N__5844));
    InMux I__1297 (
            .O(N__5866),
            .I(N__5840));
    Span4Mux_s1_v I__1296 (
            .O(N__5863),
            .I(N__5837));
    InMux I__1295 (
            .O(N__5862),
            .I(N__5832));
    InMux I__1294 (
            .O(N__5861),
            .I(N__5832));
    LocalMux I__1293 (
            .O(N__5858),
            .I(N__5828));
    LocalMux I__1292 (
            .O(N__5853),
            .I(N__5825));
    LocalMux I__1291 (
            .O(N__5850),
            .I(N__5818));
    LocalMux I__1290 (
            .O(N__5847),
            .I(N__5818));
    LocalMux I__1289 (
            .O(N__5844),
            .I(N__5818));
    InMux I__1288 (
            .O(N__5843),
            .I(N__5815));
    LocalMux I__1287 (
            .O(N__5840),
            .I(N__5808));
    Span4Mux_h I__1286 (
            .O(N__5837),
            .I(N__5808));
    LocalMux I__1285 (
            .O(N__5832),
            .I(N__5808));
    InMux I__1284 (
            .O(N__5831),
            .I(N__5805));
    Span4Mux_s3_h I__1283 (
            .O(N__5828),
            .I(N__5802));
    Span4Mux_s3_h I__1282 (
            .O(N__5825),
            .I(N__5799));
    Span12Mux_s8_h I__1281 (
            .O(N__5818),
            .I(N__5796));
    LocalMux I__1280 (
            .O(N__5815),
            .I(N__5791));
    Span4Mux_v I__1279 (
            .O(N__5808),
            .I(N__5791));
    LocalMux I__1278 (
            .O(N__5805),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1277 (
            .O(N__5802),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1276 (
            .O(N__5799),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_1 ));
    Odrv12 I__1275 (
            .O(N__5796),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1274 (
            .O(N__5791),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_1 ));
    CascadeMux I__1273 (
            .O(N__5780),
            .I(N__5777));
    InMux I__1272 (
            .O(N__5777),
            .I(N__5774));
    LocalMux I__1271 (
            .O(N__5774),
            .I(N__5771));
    IoSpan4Mux I__1270 (
            .O(N__5771),
            .I(N__5768));
    Odrv4 I__1269 (
            .O(N__5768),
            .I(A_c_14));
    InMux I__1268 (
            .O(N__5765),
            .I(N__5760));
    InMux I__1267 (
            .O(N__5764),
            .I(N__5755));
    InMux I__1266 (
            .O(N__5763),
            .I(N__5755));
    LocalMux I__1265 (
            .O(N__5760),
            .I(N__5748));
    LocalMux I__1264 (
            .O(N__5755),
            .I(N__5745));
    InMux I__1263 (
            .O(N__5754),
            .I(N__5742));
    InMux I__1262 (
            .O(N__5753),
            .I(N__5739));
    InMux I__1261 (
            .O(N__5752),
            .I(N__5736));
    InMux I__1260 (
            .O(N__5751),
            .I(N__5733));
    Span4Mux_s1_v I__1259 (
            .O(N__5748),
            .I(N__5726));
    Span4Mux_h I__1258 (
            .O(N__5745),
            .I(N__5726));
    LocalMux I__1257 (
            .O(N__5742),
            .I(N__5726));
    LocalMux I__1256 (
            .O(N__5739),
            .I(N__5717));
    LocalMux I__1255 (
            .O(N__5736),
            .I(N__5717));
    LocalMux I__1254 (
            .O(N__5733),
            .I(N__5714));
    Span4Mux_v I__1253 (
            .O(N__5726),
            .I(N__5710));
    InMux I__1252 (
            .O(N__5725),
            .I(N__5707));
    InMux I__1251 (
            .O(N__5724),
            .I(N__5702));
    InMux I__1250 (
            .O(N__5723),
            .I(N__5702));
    InMux I__1249 (
            .O(N__5722),
            .I(N__5699));
    Span4Mux_v I__1248 (
            .O(N__5717),
            .I(N__5696));
    Span4Mux_h I__1247 (
            .O(N__5714),
            .I(N__5693));
    InMux I__1246 (
            .O(N__5713),
            .I(N__5690));
    Span4Mux_h I__1245 (
            .O(N__5710),
            .I(N__5687));
    LocalMux I__1244 (
            .O(N__5707),
            .I(N__5682));
    LocalMux I__1243 (
            .O(N__5702),
            .I(N__5682));
    LocalMux I__1242 (
            .O(N__5699),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1241 (
            .O(N__5696),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1240 (
            .O(N__5693),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1239 (
            .O(N__5690),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1238 (
            .O(N__5687),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_0 ));
    Odrv12 I__1237 (
            .O(N__5682),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_0 ));
    InMux I__1236 (
            .O(N__5669),
            .I(N__5664));
    InMux I__1235 (
            .O(N__5668),
            .I(N__5661));
    InMux I__1234 (
            .O(N__5667),
            .I(N__5658));
    LocalMux I__1233 (
            .O(N__5664),
            .I(N__5655));
    LocalMux I__1232 (
            .O(N__5661),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_1 ));
    LocalMux I__1231 (
            .O(N__5658),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_1 ));
    Odrv4 I__1230 (
            .O(N__5655),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_1 ));
    InMux I__1229 (
            .O(N__5648),
            .I(N__5645));
    LocalMux I__1228 (
            .O(N__5645),
            .I(\U400_SDRAM.TA_OUT_5_0 ));
    CascadeMux I__1227 (
            .O(N__5642),
            .I(N__5639));
    InMux I__1226 (
            .O(N__5639),
            .I(N__5636));
    LocalMux I__1225 (
            .O(N__5636),
            .I(N__5633));
    Span4Mux_s2_v I__1224 (
            .O(N__5633),
            .I(N__5630));
    Sp12to4 I__1223 (
            .O(N__5630),
            .I(N__5627));
    Span12Mux_s10_h I__1222 (
            .O(N__5627),
            .I(N__5624));
    Span12Mux_v I__1221 (
            .O(N__5624),
            .I(N__5621));
    Odrv12 I__1220 (
            .O(N__5621),
            .I(A_c_24));
    IoInMux I__1219 (
            .O(N__5618),
            .I(N__5615));
    LocalMux I__1218 (
            .O(N__5615),
            .I(N__5612));
    Odrv4 I__1217 (
            .O(N__5612),
            .I(MA_c_11));
    InMux I__1216 (
            .O(N__5609),
            .I(N__5606));
    LocalMux I__1215 (
            .O(N__5606),
            .I(N__5603));
    Odrv12 I__1214 (
            .O(N__5603),
            .I(A_c_11));
    IoInMux I__1213 (
            .O(N__5600),
            .I(N__5597));
    LocalMux I__1212 (
            .O(N__5597),
            .I(N__5594));
    Span4Mux_s1_v I__1211 (
            .O(N__5594),
            .I(N__5591));
    Odrv4 I__1210 (
            .O(N__5591),
            .I(MA_c_9));
    InMux I__1209 (
            .O(N__5588),
            .I(N__5585));
    LocalMux I__1208 (
            .O(N__5585),
            .I(N__5582));
    Span12Mux_s11_v I__1207 (
            .O(N__5582),
            .I(N__5579));
    Odrv12 I__1206 (
            .O(N__5579),
            .I(A_c_25));
    CascadeMux I__1205 (
            .O(N__5576),
            .I(N__5573));
    InMux I__1204 (
            .O(N__5573),
            .I(N__5570));
    LocalMux I__1203 (
            .O(N__5570),
            .I(N__5567));
    Odrv12 I__1202 (
            .O(N__5567),
            .I(A_c_10));
    IoInMux I__1201 (
            .O(N__5564),
            .I(N__5561));
    LocalMux I__1200 (
            .O(N__5561),
            .I(N__5558));
    IoSpan4Mux I__1199 (
            .O(N__5558),
            .I(N__5555));
    Odrv4 I__1198 (
            .O(N__5555),
            .I(MA_c_8));
    InMux I__1197 (
            .O(N__5552),
            .I(N__5547));
    InMux I__1196 (
            .O(N__5551),
            .I(N__5544));
    InMux I__1195 (
            .O(N__5550),
            .I(N__5541));
    LocalMux I__1194 (
            .O(N__5547),
            .I(N__5538));
    LocalMux I__1193 (
            .O(N__5544),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_4 ));
    LocalMux I__1192 (
            .O(N__5541),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_4 ));
    Odrv4 I__1191 (
            .O(N__5538),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_4 ));
    InMux I__1190 (
            .O(N__5531),
            .I(N__5528));
    LocalMux I__1189 (
            .O(N__5528),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_5 ));
    InMux I__1188 (
            .O(N__5525),
            .I(N__5520));
    InMux I__1187 (
            .O(N__5524),
            .I(N__5515));
    InMux I__1186 (
            .O(N__5523),
            .I(N__5515));
    LocalMux I__1185 (
            .O(N__5520),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_2 ));
    LocalMux I__1184 (
            .O(N__5515),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_2 ));
    InMux I__1183 (
            .O(N__5510),
            .I(N__5506));
    InMux I__1182 (
            .O(N__5509),
            .I(N__5503));
    LocalMux I__1181 (
            .O(N__5506),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_3 ));
    LocalMux I__1180 (
            .O(N__5503),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_3 ));
    ClkMux I__1179 (
            .O(N__5498),
            .I(N__5423));
    ClkMux I__1178 (
            .O(N__5497),
            .I(N__5423));
    ClkMux I__1177 (
            .O(N__5496),
            .I(N__5423));
    ClkMux I__1176 (
            .O(N__5495),
            .I(N__5423));
    ClkMux I__1175 (
            .O(N__5494),
            .I(N__5423));
    ClkMux I__1174 (
            .O(N__5493),
            .I(N__5423));
    ClkMux I__1173 (
            .O(N__5492),
            .I(N__5423));
    ClkMux I__1172 (
            .O(N__5491),
            .I(N__5423));
    ClkMux I__1171 (
            .O(N__5490),
            .I(N__5423));
    ClkMux I__1170 (
            .O(N__5489),
            .I(N__5423));
    ClkMux I__1169 (
            .O(N__5488),
            .I(N__5423));
    ClkMux I__1168 (
            .O(N__5487),
            .I(N__5423));
    ClkMux I__1167 (
            .O(N__5486),
            .I(N__5423));
    ClkMux I__1166 (
            .O(N__5485),
            .I(N__5423));
    ClkMux I__1165 (
            .O(N__5484),
            .I(N__5423));
    ClkMux I__1164 (
            .O(N__5483),
            .I(N__5423));
    ClkMux I__1163 (
            .O(N__5482),
            .I(N__5423));
    ClkMux I__1162 (
            .O(N__5481),
            .I(N__5423));
    ClkMux I__1161 (
            .O(N__5480),
            .I(N__5423));
    ClkMux I__1160 (
            .O(N__5479),
            .I(N__5423));
    ClkMux I__1159 (
            .O(N__5478),
            .I(N__5423));
    ClkMux I__1158 (
            .O(N__5477),
            .I(N__5423));
    ClkMux I__1157 (
            .O(N__5476),
            .I(N__5423));
    ClkMux I__1156 (
            .O(N__5475),
            .I(N__5423));
    ClkMux I__1155 (
            .O(N__5474),
            .I(N__5423));
    GlobalMux I__1154 (
            .O(N__5423),
            .I(N__5420));
    gio2CtrlBuf I__1153 (
            .O(N__5420),
            .I(CLK40_c_g));
    InMux I__1152 (
            .O(N__5417),
            .I(N__5413));
    InMux I__1151 (
            .O(N__5416),
            .I(N__5410));
    LocalMux I__1150 (
            .O(N__5413),
            .I(N__5407));
    LocalMux I__1149 (
            .O(N__5410),
            .I(N__5402));
    Span4Mux_h I__1148 (
            .O(N__5407),
            .I(N__5399));
    InMux I__1147 (
            .O(N__5406),
            .I(N__5396));
    InMux I__1146 (
            .O(N__5405),
            .I(N__5393));
    Odrv12 I__1145 (
            .O(N__5402),
            .I(\U400_SDRAM.SDRAM_CMD_1_sqmuxa_1 ));
    Odrv4 I__1144 (
            .O(N__5399),
            .I(\U400_SDRAM.SDRAM_CMD_1_sqmuxa_1 ));
    LocalMux I__1143 (
            .O(N__5396),
            .I(\U400_SDRAM.SDRAM_CMD_1_sqmuxa_1 ));
    LocalMux I__1142 (
            .O(N__5393),
            .I(\U400_SDRAM.SDRAM_CMD_1_sqmuxa_1 ));
    InMux I__1141 (
            .O(N__5384),
            .I(N__5378));
    InMux I__1140 (
            .O(N__5383),
            .I(N__5375));
    InMux I__1139 (
            .O(N__5382),
            .I(N__5372));
    InMux I__1138 (
            .O(N__5381),
            .I(N__5369));
    LocalMux I__1137 (
            .O(N__5378),
            .I(\U400_SDRAM.BURSTZ0 ));
    LocalMux I__1136 (
            .O(N__5375),
            .I(\U400_SDRAM.BURSTZ0 ));
    LocalMux I__1135 (
            .O(N__5372),
            .I(\U400_SDRAM.BURSTZ0 ));
    LocalMux I__1134 (
            .O(N__5369),
            .I(\U400_SDRAM.BURSTZ0 ));
    InMux I__1133 (
            .O(N__5360),
            .I(N__5357));
    LocalMux I__1132 (
            .O(N__5357),
            .I(\U400_SDRAM.TA_COUNTER_srsts_0_a4_0_0 ));
    InMux I__1131 (
            .O(N__5354),
            .I(N__5351));
    LocalMux I__1130 (
            .O(N__5351),
            .I(\U400_SDRAM.N_243_0 ));
    InMux I__1129 (
            .O(N__5348),
            .I(N__5343));
    InMux I__1128 (
            .O(N__5347),
            .I(N__5340));
    InMux I__1127 (
            .O(N__5346),
            .I(N__5332));
    LocalMux I__1126 (
            .O(N__5343),
            .I(N__5327));
    LocalMux I__1125 (
            .O(N__5340),
            .I(N__5327));
    InMux I__1124 (
            .O(N__5339),
            .I(N__5324));
    CascadeMux I__1123 (
            .O(N__5338),
            .I(N__5319));
    InMux I__1122 (
            .O(N__5337),
            .I(N__5316));
    InMux I__1121 (
            .O(N__5336),
            .I(N__5313));
    CascadeMux I__1120 (
            .O(N__5335),
            .I(N__5310));
    LocalMux I__1119 (
            .O(N__5332),
            .I(N__5305));
    Span4Mux_v I__1118 (
            .O(N__5327),
            .I(N__5300));
    LocalMux I__1117 (
            .O(N__5324),
            .I(N__5300));
    InMux I__1116 (
            .O(N__5323),
            .I(N__5297));
    CascadeMux I__1115 (
            .O(N__5322),
            .I(N__5293));
    InMux I__1114 (
            .O(N__5319),
            .I(N__5289));
    LocalMux I__1113 (
            .O(N__5316),
            .I(N__5286));
    LocalMux I__1112 (
            .O(N__5313),
            .I(N__5283));
    InMux I__1111 (
            .O(N__5310),
            .I(N__5280));
    InMux I__1110 (
            .O(N__5309),
            .I(N__5277));
    CascadeMux I__1109 (
            .O(N__5308),
            .I(N__5274));
    Span4Mux_h I__1108 (
            .O(N__5305),
            .I(N__5266));
    Span4Mux_h I__1107 (
            .O(N__5300),
            .I(N__5266));
    LocalMux I__1106 (
            .O(N__5297),
            .I(N__5266));
    InMux I__1105 (
            .O(N__5296),
            .I(N__5263));
    InMux I__1104 (
            .O(N__5293),
            .I(N__5258));
    InMux I__1103 (
            .O(N__5292),
            .I(N__5258));
    LocalMux I__1102 (
            .O(N__5289),
            .I(N__5255));
    Span4Mux_h I__1101 (
            .O(N__5286),
            .I(N__5246));
    Span4Mux_v I__1100 (
            .O(N__5283),
            .I(N__5246));
    LocalMux I__1099 (
            .O(N__5280),
            .I(N__5246));
    LocalMux I__1098 (
            .O(N__5277),
            .I(N__5246));
    InMux I__1097 (
            .O(N__5274),
            .I(N__5241));
    InMux I__1096 (
            .O(N__5273),
            .I(N__5241));
    Span4Mux_h I__1095 (
            .O(N__5266),
            .I(N__5234));
    LocalMux I__1094 (
            .O(N__5263),
            .I(N__5234));
    LocalMux I__1093 (
            .O(N__5258),
            .I(N__5234));
    Sp12to4 I__1092 (
            .O(N__5255),
            .I(N__5231));
    Span4Mux_v I__1091 (
            .O(N__5246),
            .I(N__5228));
    LocalMux I__1090 (
            .O(N__5241),
            .I(N__5225));
    Span4Mux_v I__1089 (
            .O(N__5234),
            .I(N__5222));
    Span12Mux_s8_v I__1088 (
            .O(N__5231),
            .I(N__5219));
    Sp12to4 I__1087 (
            .O(N__5228),
            .I(N__5214));
    Span12Mux_s8_v I__1086 (
            .O(N__5225),
            .I(N__5214));
    Span4Mux_h I__1085 (
            .O(N__5222),
            .I(N__5211));
    Odrv12 I__1084 (
            .O(N__5219),
            .I(RESETn_c));
    Odrv12 I__1083 (
            .O(N__5214),
            .I(RESETn_c));
    Odrv4 I__1082 (
            .O(N__5211),
            .I(RESETn_c));
    InMux I__1081 (
            .O(N__5204),
            .I(N__5199));
    InMux I__1080 (
            .O(N__5203),
            .I(N__5196));
    InMux I__1079 (
            .O(N__5202),
            .I(N__5193));
    LocalMux I__1078 (
            .O(N__5199),
            .I(N__5190));
    LocalMux I__1077 (
            .O(N__5196),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_0 ));
    LocalMux I__1076 (
            .O(N__5193),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_0 ));
    Odrv4 I__1075 (
            .O(N__5190),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_0 ));
    CascadeMux I__1074 (
            .O(N__5183),
            .I(\U400_SDRAM.N_243_0_cascade_ ));
    InMux I__1073 (
            .O(N__5180),
            .I(N__5175));
    InMux I__1072 (
            .O(N__5179),
            .I(N__5169));
    InMux I__1071 (
            .O(N__5178),
            .I(N__5169));
    LocalMux I__1070 (
            .O(N__5175),
            .I(N__5166));
    InMux I__1069 (
            .O(N__5174),
            .I(N__5162));
    LocalMux I__1068 (
            .O(N__5169),
            .I(N__5159));
    Span4Mux_v I__1067 (
            .O(N__5166),
            .I(N__5156));
    InMux I__1066 (
            .O(N__5165),
            .I(N__5153));
    LocalMux I__1065 (
            .O(N__5162),
            .I(\U400_SDRAM.TACKZ0 ));
    Odrv4 I__1064 (
            .O(N__5159),
            .I(\U400_SDRAM.TACKZ0 ));
    Odrv4 I__1063 (
            .O(N__5156),
            .I(\U400_SDRAM.TACKZ0 ));
    LocalMux I__1062 (
            .O(N__5153),
            .I(\U400_SDRAM.TACKZ0 ));
    InMux I__1061 (
            .O(N__5144),
            .I(N__5141));
    LocalMux I__1060 (
            .O(N__5141),
            .I(\U400_SDRAM.N_241_0_en ));
    CascadeMux I__1059 (
            .O(N__5138),
            .I(N__5134));
    InMux I__1058 (
            .O(N__5137),
            .I(N__5131));
    InMux I__1057 (
            .O(N__5134),
            .I(N__5128));
    LocalMux I__1056 (
            .O(N__5131),
            .I(\U400_SDRAM.un1_TA_COUNTER_6_0_0 ));
    LocalMux I__1055 (
            .O(N__5128),
            .I(\U400_SDRAM.un1_TA_COUNTER_6_0_0 ));
    InMux I__1054 (
            .O(N__5123),
            .I(N__5119));
    InMux I__1053 (
            .O(N__5122),
            .I(N__5116));
    LocalMux I__1052 (
            .O(N__5119),
            .I(\U400_SDRAM.N_244_0 ));
    LocalMux I__1051 (
            .O(N__5116),
            .I(\U400_SDRAM.N_244_0 ));
    IoInMux I__1050 (
            .O(N__5111),
            .I(N__5107));
    CascadeMux I__1049 (
            .O(N__5110),
            .I(N__5104));
    LocalMux I__1048 (
            .O(N__5107),
            .I(N__5101));
    InMux I__1047 (
            .O(N__5104),
            .I(N__5098));
    Odrv12 I__1046 (
            .O(N__5101),
            .I(TA_OUT));
    LocalMux I__1045 (
            .O(N__5098),
            .I(TA_OUT));
    IoInMux I__1044 (
            .O(N__5093),
            .I(N__5090));
    LocalMux I__1043 (
            .O(N__5090),
            .I(N__5087));
    Odrv12 I__1042 (
            .O(N__5087),
            .I(N_53));
    CascadeMux I__1041 (
            .O(N__5084),
            .I(N__5078));
    InMux I__1040 (
            .O(N__5083),
            .I(N__5074));
    InMux I__1039 (
            .O(N__5082),
            .I(N__5069));
    InMux I__1038 (
            .O(N__5081),
            .I(N__5069));
    InMux I__1037 (
            .O(N__5078),
            .I(N__5063));
    InMux I__1036 (
            .O(N__5077),
            .I(N__5060));
    LocalMux I__1035 (
            .O(N__5074),
            .I(N__5055));
    LocalMux I__1034 (
            .O(N__5069),
            .I(N__5055));
    InMux I__1033 (
            .O(N__5068),
            .I(N__5044));
    InMux I__1032 (
            .O(N__5067),
            .I(N__5039));
    InMux I__1031 (
            .O(N__5066),
            .I(N__5039));
    LocalMux I__1030 (
            .O(N__5063),
            .I(N__5032));
    LocalMux I__1029 (
            .O(N__5060),
            .I(N__5032));
    Span4Mux_h I__1028 (
            .O(N__5055),
            .I(N__5032));
    InMux I__1027 (
            .O(N__5054),
            .I(N__5027));
    InMux I__1026 (
            .O(N__5053),
            .I(N__5027));
    InMux I__1025 (
            .O(N__5052),
            .I(N__5020));
    InMux I__1024 (
            .O(N__5051),
            .I(N__5020));
    InMux I__1023 (
            .O(N__5050),
            .I(N__5020));
    InMux I__1022 (
            .O(N__5049),
            .I(N__5017));
    InMux I__1021 (
            .O(N__5048),
            .I(N__5014));
    InMux I__1020 (
            .O(N__5047),
            .I(N__5011));
    LocalMux I__1019 (
            .O(N__5044),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1018 (
            .O(N__5039),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1017 (
            .O(N__5032),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1016 (
            .O(N__5027),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1015 (
            .O(N__5020),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1014 (
            .O(N__5017),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1013 (
            .O(N__5014),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1012 (
            .O(N__5011),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    InMux I__1011 (
            .O(N__4994),
            .I(N__4991));
    LocalMux I__1010 (
            .O(N__4991),
            .I(\U400_SDRAM.N_28 ));
    InMux I__1009 (
            .O(N__4988),
            .I(N__4985));
    LocalMux I__1008 (
            .O(N__4985),
            .I(\U400_SDRAM.N_110 ));
    CascadeMux I__1007 (
            .O(N__4982),
            .I(N__4979));
    InMux I__1006 (
            .O(N__4979),
            .I(N__4973));
    InMux I__1005 (
            .O(N__4978),
            .I(N__4973));
    LocalMux I__1004 (
            .O(N__4973),
            .I(N__4965));
    InMux I__1003 (
            .O(N__4972),
            .I(N__4958));
    InMux I__1002 (
            .O(N__4971),
            .I(N__4958));
    InMux I__1001 (
            .O(N__4970),
            .I(N__4958));
    InMux I__1000 (
            .O(N__4969),
            .I(N__4953));
    InMux I__999 (
            .O(N__4968),
            .I(N__4950));
    Span4Mux_h I__998 (
            .O(N__4965),
            .I(N__4947));
    LocalMux I__997 (
            .O(N__4958),
            .I(N__4944));
    InMux I__996 (
            .O(N__4957),
            .I(N__4939));
    InMux I__995 (
            .O(N__4956),
            .I(N__4939));
    LocalMux I__994 (
            .O(N__4953),
            .I(N__4934));
    LocalMux I__993 (
            .O(N__4950),
            .I(N__4934));
    Odrv4 I__992 (
            .O(N__4947),
            .I(\U400_SDRAM.WRITE_CYCLEZ0 ));
    Odrv4 I__991 (
            .O(N__4944),
            .I(\U400_SDRAM.WRITE_CYCLEZ0 ));
    LocalMux I__990 (
            .O(N__4939),
            .I(\U400_SDRAM.WRITE_CYCLEZ0 ));
    Odrv4 I__989 (
            .O(N__4934),
            .I(\U400_SDRAM.WRITE_CYCLEZ0 ));
    InMux I__988 (
            .O(N__4925),
            .I(N__4922));
    LocalMux I__987 (
            .O(N__4922),
            .I(\U400_SDRAM.N_13 ));
    InMux I__986 (
            .O(N__4919),
            .I(N__4909));
    InMux I__985 (
            .O(N__4918),
            .I(N__4904));
    InMux I__984 (
            .O(N__4917),
            .I(N__4904));
    InMux I__983 (
            .O(N__4916),
            .I(N__4901));
    InMux I__982 (
            .O(N__4915),
            .I(N__4897));
    InMux I__981 (
            .O(N__4914),
            .I(N__4890));
    InMux I__980 (
            .O(N__4913),
            .I(N__4890));
    InMux I__979 (
            .O(N__4912),
            .I(N__4890));
    LocalMux I__978 (
            .O(N__4909),
            .I(N__4881));
    LocalMux I__977 (
            .O(N__4904),
            .I(N__4881));
    LocalMux I__976 (
            .O(N__4901),
            .I(N__4881));
    InMux I__975 (
            .O(N__4900),
            .I(N__4878));
    LocalMux I__974 (
            .O(N__4897),
            .I(N__4873));
    LocalMux I__973 (
            .O(N__4890),
            .I(N__4873));
    InMux I__972 (
            .O(N__4889),
            .I(N__4870));
    InMux I__971 (
            .O(N__4888),
            .I(N__4867));
    Odrv4 I__970 (
            .O(N__4881),
            .I(\U400_SDRAM.N_44 ));
    LocalMux I__969 (
            .O(N__4878),
            .I(\U400_SDRAM.N_44 ));
    Odrv4 I__968 (
            .O(N__4873),
            .I(\U400_SDRAM.N_44 ));
    LocalMux I__967 (
            .O(N__4870),
            .I(\U400_SDRAM.N_44 ));
    LocalMux I__966 (
            .O(N__4867),
            .I(\U400_SDRAM.N_44 ));
    CascadeMux I__965 (
            .O(N__4856),
            .I(N__4852));
    InMux I__964 (
            .O(N__4855),
            .I(N__4847));
    InMux I__963 (
            .O(N__4852),
            .I(N__4847));
    LocalMux I__962 (
            .O(N__4847),
            .I(N__4844));
    Odrv12 I__961 (
            .O(N__4844),
            .I(\U400_SDRAM.N_8 ));
    CascadeMux I__960 (
            .O(N__4841),
            .I(\U400_SDRAM.N_13_cascade_ ));
    InMux I__959 (
            .O(N__4838),
            .I(N__4835));
    LocalMux I__958 (
            .O(N__4835),
            .I(N__4832));
    Span4Mux_h I__957 (
            .O(N__4832),
            .I(N__4829));
    Odrv4 I__956 (
            .O(N__4829),
            .I(\U400_SDRAM.N_76 ));
    InMux I__955 (
            .O(N__4826),
            .I(N__4823));
    LocalMux I__954 (
            .O(N__4823),
            .I(N__4820));
    Odrv12 I__953 (
            .O(N__4820),
            .I(\U400_SDRAM.un1_SDRAM_COUNTER59_1_1_0 ));
    CascadeMux I__952 (
            .O(N__4817),
            .I(N__4814));
    InMux I__951 (
            .O(N__4814),
            .I(N__4809));
    CascadeMux I__950 (
            .O(N__4813),
            .I(N__4806));
    InMux I__949 (
            .O(N__4812),
            .I(N__4802));
    LocalMux I__948 (
            .O(N__4809),
            .I(N__4799));
    InMux I__947 (
            .O(N__4806),
            .I(N__4796));
    InMux I__946 (
            .O(N__4805),
            .I(N__4793));
    LocalMux I__945 (
            .O(N__4802),
            .I(\U400_SDRAM.N_46 ));
    Odrv4 I__944 (
            .O(N__4799),
            .I(\U400_SDRAM.N_46 ));
    LocalMux I__943 (
            .O(N__4796),
            .I(\U400_SDRAM.N_46 ));
    LocalMux I__942 (
            .O(N__4793),
            .I(\U400_SDRAM.N_46 ));
    CascadeMux I__941 (
            .O(N__4784),
            .I(\U400_SDRAM.N_33_cascade_ ));
    InMux I__940 (
            .O(N__4781),
            .I(N__4778));
    LocalMux I__939 (
            .O(N__4778),
            .I(N__4774));
    CascadeMux I__938 (
            .O(N__4777),
            .I(N__4770));
    Span4Mux_v I__937 (
            .O(N__4774),
            .I(N__4767));
    InMux I__936 (
            .O(N__4773),
            .I(N__4762));
    InMux I__935 (
            .O(N__4770),
            .I(N__4762));
    Odrv4 I__934 (
            .O(N__4767),
            .I(\U400_SDRAM.N_67 ));
    LocalMux I__933 (
            .O(N__4762),
            .I(\U400_SDRAM.N_67 ));
    InMux I__932 (
            .O(N__4757),
            .I(N__4754));
    LocalMux I__931 (
            .O(N__4754),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_0_1_66_i_0_1 ));
    InMux I__930 (
            .O(N__4751),
            .I(N__4745));
    InMux I__929 (
            .O(N__4750),
            .I(N__4732));
    InMux I__928 (
            .O(N__4749),
            .I(N__4732));
    InMux I__927 (
            .O(N__4748),
            .I(N__4729));
    LocalMux I__926 (
            .O(N__4745),
            .I(N__4721));
    InMux I__925 (
            .O(N__4744),
            .I(N__4714));
    InMux I__924 (
            .O(N__4743),
            .I(N__4714));
    InMux I__923 (
            .O(N__4742),
            .I(N__4714));
    InMux I__922 (
            .O(N__4741),
            .I(N__4711));
    InMux I__921 (
            .O(N__4740),
            .I(N__4708));
    InMux I__920 (
            .O(N__4739),
            .I(N__4703));
    InMux I__919 (
            .O(N__4738),
            .I(N__4703));
    InMux I__918 (
            .O(N__4737),
            .I(N__4700));
    LocalMux I__917 (
            .O(N__4732),
            .I(N__4695));
    LocalMux I__916 (
            .O(N__4729),
            .I(N__4695));
    InMux I__915 (
            .O(N__4728),
            .I(N__4688));
    InMux I__914 (
            .O(N__4727),
            .I(N__4688));
    InMux I__913 (
            .O(N__4726),
            .I(N__4688));
    InMux I__912 (
            .O(N__4725),
            .I(N__4685));
    InMux I__911 (
            .O(N__4724),
            .I(N__4682));
    Span4Mux_h I__910 (
            .O(N__4721),
            .I(N__4677));
    LocalMux I__909 (
            .O(N__4714),
            .I(N__4677));
    LocalMux I__908 (
            .O(N__4711),
            .I(N__4674));
    LocalMux I__907 (
            .O(N__4708),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__906 (
            .O(N__4703),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__905 (
            .O(N__4700),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__904 (
            .O(N__4695),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__903 (
            .O(N__4688),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__902 (
            .O(N__4685),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__901 (
            .O(N__4682),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__900 (
            .O(N__4677),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__899 (
            .O(N__4674),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__898 (
            .O(N__4655),
            .I(N__4638));
    InMux I__897 (
            .O(N__4654),
            .I(N__4635));
    InMux I__896 (
            .O(N__4653),
            .I(N__4630));
    InMux I__895 (
            .O(N__4652),
            .I(N__4630));
    InMux I__894 (
            .O(N__4651),
            .I(N__4627));
    InMux I__893 (
            .O(N__4650),
            .I(N__4622));
    InMux I__892 (
            .O(N__4649),
            .I(N__4622));
    InMux I__891 (
            .O(N__4648),
            .I(N__4619));
    InMux I__890 (
            .O(N__4647),
            .I(N__4616));
    InMux I__889 (
            .O(N__4646),
            .I(N__4611));
    InMux I__888 (
            .O(N__4645),
            .I(N__4611));
    InMux I__887 (
            .O(N__4644),
            .I(N__4606));
    InMux I__886 (
            .O(N__4643),
            .I(N__4606));
    InMux I__885 (
            .O(N__4642),
            .I(N__4594));
    InMux I__884 (
            .O(N__4641),
            .I(N__4594));
    LocalMux I__883 (
            .O(N__4638),
            .I(N__4589));
    LocalMux I__882 (
            .O(N__4635),
            .I(N__4589));
    LocalMux I__881 (
            .O(N__4630),
            .I(N__4578));
    LocalMux I__880 (
            .O(N__4627),
            .I(N__4578));
    LocalMux I__879 (
            .O(N__4622),
            .I(N__4578));
    LocalMux I__878 (
            .O(N__4619),
            .I(N__4578));
    LocalMux I__877 (
            .O(N__4616),
            .I(N__4578));
    LocalMux I__876 (
            .O(N__4611),
            .I(N__4574));
    LocalMux I__875 (
            .O(N__4606),
            .I(N__4571));
    InMux I__874 (
            .O(N__4605),
            .I(N__4564));
    InMux I__873 (
            .O(N__4604),
            .I(N__4564));
    InMux I__872 (
            .O(N__4603),
            .I(N__4564));
    InMux I__871 (
            .O(N__4602),
            .I(N__4557));
    InMux I__870 (
            .O(N__4601),
            .I(N__4557));
    InMux I__869 (
            .O(N__4600),
            .I(N__4557));
    InMux I__868 (
            .O(N__4599),
            .I(N__4554));
    LocalMux I__867 (
            .O(N__4594),
            .I(N__4549));
    Span4Mux_v I__866 (
            .O(N__4589),
            .I(N__4544));
    Span4Mux_v I__865 (
            .O(N__4578),
            .I(N__4544));
    InMux I__864 (
            .O(N__4577),
            .I(N__4541));
    Span4Mux_s3_h I__863 (
            .O(N__4574),
            .I(N__4538));
    Span4Mux_h I__862 (
            .O(N__4571),
            .I(N__4535));
    LocalMux I__861 (
            .O(N__4564),
            .I(N__4528));
    LocalMux I__860 (
            .O(N__4557),
            .I(N__4528));
    LocalMux I__859 (
            .O(N__4554),
            .I(N__4528));
    InMux I__858 (
            .O(N__4553),
            .I(N__4523));
    InMux I__857 (
            .O(N__4552),
            .I(N__4523));
    Odrv12 I__856 (
            .O(N__4549),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__855 (
            .O(N__4544),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__854 (
            .O(N__4541),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__853 (
            .O(N__4538),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__852 (
            .O(N__4535),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__851 (
            .O(N__4528),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__850 (
            .O(N__4523),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__849 (
            .O(N__4508),
            .I(N__4504));
    CascadeMux I__848 (
            .O(N__4507),
            .I(N__4497));
    LocalMux I__847 (
            .O(N__4504),
            .I(N__4493));
    CascadeMux I__846 (
            .O(N__4503),
            .I(N__4490));
    CascadeMux I__845 (
            .O(N__4502),
            .I(N__4487));
    InMux I__844 (
            .O(N__4501),
            .I(N__4484));
    InMux I__843 (
            .O(N__4500),
            .I(N__4479));
    InMux I__842 (
            .O(N__4497),
            .I(N__4479));
    CascadeMux I__841 (
            .O(N__4496),
            .I(N__4472));
    Span4Mux_h I__840 (
            .O(N__4493),
            .I(N__4464));
    InMux I__839 (
            .O(N__4490),
            .I(N__4459));
    InMux I__838 (
            .O(N__4487),
            .I(N__4459));
    LocalMux I__837 (
            .O(N__4484),
            .I(N__4454));
    LocalMux I__836 (
            .O(N__4479),
            .I(N__4454));
    InMux I__835 (
            .O(N__4478),
            .I(N__4451));
    InMux I__834 (
            .O(N__4477),
            .I(N__4446));
    InMux I__833 (
            .O(N__4476),
            .I(N__4446));
    InMux I__832 (
            .O(N__4475),
            .I(N__4443));
    InMux I__831 (
            .O(N__4472),
            .I(N__4440));
    InMux I__830 (
            .O(N__4471),
            .I(N__4437));
    InMux I__829 (
            .O(N__4470),
            .I(N__4434));
    InMux I__828 (
            .O(N__4469),
            .I(N__4427));
    InMux I__827 (
            .O(N__4468),
            .I(N__4427));
    InMux I__826 (
            .O(N__4467),
            .I(N__4427));
    Odrv4 I__825 (
            .O(N__4464),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__824 (
            .O(N__4459),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__823 (
            .O(N__4454),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__822 (
            .O(N__4451),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__821 (
            .O(N__4446),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__820 (
            .O(N__4443),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__819 (
            .O(N__4440),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__818 (
            .O(N__4437),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__817 (
            .O(N__4434),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__816 (
            .O(N__4427),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    InMux I__815 (
            .O(N__4406),
            .I(N__4397));
    InMux I__814 (
            .O(N__4405),
            .I(N__4392));
    InMux I__813 (
            .O(N__4404),
            .I(N__4392));
    InMux I__812 (
            .O(N__4403),
            .I(N__4389));
    InMux I__811 (
            .O(N__4402),
            .I(N__4379));
    InMux I__810 (
            .O(N__4401),
            .I(N__4379));
    InMux I__809 (
            .O(N__4400),
            .I(N__4374));
    LocalMux I__808 (
            .O(N__4397),
            .I(N__4369));
    LocalMux I__807 (
            .O(N__4392),
            .I(N__4369));
    LocalMux I__806 (
            .O(N__4389),
            .I(N__4366));
    InMux I__805 (
            .O(N__4388),
            .I(N__4363));
    InMux I__804 (
            .O(N__4387),
            .I(N__4360));
    InMux I__803 (
            .O(N__4386),
            .I(N__4355));
    InMux I__802 (
            .O(N__4385),
            .I(N__4355));
    InMux I__801 (
            .O(N__4384),
            .I(N__4352));
    LocalMux I__800 (
            .O(N__4379),
            .I(N__4349));
    InMux I__799 (
            .O(N__4378),
            .I(N__4341));
    InMux I__798 (
            .O(N__4377),
            .I(N__4338));
    LocalMux I__797 (
            .O(N__4374),
            .I(N__4335));
    Span4Mux_v I__796 (
            .O(N__4369),
            .I(N__4328));
    Span4Mux_v I__795 (
            .O(N__4366),
            .I(N__4328));
    LocalMux I__794 (
            .O(N__4363),
            .I(N__4328));
    LocalMux I__793 (
            .O(N__4360),
            .I(N__4323));
    LocalMux I__792 (
            .O(N__4355),
            .I(N__4323));
    LocalMux I__791 (
            .O(N__4352),
            .I(N__4318));
    Span4Mux_h I__790 (
            .O(N__4349),
            .I(N__4318));
    InMux I__789 (
            .O(N__4348),
            .I(N__4311));
    InMux I__788 (
            .O(N__4347),
            .I(N__4311));
    InMux I__787 (
            .O(N__4346),
            .I(N__4311));
    InMux I__786 (
            .O(N__4345),
            .I(N__4306));
    InMux I__785 (
            .O(N__4344),
            .I(N__4306));
    LocalMux I__784 (
            .O(N__4341),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__783 (
            .O(N__4338),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__782 (
            .O(N__4335),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__781 (
            .O(N__4328),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__780 (
            .O(N__4323),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__779 (
            .O(N__4318),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__778 (
            .O(N__4311),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__777 (
            .O(N__4306),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    InMux I__776 (
            .O(N__4289),
            .I(N__4286));
    LocalMux I__775 (
            .O(N__4286),
            .I(\U400_SDRAM.N_30 ));
    InMux I__774 (
            .O(N__4283),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_0 ));
    InMux I__773 (
            .O(N__4280),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_1 ));
    CascadeMux I__772 (
            .O(N__4277),
            .I(N__4274));
    InMux I__771 (
            .O(N__4274),
            .I(N__4271));
    LocalMux I__770 (
            .O(N__4271),
            .I(\U400_SDRAM.SDRAM_COUNTER_s_3 ));
    InMux I__769 (
            .O(N__4268),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_2 ));
    InMux I__768 (
            .O(N__4265),
            .I(N__4261));
    InMux I__767 (
            .O(N__4264),
            .I(N__4258));
    LocalMux I__766 (
            .O(N__4261),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__765 (
            .O(N__4258),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__764 (
            .O(N__4253),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_3 ));
    InMux I__763 (
            .O(N__4250),
            .I(N__4245));
    InMux I__762 (
            .O(N__4249),
            .I(N__4242));
    InMux I__761 (
            .O(N__4248),
            .I(N__4239));
    LocalMux I__760 (
            .O(N__4245),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__759 (
            .O(N__4242),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__758 (
            .O(N__4239),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_5 ));
    InMux I__757 (
            .O(N__4232),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_4 ));
    InMux I__756 (
            .O(N__4229),
            .I(N__4224));
    InMux I__755 (
            .O(N__4228),
            .I(N__4221));
    InMux I__754 (
            .O(N__4227),
            .I(N__4218));
    LocalMux I__753 (
            .O(N__4224),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__752 (
            .O(N__4221),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__751 (
            .O(N__4218),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__750 (
            .O(N__4211),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_5 ));
    InMux I__749 (
            .O(N__4208),
            .I(N__4205));
    LocalMux I__748 (
            .O(N__4205),
            .I(N__4195));
    InMux I__747 (
            .O(N__4204),
            .I(N__4192));
    InMux I__746 (
            .O(N__4203),
            .I(N__4183));
    InMux I__745 (
            .O(N__4202),
            .I(N__4183));
    InMux I__744 (
            .O(N__4201),
            .I(N__4183));
    InMux I__743 (
            .O(N__4200),
            .I(N__4183));
    InMux I__742 (
            .O(N__4199),
            .I(N__4178));
    InMux I__741 (
            .O(N__4198),
            .I(N__4178));
    Odrv4 I__740 (
            .O(N__4195),
            .I(\U400_SDRAM.N_29 ));
    LocalMux I__739 (
            .O(N__4192),
            .I(\U400_SDRAM.N_29 ));
    LocalMux I__738 (
            .O(N__4183),
            .I(\U400_SDRAM.N_29 ));
    LocalMux I__737 (
            .O(N__4178),
            .I(\U400_SDRAM.N_29 ));
    InMux I__736 (
            .O(N__4169),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_6 ));
    CascadeMux I__735 (
            .O(N__4166),
            .I(N__4162));
    InMux I__734 (
            .O(N__4165),
            .I(N__4159));
    InMux I__733 (
            .O(N__4162),
            .I(N__4156));
    LocalMux I__732 (
            .O(N__4159),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__731 (
            .O(N__4156),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_7 ));
    CEMux I__730 (
            .O(N__4151),
            .I(N__4146));
    CEMux I__729 (
            .O(N__4150),
            .I(N__4143));
    CEMux I__728 (
            .O(N__4149),
            .I(N__4140));
    LocalMux I__727 (
            .O(N__4146),
            .I(N__4137));
    LocalMux I__726 (
            .O(N__4143),
            .I(N__4134));
    LocalMux I__725 (
            .O(N__4140),
            .I(N__4131));
    Span4Mux_v I__724 (
            .O(N__4137),
            .I(N__4124));
    Span4Mux_h I__723 (
            .O(N__4134),
            .I(N__4124));
    Span4Mux_h I__722 (
            .O(N__4131),
            .I(N__4124));
    Odrv4 I__721 (
            .O(N__4124),
            .I(\U400_SDRAM.SDRAM_COUNTERe_0_i ));
    InMux I__720 (
            .O(N__4121),
            .I(N__4117));
    InMux I__719 (
            .O(N__4120),
            .I(N__4114));
    LocalMux I__718 (
            .O(N__4117),
            .I(\U400_SDRAM.N_336_1 ));
    LocalMux I__717 (
            .O(N__4114),
            .I(\U400_SDRAM.N_336_1 ));
    CascadeMux I__716 (
            .O(N__4109),
            .I(\U400_SDRAM.N_56_cascade_ ));
    CascadeMux I__715 (
            .O(N__4106),
            .I(N__4103));
    InMux I__714 (
            .O(N__4103),
            .I(N__4100));
    LocalMux I__713 (
            .O(N__4100),
            .I(N__4097));
    Span4Mux_h I__712 (
            .O(N__4097),
            .I(N__4094));
    Odrv4 I__711 (
            .O(N__4094),
            .I(\U400_SDRAM.TACK_7_iv_i_0 ));
    CascadeMux I__710 (
            .O(N__4091),
            .I(\U400_SDRAM.N_8_cascade_ ));
    InMux I__709 (
            .O(N__4088),
            .I(N__4085));
    LocalMux I__708 (
            .O(N__4085),
            .I(\U400_SDRAM.un1_SDRAM_COUNTER59_4_i_1 ));
    CascadeMux I__707 (
            .O(N__4082),
            .I(\U400_SDRAM.N_15_cascade_ ));
    InMux I__706 (
            .O(N__4079),
            .I(N__4076));
    LocalMux I__705 (
            .O(N__4076),
            .I(N__4073));
    Odrv4 I__704 (
            .O(N__4073),
            .I(\U400_SDRAM.N_87 ));
    InMux I__703 (
            .O(N__4070),
            .I(N__4067));
    LocalMux I__702 (
            .O(N__4067),
            .I(\U400_SDRAM.N_25 ));
    InMux I__701 (
            .O(N__4064),
            .I(N__4061));
    LocalMux I__700 (
            .O(N__4061),
            .I(\U400_SDRAM.N_84 ));
    InMux I__699 (
            .O(N__4058),
            .I(N__4055));
    LocalMux I__698 (
            .O(N__4055),
            .I(\U400_SDRAM.N_88 ));
    InMux I__697 (
            .O(N__4052),
            .I(N__4047));
    InMux I__696 (
            .O(N__4051),
            .I(N__4044));
    InMux I__695 (
            .O(N__4050),
            .I(N__4041));
    LocalMux I__694 (
            .O(N__4047),
            .I(\U400_SDRAM.N_48 ));
    LocalMux I__693 (
            .O(N__4044),
            .I(\U400_SDRAM.N_48 ));
    LocalMux I__692 (
            .O(N__4041),
            .I(\U400_SDRAM.N_48 ));
    CascadeMux I__691 (
            .O(N__4034),
            .I(N__4031));
    InMux I__690 (
            .O(N__4031),
            .I(N__4028));
    LocalMux I__689 (
            .O(N__4028),
            .I(N__4025));
    Span4Mux_h I__688 (
            .O(N__4025),
            .I(N__4022));
    Odrv4 I__687 (
            .O(N__4022),
            .I(\U400_SDRAM.SDRAM_COUNTER_s_1 ));
    CascadeMux I__686 (
            .O(N__4019),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_3_cascade_ ));
    InMux I__685 (
            .O(N__4016),
            .I(N__4009));
    InMux I__684 (
            .O(N__4015),
            .I(N__4009));
    InMux I__683 (
            .O(N__4014),
            .I(N__4006));
    LocalMux I__682 (
            .O(N__4009),
            .I(\U400_SDRAM.N_38 ));
    LocalMux I__681 (
            .O(N__4006),
            .I(\U400_SDRAM.N_38 ));
    CascadeMux I__680 (
            .O(N__4001),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_a2_2_0_cascade_ ));
    InMux I__679 (
            .O(N__3998),
            .I(N__3995));
    LocalMux I__678 (
            .O(N__3995),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_2 ));
    InMux I__677 (
            .O(N__3992),
            .I(N__3989));
    LocalMux I__676 (
            .O(N__3989),
            .I(N__3986));
    Odrv12 I__675 (
            .O(N__3986),
            .I(A_c_5));
    InMux I__674 (
            .O(N__3983),
            .I(N__3980));
    LocalMux I__673 (
            .O(N__3980),
            .I(N__3977));
    Span4Mux_v I__672 (
            .O(N__3977),
            .I(N__3974));
    Span4Mux_v I__671 (
            .O(N__3974),
            .I(N__3971));
    Sp12to4 I__670 (
            .O(N__3971),
            .I(N__3968));
    Odrv12 I__669 (
            .O(N__3968),
            .I(A_c_16));
    IoInMux I__668 (
            .O(N__3965),
            .I(N__3962));
    LocalMux I__667 (
            .O(N__3962),
            .I(N__3959));
    Span12Mux_s3_v I__666 (
            .O(N__3959),
            .I(N__3956));
    Odrv12 I__665 (
            .O(N__3956),
            .I(MA_c_3));
    CascadeMux I__664 (
            .O(N__3953),
            .I(N__3950));
    InMux I__663 (
            .O(N__3950),
            .I(N__3947));
    LocalMux I__662 (
            .O(N__3947),
            .I(N__3944));
    Span4Mux_h I__661 (
            .O(N__3944),
            .I(N__3941));
    Sp12to4 I__660 (
            .O(N__3941),
            .I(N__3938));
    Span12Mux_v I__659 (
            .O(N__3938),
            .I(N__3935));
    Odrv12 I__658 (
            .O(N__3935),
            .I(A_c_26));
    IoInMux I__657 (
            .O(N__3932),
            .I(N__3929));
    LocalMux I__656 (
            .O(N__3929),
            .I(N__3926));
    Span4Mux_s0_v I__655 (
            .O(N__3926),
            .I(N__3923));
    Odrv4 I__654 (
            .O(N__3923),
            .I(MA_c_12));
    InMux I__653 (
            .O(N__3920),
            .I(N__3917));
    LocalMux I__652 (
            .O(N__3917),
            .I(N__3914));
    Span4Mux_v I__651 (
            .O(N__3914),
            .I(N__3911));
    Span4Mux_h I__650 (
            .O(N__3911),
            .I(N__3908));
    Odrv4 I__649 (
            .O(N__3908),
            .I(A_c_7));
    InMux I__648 (
            .O(N__3905),
            .I(N__3902));
    LocalMux I__647 (
            .O(N__3902),
            .I(N__3899));
    Odrv12 I__646 (
            .O(N__3899),
            .I(\U400_SDRAM.MA_5_iv_0_5 ));
    IoInMux I__645 (
            .O(N__3896),
            .I(N__3893));
    LocalMux I__644 (
            .O(N__3893),
            .I(N__3890));
    Span4Mux_s3_v I__643 (
            .O(N__3890),
            .I(N__3887));
    Odrv4 I__642 (
            .O(N__3887),
            .I(MA_c_5));
    CascadeMux I__641 (
            .O(N__3884),
            .I(\U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_a2_0_0_cascade_ ));
    CascadeMux I__640 (
            .O(N__3881),
            .I(\U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_1_cascade_ ));
    InMux I__639 (
            .O(N__3878),
            .I(N__3875));
    LocalMux I__638 (
            .O(N__3875),
            .I(\U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_3 ));
    CascadeMux I__637 (
            .O(N__3872),
            .I(N__3869));
    InMux I__636 (
            .O(N__3869),
            .I(N__3866));
    LocalMux I__635 (
            .O(N__3866),
            .I(\U400_SDRAM.N_60 ));
    CascadeMux I__634 (
            .O(N__3863),
            .I(\U400_SDRAM.N_97_cascade_ ));
    InMux I__633 (
            .O(N__3860),
            .I(N__3857));
    LocalMux I__632 (
            .O(N__3857),
            .I(N__3853));
    InMux I__631 (
            .O(N__3856),
            .I(N__3850));
    Odrv4 I__630 (
            .O(N__3853),
            .I(\U400_SDRAM.N_20 ));
    LocalMux I__629 (
            .O(N__3850),
            .I(\U400_SDRAM.N_20 ));
    CascadeMux I__628 (
            .O(N__3845),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_0_1_66_i_0_2_cascade_ ));
    CascadeMux I__627 (
            .O(N__3842),
            .I(N__3839));
    InMux I__626 (
            .O(N__3839),
            .I(N__3836));
    LocalMux I__625 (
            .O(N__3836),
            .I(N__3833));
    Span4Mux_v I__624 (
            .O(N__3833),
            .I(N__3830));
    Span4Mux_h I__623 (
            .O(N__3830),
            .I(N__3827));
    Odrv4 I__622 (
            .O(N__3827),
            .I(A_c_18));
    InMux I__621 (
            .O(N__3824),
            .I(N__3820));
    InMux I__620 (
            .O(N__3823),
            .I(N__3817));
    LocalMux I__619 (
            .O(N__3820),
            .I(N__3813));
    LocalMux I__618 (
            .O(N__3817),
            .I(N__3810));
    InMux I__617 (
            .O(N__3816),
            .I(N__3807));
    Odrv4 I__616 (
            .O(N__3813),
            .I(\U400_SDRAM.N_11 ));
    Odrv4 I__615 (
            .O(N__3810),
            .I(\U400_SDRAM.N_11 ));
    LocalMux I__614 (
            .O(N__3807),
            .I(\U400_SDRAM.N_11 ));
    InMux I__613 (
            .O(N__3800),
            .I(N__3797));
    LocalMux I__612 (
            .O(N__3797),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_1 ));
    CascadeMux I__611 (
            .O(N__3794),
            .I(\U400_SDRAM.N_44_cascade_ ));
    InMux I__610 (
            .O(N__3791),
            .I(N__3784));
    InMux I__609 (
            .O(N__3790),
            .I(N__3784));
    InMux I__608 (
            .O(N__3789),
            .I(N__3781));
    LocalMux I__607 (
            .O(N__3784),
            .I(N__3777));
    LocalMux I__606 (
            .O(N__3781),
            .I(N__3773));
    InMux I__605 (
            .O(N__3780),
            .I(N__3770));
    Span4Mux_h I__604 (
            .O(N__3777),
            .I(N__3767));
    InMux I__603 (
            .O(N__3776),
            .I(N__3764));
    Odrv4 I__602 (
            .O(N__3773),
            .I(\U400_SDRAM.N_108 ));
    LocalMux I__601 (
            .O(N__3770),
            .I(\U400_SDRAM.N_108 ));
    Odrv4 I__600 (
            .O(N__3767),
            .I(\U400_SDRAM.N_108 ));
    LocalMux I__599 (
            .O(N__3764),
            .I(\U400_SDRAM.N_108 ));
    CascadeMux I__598 (
            .O(N__3755),
            .I(\U400_SDRAM.N_108_cascade_ ));
    InMux I__597 (
            .O(N__3752),
            .I(N__3749));
    LocalMux I__596 (
            .O(N__3749),
            .I(N__3746));
    Span4Mux_h I__595 (
            .O(N__3746),
            .I(N__3742));
    InMux I__594 (
            .O(N__3745),
            .I(N__3739));
    Odrv4 I__593 (
            .O(N__3742),
            .I(\U400_SDRAM.N_109 ));
    LocalMux I__592 (
            .O(N__3739),
            .I(\U400_SDRAM.N_109 ));
    InMux I__591 (
            .O(N__3734),
            .I(N__3727));
    InMux I__590 (
            .O(N__3733),
            .I(N__3727));
    InMux I__589 (
            .O(N__3732),
            .I(N__3724));
    LocalMux I__588 (
            .O(N__3727),
            .I(N__3721));
    LocalMux I__587 (
            .O(N__3724),
            .I(\U400_SDRAM.N_52 ));
    Odrv4 I__586 (
            .O(N__3721),
            .I(\U400_SDRAM.N_52 ));
    InMux I__585 (
            .O(N__3716),
            .I(N__3713));
    LocalMux I__584 (
            .O(N__3713),
            .I(N__3710));
    Span4Mux_h I__583 (
            .O(N__3710),
            .I(N__3707));
    Span4Mux_s1_h I__582 (
            .O(N__3707),
            .I(N__3704));
    Odrv4 I__581 (
            .O(N__3704),
            .I(\U400_SDRAM.SDRAM_COUNTER_s_0 ));
    InMux I__580 (
            .O(N__3701),
            .I(N__3698));
    LocalMux I__579 (
            .O(N__3698),
            .I(N__3695));
    Odrv4 I__578 (
            .O(N__3695),
            .I(\U400_SDRAM.N_86 ));
    CascadeMux I__577 (
            .O(N__3692),
            .I(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_1_0_cascade_ ));
    InMux I__576 (
            .O(N__3689),
            .I(N__3684));
    InMux I__575 (
            .O(N__3688),
            .I(N__3681));
    InMux I__574 (
            .O(N__3687),
            .I(N__3678));
    LocalMux I__573 (
            .O(N__3684),
            .I(\U400_SDRAM.SDRAM_CMD_3_sqmuxa ));
    LocalMux I__572 (
            .O(N__3681),
            .I(\U400_SDRAM.SDRAM_CMD_3_sqmuxa ));
    LocalMux I__571 (
            .O(N__3678),
            .I(\U400_SDRAM.SDRAM_CMD_3_sqmuxa ));
    InMux I__570 (
            .O(N__3671),
            .I(N__3668));
    LocalMux I__569 (
            .O(N__3668),
            .I(N__3664));
    InMux I__568 (
            .O(N__3667),
            .I(N__3661));
    Span4Mux_v I__567 (
            .O(N__3664),
            .I(N__3656));
    LocalMux I__566 (
            .O(N__3661),
            .I(N__3656));
    Span4Mux_h I__565 (
            .O(N__3656),
            .I(N__3652));
    InMux I__564 (
            .O(N__3655),
            .I(N__3649));
    Odrv4 I__563 (
            .O(N__3652),
            .I(\U400_SDRAM.N_118 ));
    LocalMux I__562 (
            .O(N__3649),
            .I(\U400_SDRAM.N_118 ));
    InMux I__561 (
            .O(N__3644),
            .I(N__3641));
    LocalMux I__560 (
            .O(N__3641),
            .I(\U400_SDRAM.SDRAM_COUNTER_3_sqmuxa_0_a3_0_a2_0 ));
    CascadeMux I__559 (
            .O(N__3638),
            .I(\U400_SDRAM.N_46_cascade_ ));
    InMux I__558 (
            .O(N__3635),
            .I(N__3632));
    LocalMux I__557 (
            .O(N__3632),
            .I(N__3628));
    InMux I__556 (
            .O(N__3631),
            .I(N__3622));
    Span4Mux_s2_v I__555 (
            .O(N__3628),
            .I(N__3619));
    InMux I__554 (
            .O(N__3627),
            .I(N__3614));
    InMux I__553 (
            .O(N__3626),
            .I(N__3614));
    InMux I__552 (
            .O(N__3625),
            .I(N__3607));
    LocalMux I__551 (
            .O(N__3622),
            .I(N__3600));
    Span4Mux_v I__550 (
            .O(N__3619),
            .I(N__3600));
    LocalMux I__549 (
            .O(N__3614),
            .I(N__3600));
    InMux I__548 (
            .O(N__3613),
            .I(N__3591));
    InMux I__547 (
            .O(N__3612),
            .I(N__3591));
    InMux I__546 (
            .O(N__3611),
            .I(N__3591));
    InMux I__545 (
            .O(N__3610),
            .I(N__3591));
    LocalMux I__544 (
            .O(N__3607),
            .I(\U400_SDRAM.RAM_CYCLE_STARTZ0 ));
    Odrv4 I__543 (
            .O(N__3600),
            .I(\U400_SDRAM.RAM_CYCLE_STARTZ0 ));
    LocalMux I__542 (
            .O(N__3591),
            .I(\U400_SDRAM.RAM_CYCLE_STARTZ0 ));
    InMux I__541 (
            .O(N__3584),
            .I(N__3581));
    LocalMux I__540 (
            .O(N__3581),
            .I(\U400_SDRAM.SDRAM_COUNTER_4_sqmuxa_0_a3_0 ));
    InMux I__539 (
            .O(N__3578),
            .I(N__3575));
    LocalMux I__538 (
            .O(N__3575),
            .I(N__3572));
    Span4Mux_v I__537 (
            .O(N__3572),
            .I(N__3569));
    Span4Mux_h I__536 (
            .O(N__3569),
            .I(N__3566));
    Odrv4 I__535 (
            .O(N__3566),
            .I(RnW_c));
    InMux I__534 (
            .O(N__3563),
            .I(N__3560));
    LocalMux I__533 (
            .O(N__3560),
            .I(N__3554));
    InMux I__532 (
            .O(N__3559),
            .I(N__3549));
    InMux I__531 (
            .O(N__3558),
            .I(N__3549));
    InMux I__530 (
            .O(N__3557),
            .I(N__3546));
    Odrv4 I__529 (
            .O(N__3554),
            .I(\U400_SDRAM.N_113 ));
    LocalMux I__528 (
            .O(N__3549),
            .I(\U400_SDRAM.N_113 ));
    LocalMux I__527 (
            .O(N__3546),
            .I(\U400_SDRAM.N_113 ));
    InMux I__526 (
            .O(N__3539),
            .I(N__3536));
    LocalMux I__525 (
            .O(N__3536),
            .I(\U400_SDRAM.N_63 ));
    CascadeMux I__524 (
            .O(N__3533),
            .I(\U400_SDRAM.N_20_cascade_ ));
    InMux I__523 (
            .O(N__3530),
            .I(N__3527));
    LocalMux I__522 (
            .O(N__3527),
            .I(N__3524));
    Odrv12 I__521 (
            .O(N__3524),
            .I(\U400_SDRAM.N_35 ));
    InMux I__520 (
            .O(N__3521),
            .I(N__3518));
    LocalMux I__519 (
            .O(N__3518),
            .I(N__3514));
    InMux I__518 (
            .O(N__3517),
            .I(N__3511));
    Odrv12 I__517 (
            .O(N__3514),
            .I(\U400_SDRAM.N_39 ));
    LocalMux I__516 (
            .O(N__3511),
            .I(\U400_SDRAM.N_39 ));
    CascadeMux I__515 (
            .O(N__3506),
            .I(\U400_SDRAM.N_35_cascade_ ));
    CascadeMux I__514 (
            .O(N__3503),
            .I(\U400_SDRAM.N_12_cascade_ ));
    CascadeMux I__513 (
            .O(N__3500),
            .I(\U400_SDRAM.N_91_cascade_ ));
    InMux I__512 (
            .O(N__3497),
            .I(N__3494));
    LocalMux I__511 (
            .O(N__3494),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_0_0_103_i_i_a3_0_0 ));
    InMux I__510 (
            .O(N__3491),
            .I(N__3488));
    LocalMux I__509 (
            .O(N__3488),
            .I(\U400_SDRAM.N_89 ));
    CascadeMux I__508 (
            .O(N__3485),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_0_0_103_i_i_0_cascade_ ));
    InMux I__507 (
            .O(N__3482),
            .I(N__3479));
    LocalMux I__506 (
            .O(N__3479),
            .I(N__3476));
    Span4Mux_v I__505 (
            .O(N__3476),
            .I(N__3473));
    Span4Mux_h I__504 (
            .O(N__3473),
            .I(N__3470));
    Odrv4 I__503 (
            .O(N__3470),
            .I(A_c_8));
    CascadeMux I__502 (
            .O(N__3467),
            .I(N__3464));
    InMux I__501 (
            .O(N__3464),
            .I(N__3461));
    LocalMux I__500 (
            .O(N__3461),
            .I(N__3458));
    Span4Mux_v I__499 (
            .O(N__3458),
            .I(N__3455));
    Span4Mux_v I__498 (
            .O(N__3455),
            .I(N__3452));
    Odrv4 I__497 (
            .O(N__3452),
            .I(A_c_19));
    IoInMux I__496 (
            .O(N__3449),
            .I(N__3446));
    LocalMux I__495 (
            .O(N__3446),
            .I(N__3443));
    Odrv12 I__494 (
            .O(N__3443),
            .I(MA_c_6));
    InMux I__493 (
            .O(N__3440),
            .I(N__3437));
    LocalMux I__492 (
            .O(N__3437),
            .I(N__3434));
    Odrv12 I__491 (
            .O(N__3434),
            .I(A_c_6));
    CascadeMux I__490 (
            .O(N__3431),
            .I(N__3428));
    InMux I__489 (
            .O(N__3428),
            .I(N__3425));
    LocalMux I__488 (
            .O(N__3425),
            .I(N__3422));
    Span12Mux_s8_v I__487 (
            .O(N__3422),
            .I(N__3419));
    Odrv12 I__486 (
            .O(N__3419),
            .I(A_c_17));
    IoInMux I__485 (
            .O(N__3416),
            .I(N__3413));
    LocalMux I__484 (
            .O(N__3413),
            .I(N__3410));
    Span4Mux_s3_v I__483 (
            .O(N__3410),
            .I(N__3407));
    Odrv4 I__482 (
            .O(N__3407),
            .I(MA_c_4));
    InMux I__481 (
            .O(N__3404),
            .I(N__3401));
    LocalMux I__480 (
            .O(N__3401),
            .I(N__3398));
    Span4Mux_v I__479 (
            .O(N__3398),
            .I(N__3395));
    Span4Mux_v I__478 (
            .O(N__3395),
            .I(N__3392));
    Span4Mux_v I__477 (
            .O(N__3392),
            .I(N__3389));
    Odrv4 I__476 (
            .O(N__3389),
            .I(A_c_20));
    CascadeMux I__475 (
            .O(N__3386),
            .I(N__3383));
    InMux I__474 (
            .O(N__3383),
            .I(N__3380));
    LocalMux I__473 (
            .O(N__3380),
            .I(N__3377));
    Span12Mux_s4_v I__472 (
            .O(N__3377),
            .I(N__3374));
    Odrv12 I__471 (
            .O(N__3374),
            .I(A_c_9));
    IoInMux I__470 (
            .O(N__3371),
            .I(N__3368));
    LocalMux I__469 (
            .O(N__3368),
            .I(N__3365));
    Odrv12 I__468 (
            .O(N__3365),
            .I(MA_c_7));
    CascadeMux I__467 (
            .O(N__3362),
            .I(\U400_SDRAM.N_113_cascade_ ));
    CascadeMux I__466 (
            .O(N__3359),
            .I(\U400_SDRAM.N_39_cascade_ ));
    InMux I__465 (
            .O(N__3356),
            .I(N__3353));
    LocalMux I__464 (
            .O(N__3353),
            .I(N__3350));
    Odrv4 I__463 (
            .O(N__3350),
            .I(\U400_SDRAM.SDRAM_COUNTER_1_sqmuxa_i_0_1 ));
    InMux I__462 (
            .O(N__3347),
            .I(N__3344));
    LocalMux I__461 (
            .O(N__3344),
            .I(N__3341));
    Span4Mux_s2_h I__460 (
            .O(N__3341),
            .I(N__3338));
    Odrv4 I__459 (
            .O(N__3338),
            .I(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_a2_1_0_0 ));
    CascadeMux I__458 (
            .O(N__3335),
            .I(\U400_SDRAM.N_78_cascade_ ));
    InMux I__457 (
            .O(N__3332),
            .I(N__3326));
    InMux I__456 (
            .O(N__3331),
            .I(N__3326));
    LocalMux I__455 (
            .O(N__3326),
            .I(N__3321));
    CascadeMux I__454 (
            .O(N__3325),
            .I(N__3318));
    InMux I__453 (
            .O(N__3324),
            .I(N__3314));
    Span4Mux_v I__452 (
            .O(N__3321),
            .I(N__3311));
    InMux I__451 (
            .O(N__3318),
            .I(N__3306));
    InMux I__450 (
            .O(N__3317),
            .I(N__3306));
    LocalMux I__449 (
            .O(N__3314),
            .I(\U400_SDRAM.N_337_1 ));
    Odrv4 I__448 (
            .O(N__3311),
            .I(\U400_SDRAM.N_337_1 ));
    LocalMux I__447 (
            .O(N__3306),
            .I(\U400_SDRAM.N_337_1 ));
    IoInMux I__446 (
            .O(N__3299),
            .I(N__3296));
    LocalMux I__445 (
            .O(N__3296),
            .I(N__3293));
    Odrv4 I__444 (
            .O(N__3293),
            .I(RASn_c));
    CascadeMux I__443 (
            .O(N__3290),
            .I(N__3287));
    InMux I__442 (
            .O(N__3287),
            .I(N__3284));
    LocalMux I__441 (
            .O(N__3284),
            .I(N__3280));
    InMux I__440 (
            .O(N__3283),
            .I(N__3277));
    Odrv12 I__439 (
            .O(N__3280),
            .I(\U400_SDRAM.CS0_ENZ0 ));
    LocalMux I__438 (
            .O(N__3277),
            .I(\U400_SDRAM.CS0_ENZ0 ));
    IoInMux I__437 (
            .O(N__3272),
            .I(N__3269));
    LocalMux I__436 (
            .O(N__3269),
            .I(N__3266));
    Odrv4 I__435 (
            .O(N__3266),
            .I(CS0n_c));
    InMux I__434 (
            .O(N__3263),
            .I(N__3260));
    LocalMux I__433 (
            .O(N__3260),
            .I(N__3257));
    Span4Mux_h I__432 (
            .O(N__3257),
            .I(N__3254));
    Odrv4 I__431 (
            .O(N__3254),
            .I(A_c_31));
    InMux I__430 (
            .O(N__3251),
            .I(N__3248));
    LocalMux I__429 (
            .O(N__3248),
            .I(N__3245));
    Span4Mux_h I__428 (
            .O(N__3245),
            .I(N__3242));
    Odrv4 I__427 (
            .O(N__3242),
            .I(A_c_30));
    InMux I__426 (
            .O(N__3239),
            .I(N__3236));
    LocalMux I__425 (
            .O(N__3236),
            .I(N__3233));
    Span4Mux_h I__424 (
            .O(N__3233),
            .I(N__3230));
    Odrv4 I__423 (
            .O(N__3230),
            .I(A_c_29));
    InMux I__422 (
            .O(N__3227),
            .I(N__3224));
    LocalMux I__421 (
            .O(N__3224),
            .I(A_c_28));
    InMux I__420 (
            .O(N__3221),
            .I(N__3218));
    LocalMux I__419 (
            .O(N__3218),
            .I(N__3215));
    Span12Mux_s6_v I__418 (
            .O(N__3215),
            .I(N__3212));
    Odrv12 I__417 (
            .O(N__3212),
            .I(TSn_c));
    InMux I__416 (
            .O(N__3209),
            .I(N__3206));
    LocalMux I__415 (
            .O(N__3206),
            .I(N__3203));
    Span4Mux_v I__414 (
            .O(N__3203),
            .I(N__3200));
    Odrv4 I__413 (
            .O(N__3200),
            .I(\U400_SDRAM.N_101 ));
    InMux I__412 (
            .O(N__3197),
            .I(N__3193));
    InMux I__411 (
            .O(N__3196),
            .I(N__3190));
    LocalMux I__410 (
            .O(N__3193),
            .I(N__3185));
    LocalMux I__409 (
            .O(N__3190),
            .I(N__3185));
    Odrv4 I__408 (
            .O(N__3185),
            .I(U400_ADDRESS_DECODE_RAM_SPACE_i_o3_2));
    CascadeMux I__407 (
            .O(N__3182),
            .I(N__3178));
    InMux I__406 (
            .O(N__3181),
            .I(N__3173));
    InMux I__405 (
            .O(N__3178),
            .I(N__3173));
    LocalMux I__404 (
            .O(N__3173),
            .I(N__3170));
    Span12Mux_v I__403 (
            .O(N__3170),
            .I(N__3167));
    Odrv12 I__402 (
            .O(N__3167),
            .I(A_c_27));
    CascadeMux I__401 (
            .O(N__3164),
            .I(N__3161));
    InMux I__400 (
            .O(N__3161),
            .I(N__3155));
    InMux I__399 (
            .O(N__3160),
            .I(N__3155));
    LocalMux I__398 (
            .O(N__3155),
            .I(N__3152));
    Odrv4 I__397 (
            .O(N__3152),
            .I(U400_ADDRESS_DECODE_RAM_SPACE_i_o3_1));
    CascadeMux I__396 (
            .O(N__3149),
            .I(\U400_SDRAM.N_72_cascade_ ));
    InMux I__395 (
            .O(N__3146),
            .I(N__3143));
    LocalMux I__394 (
            .O(N__3143),
            .I(\U400_SDRAM.N_40 ));
    CascadeMux I__393 (
            .O(N__3140),
            .I(N__3137));
    InMux I__392 (
            .O(N__3137),
            .I(N__3131));
    InMux I__391 (
            .O(N__3136),
            .I(N__3131));
    LocalMux I__390 (
            .O(N__3131),
            .I(N__3128));
    Span4Mux_h I__389 (
            .O(N__3128),
            .I(N__3125));
    Span4Mux_v I__388 (
            .O(N__3125),
            .I(N__3122));
    Odrv4 I__387 (
            .O(N__3122),
            .I(A_c_23));
    CascadeMux I__386 (
            .O(N__3119),
            .I(\U400_SDRAM.N_40_cascade_ ));
    InMux I__385 (
            .O(N__3116),
            .I(N__3113));
    LocalMux I__384 (
            .O(N__3113),
            .I(\U400_SDRAM.CS0_EN_0 ));
    CascadeMux I__383 (
            .O(N__3110),
            .I(N__3105));
    InMux I__382 (
            .O(N__3109),
            .I(N__3102));
    InMux I__381 (
            .O(N__3108),
            .I(N__3097));
    InMux I__380 (
            .O(N__3105),
            .I(N__3097));
    LocalMux I__379 (
            .O(N__3102),
            .I(\U400_SDRAM.N_115 ));
    LocalMux I__378 (
            .O(N__3097),
            .I(\U400_SDRAM.N_115 ));
    CascadeMux I__377 (
            .O(N__3092),
            .I(N__3089));
    InMux I__376 (
            .O(N__3089),
            .I(N__3085));
    InMux I__375 (
            .O(N__3088),
            .I(N__3082));
    LocalMux I__374 (
            .O(N__3085),
            .I(\U400_SDRAM.RAM_CYCLEZ0 ));
    LocalMux I__373 (
            .O(N__3082),
            .I(\U400_SDRAM.RAM_CYCLEZ0 ));
    CascadeMux I__372 (
            .O(N__3077),
            .I(N__3074));
    InMux I__371 (
            .O(N__3074),
            .I(N__3071));
    LocalMux I__370 (
            .O(N__3071),
            .I(N__3067));
    InMux I__369 (
            .O(N__3070),
            .I(N__3064));
    Span4Mux_v I__368 (
            .O(N__3067),
            .I(N__3061));
    LocalMux I__367 (
            .O(N__3064),
            .I(N__3058));
    Odrv4 I__366 (
            .O(N__3061),
            .I(\U400_SDRAM.CS1_ENZ0 ));
    Odrv4 I__365 (
            .O(N__3058),
            .I(\U400_SDRAM.CS1_ENZ0 ));
    IoInMux I__364 (
            .O(N__3053),
            .I(N__3050));
    LocalMux I__363 (
            .O(N__3050),
            .I(N__3047));
    Span4Mux_s3_v I__362 (
            .O(N__3047),
            .I(N__3044));
    Span4Mux_v I__361 (
            .O(N__3044),
            .I(N__3041));
    Odrv4 I__360 (
            .O(N__3041),
            .I(CS1n_c));
    IoInMux I__359 (
            .O(N__3038),
            .I(N__3035));
    LocalMux I__358 (
            .O(N__3035),
            .I(N__3032));
    Odrv4 I__357 (
            .O(N__3032),
            .I(CASn_c));
    IoInMux I__356 (
            .O(N__3029),
            .I(N__3026));
    LocalMux I__355 (
            .O(N__3026),
            .I(N__3023));
    Odrv12 I__354 (
            .O(N__3023),
            .I(WEn_c));
    InMux I__353 (
            .O(N__3020),
            .I(\U400_SDRAM.un3_REFRESH_COUNTER_cry_7 ));
    SRMux I__352 (
            .O(N__3017),
            .I(N__3014));
    LocalMux I__351 (
            .O(N__3014),
            .I(N__3010));
    SRMux I__350 (
            .O(N__3013),
            .I(N__3007));
    Span4Mux_h I__349 (
            .O(N__3010),
            .I(N__3004));
    LocalMux I__348 (
            .O(N__3007),
            .I(N__3001));
    Span4Mux_s0_h I__347 (
            .O(N__3004),
            .I(N__2996));
    Span4Mux_h I__346 (
            .O(N__3001),
            .I(N__2996));
    Odrv4 I__345 (
            .O(N__2996),
            .I(\U400_SDRAM.SDRAM_COUNTER_RNIV59H2Z0Z_1 ));
    InMux I__344 (
            .O(N__2993),
            .I(N__2989));
    InMux I__343 (
            .O(N__2992),
            .I(N__2986));
    LocalMux I__342 (
            .O(N__2989),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__341 (
            .O(N__2986),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__340 (
            .O(N__2981),
            .I(N__2977));
    InMux I__339 (
            .O(N__2980),
            .I(N__2974));
    LocalMux I__338 (
            .O(N__2977),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__337 (
            .O(N__2974),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__336 (
            .O(N__2969),
            .I(N__2965));
    InMux I__335 (
            .O(N__2968),
            .I(N__2962));
    LocalMux I__334 (
            .O(N__2965),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__333 (
            .O(N__2962),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__332 (
            .O(N__2957),
            .I(N__2953));
    InMux I__331 (
            .O(N__2956),
            .I(N__2950));
    LocalMux I__330 (
            .O(N__2953),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__329 (
            .O(N__2950),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__328 (
            .O(N__2945),
            .I(N__2941));
    InMux I__327 (
            .O(N__2944),
            .I(N__2938));
    LocalMux I__326 (
            .O(N__2941),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_8 ));
    LocalMux I__325 (
            .O(N__2938),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_8 ));
    CascadeMux I__324 (
            .O(N__2933),
            .I(\U400_SDRAM.un1_REFRESH_COUNTERlt7_0_cascade_ ));
    InMux I__323 (
            .O(N__2930),
            .I(N__2926));
    InMux I__322 (
            .O(N__2929),
            .I(N__2923));
    LocalMux I__321 (
            .O(N__2926),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_7 ));
    LocalMux I__320 (
            .O(N__2923),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_7 ));
    CascadeMux I__319 (
            .O(N__2918),
            .I(\U400_SDRAM.N_337_1_cascade_ ));
    CascadeMux I__318 (
            .O(N__2915),
            .I(\U400_SDRAM.N_64_cascade_ ));
    InMux I__317 (
            .O(N__2912),
            .I(N__2909));
    LocalMux I__316 (
            .O(N__2909),
            .I(\U400_SDRAM.CS1_EN_0 ));
    InMux I__315 (
            .O(N__2906),
            .I(N__2901));
    InMux I__314 (
            .O(N__2905),
            .I(N__2898));
    InMux I__313 (
            .O(N__2904),
            .I(N__2895));
    LocalMux I__312 (
            .O(N__2901),
            .I(N__2892));
    LocalMux I__311 (
            .O(N__2898),
            .I(\U400_SDRAM.N_64 ));
    LocalMux I__310 (
            .O(N__2895),
            .I(\U400_SDRAM.N_64 ));
    Odrv4 I__309 (
            .O(N__2892),
            .I(\U400_SDRAM.N_64 ));
    IoInMux I__308 (
            .O(N__2885),
            .I(N__2882));
    LocalMux I__307 (
            .O(N__2882),
            .I(RESETn_c_i));
    InMux I__306 (
            .O(N__2879),
            .I(N__2875));
    InMux I__305 (
            .O(N__2878),
            .I(N__2872));
    LocalMux I__304 (
            .O(N__2875),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_1 ));
    LocalMux I__303 (
            .O(N__2872),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_1 ));
    CascadeMux I__302 (
            .O(N__2867),
            .I(N__2862));
    InMux I__301 (
            .O(N__2866),
            .I(N__2857));
    InMux I__300 (
            .O(N__2865),
            .I(N__2857));
    InMux I__299 (
            .O(N__2862),
            .I(N__2854));
    LocalMux I__298 (
            .O(N__2857),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_0 ));
    LocalMux I__297 (
            .O(N__2854),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_0 ));
    InMux I__296 (
            .O(N__2849),
            .I(N__2846));
    LocalMux I__295 (
            .O(N__2846),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_2 ));
    InMux I__294 (
            .O(N__2843),
            .I(\U400_SDRAM.un3_REFRESH_COUNTER_cry_1 ));
    InMux I__293 (
            .O(N__2840),
            .I(\U400_SDRAM.un3_REFRESH_COUNTER_cry_2 ));
    InMux I__292 (
            .O(N__2837),
            .I(\U400_SDRAM.un3_REFRESH_COUNTER_cry_3 ));
    InMux I__291 (
            .O(N__2834),
            .I(\U400_SDRAM.un3_REFRESH_COUNTER_cry_4 ));
    InMux I__290 (
            .O(N__2831),
            .I(\U400_SDRAM.un3_REFRESH_COUNTER_cry_5 ));
    InMux I__289 (
            .O(N__2828),
            .I(\U400_SDRAM.un3_REFRESH_COUNTER_cry_6 ));
    CascadeMux I__288 (
            .O(N__2825),
            .I(N__2822));
    InMux I__287 (
            .O(N__2822),
            .I(N__2819));
    LocalMux I__286 (
            .O(N__2819),
            .I(A_c_21));
    IoInMux I__285 (
            .O(N__2816),
            .I(N__2813));
    LocalMux I__284 (
            .O(N__2813),
            .I(N__2810));
    IoSpan4Mux I__283 (
            .O(N__2810),
            .I(N__2807));
    Span4Mux_s0_h I__282 (
            .O(N__2807),
            .I(N__2804));
    Span4Mux_v I__281 (
            .O(N__2804),
            .I(N__2800));
    InMux I__280 (
            .O(N__2803),
            .I(N__2797));
    Odrv4 I__279 (
            .O(N__2800),
            .I(BANK0_c));
    LocalMux I__278 (
            .O(N__2797),
            .I(BANK0_c));
    IoInMux I__277 (
            .O(N__2792),
            .I(N__2789));
    LocalMux I__276 (
            .O(N__2789),
            .I(N__2786));
    Span4Mux_s0_h I__275 (
            .O(N__2786),
            .I(N__2783));
    Span4Mux_v I__274 (
            .O(N__2783),
            .I(N__2779));
    InMux I__273 (
            .O(N__2782),
            .I(N__2776));
    Span4Mux_v I__272 (
            .O(N__2779),
            .I(N__2771));
    LocalMux I__271 (
            .O(N__2776),
            .I(N__2771));
    Odrv4 I__270 (
            .O(N__2771),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__269 (
            .O(N__2768),
            .I(N__2765));
    InMux I__268 (
            .O(N__2765),
            .I(N__2762));
    LocalMux I__267 (
            .O(N__2762),
            .I(N__2759));
    Span12Mux_s2_h I__266 (
            .O(N__2759),
            .I(N__2756));
    Odrv12 I__265 (
            .O(N__2756),
            .I(A_c_22));
    IoInMux I__264 (
            .O(N__2753),
            .I(N__2750));
    LocalMux I__263 (
            .O(N__2750),
            .I(N__2747));
    IoSpan4Mux I__262 (
            .O(N__2747),
            .I(N__2744));
    IoSpan4Mux I__261 (
            .O(N__2744),
            .I(N__2740));
    InMux I__260 (
            .O(N__2743),
            .I(N__2737));
    Odrv4 I__259 (
            .O(N__2740),
            .I(BANK1_c));
    LocalMux I__258 (
            .O(N__2737),
            .I(BANK1_c));
    InMux I__257 (
            .O(N__2732),
            .I(N__2726));
    InMux I__256 (
            .O(N__2731),
            .I(N__2726));
    LocalMux I__255 (
            .O(N__2726),
            .I(\U400_SDRAM.un1_SDRAM_COUNTER59_0 ));
    InMux I__254 (
            .O(N__2723),
            .I(N__2720));
    LocalMux I__253 (
            .O(N__2720),
            .I(\U400_SDRAM.SDRAM_CMD_5_sqmuxa ));
    IoInMux I__252 (
            .O(N__2717),
            .I(N__2714));
    LocalMux I__251 (
            .O(N__2714),
            .I(N__2711));
    IoSpan4Mux I__250 (
            .O(N__2711),
            .I(N__2708));
    IoSpan4Mux I__249 (
            .O(N__2708),
            .I(N__2705));
    Span4Mux_s2_h I__248 (
            .O(N__2705),
            .I(N__2702));
    Sp12to4 I__247 (
            .O(N__2702),
            .I(N__2699));
    Odrv12 I__246 (
            .O(N__2699),
            .I(CLK40_ibuf_gb_io_gb_input));
    INV \INVU400_SDRAM.MA_nesr_1C  (
            .O(\INVU400_SDRAM.MA_nesr_1C_net ),
            .I(N__5498));
    INV \INVU400_SDRAM.MA_nesr_10C  (
            .O(\INVU400_SDRAM.MA_nesr_10C_net ),
            .I(N__5497));
    INV \INVU400_SDRAM.BURSTC  (
            .O(\INVU400_SDRAM.BURSTC_net ),
            .I(N__5493));
    INV \INVU400_SDRAM.MA_nesr_11C  (
            .O(\INVU400_SDRAM.MA_nesr_11C_net ),
            .I(N__5496));
    INV \INVU400_SDRAM.SDRAM_COUNTER_2C  (
            .O(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .I(N__5490));
    INV \INVU400_SDRAM.MA_nesr_3C  (
            .O(\INVU400_SDRAM.MA_nesr_3C_net ),
            .I(N__5489));
    INV \INVU400_SDRAM.SDRAM_CMD_0C  (
            .O(\INVU400_SDRAM.SDRAM_CMD_0C_net ),
            .I(N__5483));
    INV \INVU400_SDRAM.SDRAM_COUNTER_0C  (
            .O(\INVU400_SDRAM.SDRAM_COUNTER_0C_net ),
            .I(N__5487));
    INV \INVU400_SDRAM.TACKC  (
            .O(\INVU400_SDRAM.TACKC_net ),
            .I(N__5491));
    INV \INVU400_SDRAM.MA_nesr_6C  (
            .O(\INVU400_SDRAM.MA_nesr_6C_net ),
            .I(N__5485));
    INV \INVU400_SDRAM.SDRAM_CMD_1C  (
            .O(\INVU400_SDRAM.SDRAM_CMD_1C_net ),
            .I(N__5480));
    INV \INVU400_SDRAM.SDRAM_CONFIGUREDC  (
            .O(\INVU400_SDRAM.SDRAM_CONFIGUREDC_net ),
            .I(N__5486));
    INV \INVU400_SDRAM.SDRAM_COUNTER_1C  (
            .O(\INVU400_SDRAM.SDRAM_COUNTER_1C_net ),
            .I(N__5488));
    INV \INVU400_SDRAM.RASnC  (
            .O(\INVU400_SDRAM.RASnC_net ),
            .I(N__5476));
    INV \INVU400_SDRAM.CS1nC  (
            .O(\INVU400_SDRAM.CS1nC_net ),
            .I(N__5474));
    INV \INVU400_SDRAM.CS0_ENC  (
            .O(\INVU400_SDRAM.CS0_ENC_net ),
            .I(N__5482));
    INV \INVU400_SDRAM.REFRESH_COUNTER_2C  (
            .O(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .I(N__5484));
    INV \INVU400_SDRAM.RAM_CYCLEC  (
            .O(\INVU400_SDRAM.RAM_CYCLEC_net ),
            .I(N__5475));
    INV \INVU400_SDRAM.CS1_ENC  (
            .O(\INVU400_SDRAM.CS1_ENC_net ),
            .I(N__5477));
    INV \INVU400_SDRAM.BANK0C  (
            .O(\INVU400_SDRAM.BANK0C_net ),
            .I(N__5479));
    INV \INVU400_SDRAM.REFRESH_COUNTER_1C  (
            .O(\INVU400_SDRAM.REFRESH_COUNTER_1C_net ),
            .I(N__5481));
    defparam IN_MUX_bfv_2_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_4_0_));
    defparam IN_MUX_bfv_6_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_6_0_));
    ICE_GB CLK40_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__2717),
            .GLOBALBUFFEROUTPUT(CLK40_c_g));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__2885),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_1_3_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_1_3_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_1_3_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_1_3_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_1_LC_1_4_0 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_1_LC_1_4_0 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_1_LC_1_4_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_1_LC_1_4_0  (
            .in0(N__2866),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2879),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_1C_net ),
            .ce(),
            .sr(N__3013));
    defparam \U400_SDRAM.REFRESH_COUNTER_0_LC_1_4_1 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_0_LC_1_4_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_0_LC_1_4_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_0_LC_1_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2865),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_1C_net ),
            .ce(),
            .sr(N__3013));
    defparam \U400_SDRAM.BANK0_LC_1_5_0 .C_ON=1'b0;
    defparam \U400_SDRAM.BANK0_LC_1_5_0 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.BANK0_LC_1_5_0 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \U400_SDRAM.BANK0_LC_1_5_0  (
            .in0(N__2803),
            .in1(N__5082),
            .in2(N__2825),
            .in3(N__2731),
            .lcout(BANK0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.BANK0C_net ),
            .ce(),
            .sr(N__6348));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_2_0_LC_1_5_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_2_0_LC_1_5_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_2_0_LC_1_5_2 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_2_0_LC_1_5_2  (
            .in0(N__2782),
            .in1(N__5081),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.BANK1_LC_1_5_5 .C_ON=1'b0;
    defparam \U400_SDRAM.BANK1_LC_1_5_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.BANK1_LC_1_5_5 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \U400_SDRAM.BANK1_LC_1_5_5  (
            .in0(N__2732),
            .in1(N__2743),
            .in2(N__2768),
            .in3(N__5083),
            .lcout(BANK1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.BANK0C_net ),
            .ce(),
            .sr(N__6348));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIV59H2_1_LC_1_5_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIV59H2_1_LC_1_5_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIV59H2_1_LC_1_5_7 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIV59H2_1_LC_1_5_7  (
            .in0(N__5337),
            .in1(N__3530),
            .in2(_gnd_net_),
            .in3(N__4655),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_RNIV59H2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.CS1_EN_LC_1_6_1 .C_ON=1'b0;
    defparam \U400_SDRAM.CS1_EN_LC_1_6_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.CS1_EN_LC_1_6_1 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \U400_SDRAM.CS1_EN_LC_1_6_1  (
            .in0(N__3108),
            .in1(N__2905),
            .in2(_gnd_net_),
            .in3(N__2912),
            .lcout(\U400_SDRAM.CS1_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS1_ENC_net ),
            .ce(),
            .sr(N__6345));
    defparam \U400_SDRAM.RAM_CYCLE_RNO_0_LC_1_6_3 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_0_LC_1_6_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_0_LC_1_6_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_RNO_0_LC_1_6_3  (
            .in0(N__4406),
            .in1(N__3324),
            .in2(N__3110),
            .in3(N__3625),
            .lcout(\U400_SDRAM.SDRAM_CMD_5_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.WRITE_CYCLE_RNIF1VQ5_LC_1_6_7 .C_ON=1'b0;
    defparam \U400_SDRAM.WRITE_CYCLE_RNIF1VQ5_LC_1_6_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.WRITE_CYCLE_RNIF1VQ5_LC_1_6_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U400_SDRAM.WRITE_CYCLE_RNIF1VQ5_LC_1_6_7  (
            .in0(_gnd_net_),
            .in1(N__3521),
            .in2(_gnd_net_),
            .in3(N__5405),
            .lcout(\U400_SDRAM.un1_SDRAM_COUNTER59_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_LC_1_7_2 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_LC_1_7_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.RAM_CYCLE_LC_1_7_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_LC_1_7_2  (
            .in0(N__4826),
            .in1(N__5406),
            .in2(N__3092),
            .in3(N__2723),
            .lcout(\U400_SDRAM.RAM_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.RAM_CYCLEC_net ),
            .ce(),
            .sr(N__6344));
    defparam RESETn_ibuf_RNIM9SF_LC_1_8_3.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_1_8_3.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_1_8_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_1_8_3 (
            .in0(N__5347),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.un3_REFRESH_COUNTER_cry_1_c_LC_2_4_0 .C_ON=1'b1;
    defparam \U400_SDRAM.un3_REFRESH_COUNTER_cry_1_c_LC_2_4_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.un3_REFRESH_COUNTER_cry_1_c_LC_2_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U400_SDRAM.un3_REFRESH_COUNTER_cry_1_c_LC_2_4_0  (
            .in0(_gnd_net_),
            .in1(N__2878),
            .in2(N__2867),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_4_0_),
            .carryout(\U400_SDRAM.un3_REFRESH_COUNTER_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_2_LC_2_4_1 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_2_LC_2_4_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_2_LC_2_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_2_LC_2_4_1  (
            .in0(_gnd_net_),
            .in1(N__2849),
            .in2(_gnd_net_),
            .in3(N__2843),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U400_SDRAM.un3_REFRESH_COUNTER_cry_1 ),
            .carryout(\U400_SDRAM.un3_REFRESH_COUNTER_cry_2 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3017));
    defparam \U400_SDRAM.REFRESH_COUNTER_3_LC_2_4_2 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_3_LC_2_4_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_3_LC_2_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_3_LC_2_4_2  (
            .in0(_gnd_net_),
            .in1(N__2993),
            .in2(_gnd_net_),
            .in3(N__2840),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U400_SDRAM.un3_REFRESH_COUNTER_cry_2 ),
            .carryout(\U400_SDRAM.un3_REFRESH_COUNTER_cry_3 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3017));
    defparam \U400_SDRAM.REFRESH_COUNTER_4_LC_2_4_3 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_4_LC_2_4_3 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_4_LC_2_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_4_LC_2_4_3  (
            .in0(_gnd_net_),
            .in1(N__2969),
            .in2(_gnd_net_),
            .in3(N__2837),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U400_SDRAM.un3_REFRESH_COUNTER_cry_3 ),
            .carryout(\U400_SDRAM.un3_REFRESH_COUNTER_cry_4 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3017));
    defparam \U400_SDRAM.REFRESH_COUNTER_5_LC_2_4_4 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_5_LC_2_4_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_5_LC_2_4_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_5_LC_2_4_4  (
            .in0(_gnd_net_),
            .in1(N__2981),
            .in2(_gnd_net_),
            .in3(N__2834),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U400_SDRAM.un3_REFRESH_COUNTER_cry_4 ),
            .carryout(\U400_SDRAM.un3_REFRESH_COUNTER_cry_5 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3017));
    defparam \U400_SDRAM.REFRESH_COUNTER_6_LC_2_4_5 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_6_LC_2_4_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_6_LC_2_4_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_6_LC_2_4_5  (
            .in0(_gnd_net_),
            .in1(N__2957),
            .in2(_gnd_net_),
            .in3(N__2831),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U400_SDRAM.un3_REFRESH_COUNTER_cry_5 ),
            .carryout(\U400_SDRAM.un3_REFRESH_COUNTER_cry_6 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3017));
    defparam \U400_SDRAM.REFRESH_COUNTER_7_LC_2_4_6 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_7_LC_2_4_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_7_LC_2_4_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_7_LC_2_4_6  (
            .in0(_gnd_net_),
            .in1(N__2930),
            .in2(_gnd_net_),
            .in3(N__2828),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(\U400_SDRAM.un3_REFRESH_COUNTER_cry_6 ),
            .carryout(\U400_SDRAM.un3_REFRESH_COUNTER_cry_7 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3017));
    defparam \U400_SDRAM.REFRESH_COUNTER_8_LC_2_4_7 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_8_LC_2_4_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_8_LC_2_4_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_8_LC_2_4_7  (
            .in0(_gnd_net_),
            .in1(N__2945),
            .in2(_gnd_net_),
            .in3(N__3020),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3017));
    defparam \U400_SDRAM.CS0_EN_LC_2_5_1 .C_ON=1'b0;
    defparam \U400_SDRAM.CS0_EN_LC_2_5_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.CS0_EN_LC_2_5_1 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \U400_SDRAM.CS0_EN_LC_2_5_1  (
            .in0(N__3109),
            .in1(N__2904),
            .in2(_gnd_net_),
            .in3(N__3116),
            .lcout(\U400_SDRAM.CS0_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS0_ENC_net ),
            .ce(),
            .sr(N__6350));
    defparam \U400_SDRAM.REFRESH_COUNTER_RNILA301_3_LC_2_5_2 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNILA301_3_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNILA301_3_LC_2_5_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_RNILA301_3_LC_2_5_2  (
            .in0(N__2992),
            .in1(N__2980),
            .in2(_gnd_net_),
            .in3(N__2968),
            .lcout(),
            .ltout(\U400_SDRAM.un1_REFRESH_COUNTERlt7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIJU602_8_LC_2_5_3 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIJU602_8_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIJU602_8_LC_2_5_3 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_RNIJU602_8_LC_2_5_3  (
            .in0(N__2956),
            .in1(N__2944),
            .in2(N__2933),
            .in3(N__2929),
            .lcout(\U400_SDRAM.N_337_1 ),
            .ltout(\U400_SDRAM.N_337_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIS9I32_LC_2_5_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIS9I32_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIS9I32_LC_2_5_4 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNIS9I32_LC_2_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2918),
            .in3(N__4388),
            .lcout(\U400_SDRAM.N_64 ),
            .ltout(\U400_SDRAM.N_64_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI6JJA4_1_LC_2_5_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI6JJA4_1_LC_2_5_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI6JJA4_1_LC_2_5_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI6JJA4_1_LC_2_5_5  (
            .in0(N__5346),
            .in1(N__3789),
            .in2(N__2915),
            .in3(N__4654),
            .lcout(\U400_SDRAM.N_118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.CS1_EN_RNO_0_LC_2_6_0 .C_ON=1'b0;
    defparam \U400_SDRAM.CS1_EN_RNO_0_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.CS1_EN_RNO_0_LC_2_6_0 .LUT_INIT=16'b0000001110101010;
    LogicCell40 \U400_SDRAM.CS1_EN_RNO_0_LC_2_6_0  (
            .in0(N__3070),
            .in1(N__3734),
            .in2(N__3140),
            .in3(N__3146),
            .lcout(\U400_SDRAM.CS1_EN_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIP6F34_LC_2_6_1 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIP6F34_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIP6F34_LC_2_6_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_RNIP6F34_LC_2_6_1  (
            .in0(N__4405),
            .in1(N__3752),
            .in2(N__3325),
            .in3(N__3611),
            .lcout(\U400_SDRAM.SDRAM_CMD_1_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_0_LC_2_6_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_0_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_0_LC_2_6_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_0_0_LC_2_6_2  (
            .in0(N__3612),
            .in1(N__3347),
            .in2(_gnd_net_),
            .in3(N__2906),
            .lcout(\U400_SDRAM.N_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_RNI8DRF2_LC_2_6_3 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNI8DRF2_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNI8DRF2_LC_2_6_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_RNI8DRF2_LC_2_6_3  (
            .in0(N__3317),
            .in1(N__4645),
            .in2(_gnd_net_),
            .in3(N__3610),
            .lcout(),
            .ltout(\U400_SDRAM.N_72_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNI9NVF9_LC_2_6_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNI9NVF9_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNI9NVF9_LC_2_6_4 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNI9NVF9_LC_2_6_4  (
            .in0(N__3356),
            .in1(N__3791),
            .in2(N__3149),
            .in3(N__4404),
            .lcout(\U400_SDRAM.N_40 ),
            .ltout(\U400_SDRAM.N_40_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.CS0_EN_RNO_0_LC_2_6_5 .C_ON=1'b0;
    defparam \U400_SDRAM.CS0_EN_RNO_0_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.CS0_EN_RNO_0_LC_2_6_5 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \U400_SDRAM.CS0_EN_RNO_0_LC_2_6_5  (
            .in0(N__3733),
            .in1(N__3136),
            .in2(N__3119),
            .in3(N__3283),
            .lcout(\U400_SDRAM.CS0_EN_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIA9172_1_LC_2_6_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIA9172_1_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIA9172_1_LC_2_6_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIA9172_1_LC_2_6_6  (
            .in0(N__4646),
            .in1(N__5348),
            .in2(_gnd_net_),
            .in3(N__3790),
            .lcout(\U400_SDRAM.N_115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIFGBJ4_LC_2_6_7 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIFGBJ4_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIFGBJ4_LC_2_6_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_RNIFGBJ4_LC_2_6_7  (
            .in0(N__3655),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3613),
            .lcout(\U400_SDRAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_LC_2_7_6 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_LC_2_7_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.RAM_CYCLE_START_LC_2_7_6 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_LC_2_7_6  (
            .in0(N__3209),
            .in1(N__3088),
            .in2(_gnd_net_),
            .in3(N__3631),
            .lcout(\U400_SDRAM.RAM_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5478),
            .ce(),
            .sr(N__6346));
    defparam \U400_SDRAM.CS1n_LC_2_9_0 .C_ON=1'b0;
    defparam \U400_SDRAM.CS1n_LC_2_9_0 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.CS1n_LC_2_9_0 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \U400_SDRAM.CS1n_LC_2_9_0  (
            .in0(N__6593),
            .in1(N__5872),
            .in2(N__3077),
            .in3(N__5753),
            .lcout(CS1n_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS1nC_net ),
            .ce(),
            .sr(N__6347));
    defparam \U400_SDRAM.CASn_LC_2_9_4 .C_ON=1'b0;
    defparam \U400_SDRAM.CASn_LC_2_9_4 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.CASn_LC_2_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U400_SDRAM.CASn_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5873),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS1nC_net ),
            .ce(),
            .sr(N__6347));
    defparam \U400_SDRAM.WEn_LC_2_9_5 .C_ON=1'b0;
    defparam \U400_SDRAM.WEn_LC_2_9_5 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.WEn_LC_2_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U400_SDRAM.WEn_LC_2_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5751),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS1nC_net ),
            .ce(),
            .sr(N__6347));
    defparam \U400_SDRAM.RASn_LC_2_10_1 .C_ON=1'b0;
    defparam \U400_SDRAM.RASn_LC_2_10_1 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.RASn_LC_2_10_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U400_SDRAM.RASn_LC_2_10_1  (
            .in0(N__6595),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.RASnC_net ),
            .ce(),
            .sr(N__6349));
    defparam \U400_SDRAM.CS0n_LC_2_10_5 .C_ON=1'b0;
    defparam \U400_SDRAM.CS0n_LC_2_10_5 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.CS0n_LC_2_10_5 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \U400_SDRAM.CS0n_LC_2_10_5  (
            .in0(N__6594),
            .in1(N__5874),
            .in2(N__3290),
            .in3(N__5752),
            .lcout(CS0n_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.RASnC_net ),
            .ce(),
            .sr(N__6349));
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_2_LC_4_1_0 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_2_LC_4_1_0 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_2_LC_4_1_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_2_LC_4_1_0  (
            .in0(_gnd_net_),
            .in1(N__3263),
            .in2(_gnd_net_),
            .in3(N__3251),
            .lcout(U400_ADDRESS_DECODE_RAM_SPACE_i_o3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_1_LC_4_1_2 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_1_LC_4_1_2 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_1_LC_4_1_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_1_LC_4_1_2  (
            .in0(N__3239),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3227),
            .lcout(U400_ADDRESS_DECODE_RAM_SPACE_i_o3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_RNO_0_LC_4_3_4 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNO_0_LC_4_3_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNO_0_LC_4_3_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_RNO_0_LC_4_3_4  (
            .in0(N__3197),
            .in1(N__3181),
            .in2(N__3164),
            .in3(N__3221),
            .lcout(\U400_SDRAM.N_101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_i_o3dup_LC_4_3_7 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_i_o3dup_LC_4_3_7 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_i_o3dup_LC_4_3_7 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \U400_ADDRESS_DECODE.RAM_SPACE_i_o3dup_LC_4_3_7  (
            .in0(N__3196),
            .in1(N__5336),
            .in2(N__3182),
            .in3(N__3160),
            .lcout(RAM_SPACE_i_o3dup),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_1_LC_4_4_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_1_LC_4_4_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_1_LC_4_4_7 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_1_LC_4_4_7  (
            .in0(N__3584),
            .in1(N__4204),
            .in2(N__4034),
            .in3(N__3667),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_1C_net ),
            .ce(N__4151),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_LC_4_5_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_LC_4_5_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_LC_4_5_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_LC_4_5_5  (
            .in0(_gnd_net_),
            .in1(N__4378),
            .in2(_gnd_net_),
            .in3(N__3689),
            .lcout(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_CONFIGUREDC_net ),
            .ce(),
            .sr(N__6351));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIQQB91_0_LC_4_6_0 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIQQB91_0_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIQQB91_0_LC_4_6_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIQQB91_0_LC_4_6_0  (
            .in0(N__4741),
            .in1(N__5049),
            .in2(_gnd_net_),
            .in3(N__4889),
            .lcout(\U400_SDRAM.N_113 ),
            .ltout(\U400_SDRAM.N_113_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.WRITE_CYCLE_RNIMQFN1_LC_4_6_1 .C_ON=1'b0;
    defparam \U400_SDRAM.WRITE_CYCLE_RNIMQFN1_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.WRITE_CYCLE_RNIMQFN1_LC_4_6_1 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \U400_SDRAM.WRITE_CYCLE_RNIMQFN1_LC_4_6_1  (
            .in0(N__4968),
            .in1(N__4600),
            .in2(N__3362),
            .in3(N__4347),
            .lcout(\U400_SDRAM.N_39 ),
            .ltout(\U400_SDRAM.N_39_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIGGGC5_LC_4_6_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIGGGC5_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIGGGC5_LC_4_6_2 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNIGGGC5_LC_4_6_2  (
            .in0(N__4348),
            .in1(N__3745),
            .in2(N__3359),
            .in3(N__3687),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_1_sqmuxa_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_3_0_LC_4_6_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_3_0_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_3_0_LC_4_6_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_3_0_LC_4_6_3  (
            .in0(N__6190),
            .in1(N__3780),
            .in2(N__6119),
            .in3(N__4601),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_a2_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNINU7A_3_LC_4_6_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNINU7A_3_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNINU7A_3_LC_4_6_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNINU7A_3_LC_4_6_6  (
            .in0(N__4346),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4471),
            .lcout(\U400_SDRAM.N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI6C8G1_1_LC_4_6_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI6C8G1_1_LC_4_6_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI6C8G1_1_LC_4_6_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI6C8G1_1_LC_4_6_7  (
            .in0(_gnd_net_),
            .in1(N__3557),
            .in2(_gnd_net_),
            .in3(N__4602),
            .lcout(\U400_SDRAM.N_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_5_2_LC_4_7_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_5_2_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_5_2_LC_4_7_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_5_2_LC_4_7_1  (
            .in0(_gnd_net_),
            .in1(N__4475),
            .in2(_gnd_net_),
            .in3(N__4603),
            .lcout(\U400_SDRAM.N_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_1_LC_4_7_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_1_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_1_LC_4_7_3 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_2_1_LC_4_7_3  (
            .in0(N__3332),
            .in1(N__4604),
            .in2(_gnd_net_),
            .in3(N__5066),
            .lcout(),
            .ltout(\U400_SDRAM.N_78_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_1_LC_4_7_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_1_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_1_LC_4_7_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_0_1_LC_4_7_4  (
            .in0(N__5309),
            .in1(N__4751),
            .in2(N__3335),
            .in3(N__4384),
            .lcout(\U400_SDRAM.N_89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_RNI2IKT2_LC_4_7_5 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNI2IKT2_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNI2IKT2_LC_4_7_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_RNI2IKT2_LC_4_7_5  (
            .in0(N__3331),
            .in1(N__5067),
            .in2(N__4813),
            .in3(N__3626),
            .lcout(),
            .ltout(\U400_SDRAM.N_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI4LJ09_1_LC_4_7_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI4LJ09_1_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI4LJ09_1_LC_4_7_6 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI4LJ09_1_LC_4_7_6  (
            .in0(N__4605),
            .in1(N__3878),
            .in2(N__3503),
            .in3(N__4916),
            .lcout(\U400_SDRAM.N_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_4_7_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_4_7_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_4_7_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_4_7_7  (
            .in0(N__6114),
            .in1(N__6170),
            .in2(_gnd_net_),
            .in3(N__3627),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_3_sqmuxa_0_a3_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_4_1_LC_4_8_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_4_1_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_4_1_LC_4_8_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_4_1_LC_4_8_2  (
            .in0(N__4120),
            .in1(N__4508),
            .in2(_gnd_net_),
            .in3(N__4641),
            .lcout(\U400_SDRAM.SDRAM_CMD_cnst_0_0_103_i_i_a3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_3_1_LC_4_8_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_3_1_LC_4_8_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_3_1_LC_4_8_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_3_1_LC_4_8_5  (
            .in0(N__4642),
            .in1(N__3563),
            .in2(N__5308),
            .in3(N__3823),
            .lcout(),
            .ltout(\U400_SDRAM.N_91_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_1_LC_4_8_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_1_LC_4_8_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_1_LC_4_8_6 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_1_1_LC_4_8_6  (
            .in0(N__4919),
            .in1(N__5273),
            .in2(N__3500),
            .in3(N__3497),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_cnst_0_0_103_i_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_1_LC_4_8_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_1_LC_4_8_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_CMD_1_LC_4_8_7 .LUT_INIT=16'b0000010111001100;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_1_LC_4_8_7  (
            .in0(N__3491),
            .in1(N__5831),
            .in2(N__3485),
            .in3(N__4014),
            .lcout(\U400_SDRAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_CMD_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_6_LC_4_13_0 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_6_LC_4_13_0 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_6_LC_4_13_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \U400_SDRAM.MA_nesr_6_LC_4_13_0  (
            .in0(N__3482),
            .in1(N__6591),
            .in2(N__3467),
            .in3(N__6461),
            .lcout(MA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_6C_net ),
            .ce(N__6421),
            .sr(N__6352));
    defparam \U400_SDRAM.MA_nesr_4_LC_4_13_4 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_4_LC_4_13_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_4_LC_4_13_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \U400_SDRAM.MA_nesr_4_LC_4_13_4  (
            .in0(N__3440),
            .in1(N__6590),
            .in2(N__3431),
            .in3(N__6460),
            .lcout(MA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_6C_net ),
            .ce(N__6421),
            .sr(N__6352));
    defparam \U400_SDRAM.MA_nesr_7_LC_4_13_7 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_7_LC_4_13_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_7_LC_4_13_7 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \U400_SDRAM.MA_nesr_7_LC_4_13_7  (
            .in0(N__6462),
            .in1(N__3404),
            .in2(N__3386),
            .in3(N__6592),
            .lcout(MA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_6C_net ),
            .ce(N__6421),
            .sr(N__6352));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_5_3_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_5_3_1 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_5_3_1  (
            .in0(N__6118),
            .in1(N__6191),
            .in2(_gnd_net_),
            .in3(N__3635),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_4_sqmuxa_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_LC_5_4_4 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_LC_5_4_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TACK_LC_5_4_4 .LUT_INIT=16'b1100110011111010;
    LogicCell40 \U400_SDRAM.TACK_LC_5_4_4  (
            .in0(N__3539),
            .in1(N__5174),
            .in2(N__4106),
            .in3(N__4070),
            .lcout(\U400_SDRAM.TACKZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.TACKC_net ),
            .ce(),
            .sr(N__6353));
    defparam \U400_SDRAM.WRITE_CYCLE_RNIJKOA_LC_5_4_6 .C_ON=1'b0;
    defparam \U400_SDRAM.WRITE_CYCLE_RNIJKOA_LC_5_4_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.WRITE_CYCLE_RNIJKOA_LC_5_4_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U400_SDRAM.WRITE_CYCLE_RNIJKOA_LC_5_4_6  (
            .in0(_gnd_net_),
            .in1(N__4956),
            .in2(_gnd_net_),
            .in3(N__4577),
            .lcout(\U400_SDRAM.N_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.WRITE_CYCLE_LC_5_4_7 .C_ON=1'b0;
    defparam \U400_SDRAM.WRITE_CYCLE_LC_5_4_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.WRITE_CYCLE_LC_5_4_7 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \U400_SDRAM.WRITE_CYCLE_LC_5_4_7  (
            .in0(N__4957),
            .in1(N__3578),
            .in2(_gnd_net_),
            .in3(N__5417),
            .lcout(\U400_SDRAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.TACKC_net ),
            .ce(),
            .sr(N__6353));
    defparam \U400_SDRAM.RAM_CYCLE_RNO_2_LC_5_5_0 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_2_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_2_LC_5_5_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_RNO_2_LC_5_5_0  (
            .in0(N__4468),
            .in1(N__3558),
            .in2(N__4777),
            .in3(N__4345),
            .lcout(\U400_SDRAM.N_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_1_LC_5_5_1 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_1_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_1_LC_5_5_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U400_SDRAM.TACK_RNO_1_LC_5_5_1  (
            .in0(N__3559),
            .in1(N__4773),
            .in2(_gnd_net_),
            .in3(N__4469),
            .lcout(\U400_SDRAM.N_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNILS7A_LC_5_5_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNILS7A_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNILS7A_LC_5_5_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNILS7A_LC_5_5_2  (
            .in0(N__4552),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4344),
            .lcout(\U400_SDRAM.N_20 ),
            .ltout(\U400_SDRAM.N_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNITAGQ1_LC_5_5_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNITAGQ1_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNITAGQ1_LC_5_5_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNITAGQ1_LC_5_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3533),
            .in3(N__3776),
            .lcout(\U400_SDRAM.N_35 ),
            .ltout(\U400_SDRAM.N_35_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.WRITE_CYCLE_RNI6QCS5_LC_5_5_4 .C_ON=1'b0;
    defparam \U400_SDRAM.WRITE_CYCLE_RNI6QCS5_LC_5_5_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.WRITE_CYCLE_RNI6QCS5_LC_5_5_4 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U400_SDRAM.WRITE_CYCLE_RNI6QCS5_LC_5_5_4  (
            .in0(N__5339),
            .in1(N__3517),
            .in2(N__3506),
            .in3(N__3688),
            .lcout(\U400_SDRAM.N_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_5_5_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_5_5_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_5_5_5  (
            .in0(N__4227),
            .in1(N__4248),
            .in2(N__4166),
            .in3(N__4264),
            .lcout(\U400_SDRAM.N_44 ),
            .ltout(\U400_SDRAM.N_44_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_0_LC_5_5_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_0_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_0_LC_5_5_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_0_LC_5_5_6  (
            .in0(N__4467),
            .in1(N__4724),
            .in2(N__3794),
            .in3(N__5048),
            .lcout(\U400_SDRAM.N_108 ),
            .ltout(\U400_SDRAM.N_108_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIKV4N1_1_LC_5_5_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIKV4N1_1_LC_5_5_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIKV4N1_1_LC_5_5_7 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIKV4N1_1_LC_5_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3755),
            .in3(N__4553),
            .lcout(\U400_SDRAM.N_109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_1_0_LC_5_6_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_1_0_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_1_0_LC_5_6_1 .LUT_INIT=16'b1110111111001111;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_1_0_LC_5_6_1  (
            .in0(N__3732),
            .in1(N__4064),
            .in2(N__5335),
            .in3(N__4377),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_0_LC_5_6_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_0_LC_5_6_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_0_LC_5_6_2 .LUT_INIT=16'b0000001110101010;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_0_LC_5_6_2  (
            .in0(N__3716),
            .in1(N__3701),
            .in2(N__3692),
            .in3(N__4199),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_0C_net ),
            .ce(N__4149),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNITAGQ1_3_LC_5_6_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNITAGQ1_3_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNITAGQ1_3_LC_5_6_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNITAGQ1_3_LC_5_6_4  (
            .in0(N__4725),
            .in1(N__3856),
            .in2(N__4496),
            .in3(N__4050),
            .lcout(\U400_SDRAM.SDRAM_CMD_3_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_3_LC_5_6_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_3_LC_5_6_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_3_LC_5_6_7 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_3_LC_5_6_7  (
            .in0(N__4198),
            .in1(N__3671),
            .in2(N__4277),
            .in3(N__3644),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_0C_net ),
            .ce(N__4149),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIR5PD_3_LC_5_7_0 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIR5PD_3_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIR5PD_3_LC_5_7_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIR5PD_3_LC_5_7_0  (
            .in0(_gnd_net_),
            .in1(N__4470),
            .in2(_gnd_net_),
            .in3(N__4742),
            .lcout(\U400_SDRAM.N_46 ),
            .ltout(\U400_SDRAM.N_46_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNII7IR_0_LC_5_7_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNII7IR_0_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNII7IR_0_LC_5_7_1 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNII7IR_0_LC_5_7_1  (
            .in0(N__4599),
            .in1(_gnd_net_),
            .in2(N__3638),
            .in3(N__5053),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI189H2_0_LC_5_7_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI189H2_0_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI189H2_0_LC_5_7_2 .LUT_INIT=16'b0111001111111111;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI189H2_0_LC_5_7_2  (
            .in0(N__4915),
            .in1(N__5296),
            .in2(N__3884),
            .in3(N__3816),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIKPF05_LC_5_7_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIKPF05_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIKPF05_LC_5_7_3 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNIKPF05_LC_5_7_3  (
            .in0(N__4386),
            .in1(N__4051),
            .in2(N__3881),
            .in3(N__4988),
            .lcout(\U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIO2PD_0_LC_5_7_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIO2PD_0_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIO2PD_0_LC_5_7_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIO2PD_0_LC_5_7_5  (
            .in0(N__4743),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5054),
            .lcout(\U400_SDRAM.N_336_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_4_2_LC_5_7_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_4_2_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_4_2_LC_5_7_6 .LUT_INIT=16'b0000011100000000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_4_2_LC_5_7_6  (
            .in0(N__4969),
            .in1(N__4744),
            .in2(N__3872),
            .in3(N__4385),
            .lcout(),
            .ltout(\U400_SDRAM.N_97_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_3_2_LC_5_7_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_3_2_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_3_2_LC_5_7_7 .LUT_INIT=16'b1111000011111100;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_3_2_LC_5_7_7  (
            .in0(_gnd_net_),
            .in1(N__4812),
            .in2(N__3863),
            .in3(N__3860),
            .lcout(\U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_0_LC_5_8_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_0_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_0_LC_5_8_1 .LUT_INIT=16'b1111111110101111;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_1_0_LC_5_8_1  (
            .in0(N__4757),
            .in1(_gnd_net_),
            .in2(N__5322),
            .in3(N__4918),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_cnst_0_1_66_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_0_LC_5_8_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_0_LC_5_8_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_CMD_0_LC_5_8_2 .LUT_INIT=16'b1110111011100100;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_0_LC_5_8_2  (
            .in0(N__4016),
            .in1(N__5722),
            .in2(N__3845),
            .in3(N__4994),
            .lcout(\U400_SDRAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_CMD_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_RNO_0_5_LC_5_8_3 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_RNO_0_5_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.MA_nesr_RNO_0_5_LC_5_8_3 .LUT_INIT=16'b0011111100101110;
    LogicCell40 \U400_SDRAM.MA_nesr_RNO_0_5_LC_5_8_3  (
            .in0(N__5843),
            .in1(N__6529),
            .in2(N__3842),
            .in3(N__5713),
            .lcout(\U400_SDRAM.MA_5_iv_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_2_LC_5_8_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_2_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_2_LC_5_8_4 .LUT_INIT=16'b1111111111010000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_1_2_LC_5_8_4  (
            .in0(N__4750),
            .in1(N__3824),
            .in2(N__5084),
            .in3(N__3800),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_2_LC_5_8_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_2_LC_5_8_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_CMD_2_LC_5_8_5 .LUT_INIT=16'b1111110010101010;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_2_LC_5_8_5  (
            .in0(N__6538),
            .in1(N__3998),
            .in2(N__4019),
            .in3(N__4015),
            .lcout(\U400_SDRAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_CMD_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_2_LC_5_8_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_2_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_2_LC_5_8_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_2_2_LC_5_8_6  (
            .in0(N__4749),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5077),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_a2_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_2_LC_5_8_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_2_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_2_LC_5_8_7 .LUT_INIT=16'b0111011101110101;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_0_2_LC_5_8_7  (
            .in0(N__5292),
            .in1(N__4387),
            .in2(N__4001),
            .in3(N__4917),
            .lcout(\U400_SDRAM.SDRAM_CMD_cnst_0_143_i_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_3_LC_5_13_0 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_3_LC_5_13_0 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_3_LC_5_13_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U400_SDRAM.MA_nesr_3_LC_5_13_0  (
            .in0(N__6456),
            .in1(N__3992),
            .in2(N__6578),
            .in3(N__3983),
            .lcout(MA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_3C_net ),
            .ce(N__6418),
            .sr(N__6355));
    defparam \U400_SDRAM.MA_nesr_12_LC_5_13_6 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_12_LC_5_13_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_12_LC_5_13_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U400_SDRAM.MA_nesr_12_LC_5_13_6  (
            .in0(N__6549),
            .in1(N__5866),
            .in2(N__3953),
            .in3(N__5725),
            .lcout(MA_c_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_3C_net ),
            .ce(N__6418),
            .sr(N__6355));
    defparam \U400_SDRAM.MA_nesr_5_LC_5_13_7 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_5_LC_5_13_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_5_LC_5_13_7 .LUT_INIT=16'b1011101100110011;
    LogicCell40 \U400_SDRAM.MA_nesr_5_LC_5_13_7  (
            .in0(N__3920),
            .in1(N__3905),
            .in2(_gnd_net_),
            .in3(N__6455),
            .lcout(MA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_3C_net ),
            .ce(N__6418),
            .sr(N__6355));
    defparam \U400_SDRAM.SDRAM_CMD_RNIMFKP_0_LC_5_14_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNIMFKP_0_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNIMFKP_0_LC_5_14_1 .LUT_INIT=16'b1111011011110111;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNIMFKP_0_LC_5_14_1  (
            .in0(N__6577),
            .in1(N__5861),
            .in2(N__6371),
            .in3(N__5723),
            .lcout(\U400_SDRAM.un1_MA21_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNI06O9_0_LC_5_14_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNI06O9_0_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNI06O9_0_LC_5_14_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNI06O9_0_LC_5_14_3  (
            .in0(N__6576),
            .in1(N__5862),
            .in2(_gnd_net_),
            .in3(N__5724),
            .lcout(\U400_SDRAM.MA20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_6_LC_6_5_0 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_6_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_6_LC_6_5_0 .LUT_INIT=16'b1111111110110011;
    LogicCell40 \U400_SDRAM.TACK_RNO_6_LC_6_5_0  (
            .in0(N__4738),
            .in1(N__4400),
            .in2(N__4502),
            .in3(N__4900),
            .lcout(\U400_SDRAM.un1_SDRAM_COUNTER59_4_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI5LLK_0_LC_6_5_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI5LLK_0_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI5LLK_0_LC_6_5_1 .LUT_INIT=16'b0100010000100010;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI5LLK_0_LC_6_5_1  (
            .in0(N__4476),
            .in1(N__4643),
            .in2(_gnd_net_),
            .in3(N__5050),
            .lcout(\U400_SDRAM.N_8 ),
            .ltout(\U400_SDRAM.N_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_4_LC_6_5_2 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_4_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_4_LC_6_5_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U400_SDRAM.TACK_RNO_4_LC_6_5_2  (
            .in0(N__4249),
            .in1(N__4978),
            .in2(N__4091),
            .in3(N__4228),
            .lcout(\U400_SDRAM.N_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_RNIPSFM_0_LC_6_5_3 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_RNIPSFM_0_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_COUNTER_RNIPSFM_0_LC_6_5_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_RNIPSFM_0_LC_6_5_3  (
            .in0(_gnd_net_),
            .in1(N__5204),
            .in2(_gnd_net_),
            .in3(N__5165),
            .lcout(\U400_SDRAM.N_244_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_3_LC_6_5_4 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_3_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_3_LC_6_5_4 .LUT_INIT=16'b0111001011110000;
    LogicCell40 \U400_SDRAM.TACK_RNO_3_LC_6_5_4  (
            .in0(N__5052),
            .in1(N__4737),
            .in2(N__4817),
            .in3(N__4649),
            .lcout(),
            .ltout(\U400_SDRAM.N_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_0_LC_6_5_5 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_0_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_0_LC_6_5_5 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U400_SDRAM.TACK_RNO_0_LC_6_5_5  (
            .in0(N__4058),
            .in1(N__4088),
            .in2(N__4082),
            .in3(N__4079),
            .lcout(\U400_SDRAM.N_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_4_0_LC_6_5_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_4_0_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_4_0_LC_6_5_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_4_0_LC_6_5_6  (
            .in0(N__4739),
            .in1(N__4650),
            .in2(N__4503),
            .in3(N__4052),
            .lcout(\U400_SDRAM.N_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_5_LC_6_5_7 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_5_LC_6_5_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_5_LC_6_5_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U400_SDRAM.TACK_RNO_5_LC_6_5_7  (
            .in0(N__4477),
            .in1(N__4644),
            .in2(N__4982),
            .in3(N__5051),
            .lcout(\U400_SDRAM.N_88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNID8F21_0_LC_6_6_0 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNID8F21_0_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNID8F21_0_LC_6_6_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNID8F21_0_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(N__5047),
            .in2(_gnd_net_),
            .in3(N__4888),
            .lcout(\U400_SDRAM.N_48 ),
            .ltout(),
            .carryin(bfn_6_6_0_),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_1_1_LC_6_6_1 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_1_1_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_1_1_LC_6_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_1_1_LC_6_6_1  (
            .in0(_gnd_net_),
            .in1(N__4651),
            .in2(_gnd_net_),
            .in3(N__4283),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_s_1 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_2_LC_6_6_2 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_2_LC_6_6_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_2_LC_6_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_2_LC_6_6_2  (
            .in0(N__4200),
            .in1(N__4740),
            .in2(_gnd_net_),
            .in3(N__4280),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_2 ),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__4150),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_1_3_LC_6_6_3 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_1_3_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_1_3_LC_6_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_1_3_LC_6_6_3  (
            .in0(_gnd_net_),
            .in1(N__4501),
            .in2(_gnd_net_),
            .in3(N__4268),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_s_3 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_4_LC_6_6_4 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_4_LC_6_6_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_4_LC_6_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_4_LC_6_6_4  (
            .in0(N__4201),
            .in1(N__4265),
            .in2(_gnd_net_),
            .in3(N__4253),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_4 ),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__4150),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_5_LC_6_6_5 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_5_LC_6_6_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_5_LC_6_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_5_LC_6_6_5  (
            .in0(N__4208),
            .in1(N__4250),
            .in2(_gnd_net_),
            .in3(N__4232),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_5 ),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__4150),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_6_LC_6_6_6 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_6_LC_6_6_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_6_LC_6_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_6_LC_6_6_6  (
            .in0(N__4202),
            .in1(N__4229),
            .in2(_gnd_net_),
            .in3(N__4211),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_6 ),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__4150),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_7_LC_6_6_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_7_LC_6_6_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_7_LC_6_6_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_7_LC_6_6_7  (
            .in0(N__4165),
            .in1(N__4203),
            .in2(_gnd_net_),
            .in3(N__4169),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__4150),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_7_LC_6_7_0 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_7_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_7_LC_6_7_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U400_SDRAM.TACK_RNO_7_LC_6_7_0  (
            .in0(N__4971),
            .in1(N__4728),
            .in2(N__4856),
            .in3(N__4913),
            .lcout(),
            .ltout(\U400_SDRAM.N_56_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_2_LC_6_7_1 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_2_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_2_LC_6_7_1 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \U400_SDRAM.TACK_RNO_2_LC_6_7_1  (
            .in0(N__4121),
            .in1(N__4972),
            .in2(N__4109),
            .in3(N__4653),
            .lcout(\U400_SDRAM.TACK_7_iv_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_0_LC_6_7_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_0_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_0_LC_6_7_3 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_0_0_LC_6_7_3  (
            .in0(N__4925),
            .in1(N__4652),
            .in2(_gnd_net_),
            .in3(N__5068),
            .lcout(\U400_SDRAM.N_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNITTB91_3_LC_6_7_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNITTB91_3_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNITTB91_3_LC_6_7_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNITTB91_3_LC_6_7_4  (
            .in0(N__4478),
            .in1(N__4726),
            .in2(_gnd_net_),
            .in3(N__4912),
            .lcout(\U400_SDRAM.N_110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.WRITE_CYCLE_RNIT04E_LC_6_7_6 .C_ON=1'b0;
    defparam \U400_SDRAM.WRITE_CYCLE_RNIT04E_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.WRITE_CYCLE_RNIT04E_LC_6_7_6 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \U400_SDRAM.WRITE_CYCLE_RNIT04E_LC_6_7_6  (
            .in0(N__4970),
            .in1(N__4727),
            .in2(_gnd_net_),
            .in3(N__4403),
            .lcout(\U400_SDRAM.N_13 ),
            .ltout(\U400_SDRAM.N_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_RNO_1_LC_6_7_7 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_1_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_1_LC_6_7_7 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_RNO_1_LC_6_7_7  (
            .in0(N__4914),
            .in1(N__4855),
            .in2(N__4841),
            .in3(N__4838),
            .lcout(\U400_SDRAM.un1_SDRAM_COUNTER59_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_4_0_LC_6_8_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_4_0_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_4_0_LC_6_8_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_4_0_LC_6_8_3  (
            .in0(N__4402),
            .in1(N__4805),
            .in2(_gnd_net_),
            .in3(N__4648),
            .lcout(),
            .ltout(\U400_SDRAM.N_33_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_0_LC_6_8_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_0_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_0_LC_6_8_4 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_2_0_LC_6_8_4  (
            .in0(N__4500),
            .in1(N__4289),
            .in2(N__4784),
            .in3(N__4781),
            .lcout(\U400_SDRAM.SDRAM_CMD_cnst_0_1_66_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_3_0_LC_6_8_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_3_0_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_3_0_LC_6_8_6 .LUT_INIT=16'b0000000011011010;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_3_0_LC_6_8_6  (
            .in0(N__4748),
            .in1(N__4647),
            .in2(N__4507),
            .in3(N__4401),
            .lcout(\U400_SDRAM.N_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_0_LC_7_4_0 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_0_LC_7_4_0 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.TA_COUNTER_0_LC_7_4_0 .LUT_INIT=16'b0010000011111111;
    LogicCell40 \U400_SDRAM.TA_COUNTER_0_LC_7_4_0  (
            .in0(N__5360),
            .in1(N__5179),
            .in2(N__5138),
            .in3(N__5354),
            .lcout(\U400_SDRAM.TA_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5494),
            .ce(),
            .sr(N__6357));
    defparam \U400_SDRAM.TA_EN_i_LC_7_4_2 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_EN_i_LC_7_4_2 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.TA_EN_i_LC_7_4_2 .LUT_INIT=16'b0011111110101010;
    LogicCell40 \U400_SDRAM.TA_EN_i_LC_7_4_2  (
            .in0(N__6223),
            .in1(N__5122),
            .in2(N__5338),
            .in3(N__5144),
            .lcout(TA_EN_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5494),
            .ce(),
            .sr(N__6357));
    defparam \U400_SDRAM.TA_COUNTER_2_LC_7_4_3 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_2_LC_7_4_3 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_2_LC_7_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_2_LC_7_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5668),
            .lcout(\U400_SDRAM.TA_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5494),
            .ce(),
            .sr(N__6357));
    defparam \U400_SDRAM.TA_COUNTER_1_LC_7_4_4 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_1_LC_7_4_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_1_LC_7_4_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_1_LC_7_4_4  (
            .in0(_gnd_net_),
            .in1(N__5203),
            .in2(_gnd_net_),
            .in3(N__5178),
            .lcout(\U400_SDRAM.TA_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5494),
            .ce(),
            .sr(N__6357));
    defparam \U400_SDRAM.TA_COUNTER_RNO_0_0_LC_7_5_0 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_RNO_0_0_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_COUNTER_RNO_0_0_LC_7_5_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U400_SDRAM.TA_COUNTER_RNO_0_0_LC_7_5_0  (
            .in0(N__5524),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5509),
            .lcout(\U400_SDRAM.TA_COUNTER_srsts_0_a4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_RNINB8O_1_LC_7_5_2 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_RNINB8O_1_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_COUNTER_RNINB8O_1_LC_7_5_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U400_SDRAM.TA_COUNTER_RNINB8O_1_LC_7_5_2  (
            .in0(N__5550),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5667),
            .lcout(\U400_SDRAM.un1_TA_COUNTER_6_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_RNIMKDP_5_LC_7_5_3 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_RNIMKDP_5_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_COUNTER_RNIMKDP_5_LC_7_5_3 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \U400_SDRAM.TA_COUNTER_RNIMKDP_5_LC_7_5_3  (
            .in0(N__5531),
            .in1(N__5523),
            .in2(_gnd_net_),
            .in3(N__5381),
            .lcout(\U400_SDRAM.N_243_0 ),
            .ltout(\U400_SDRAM.N_243_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_EN_i_RNO_0_LC_7_5_4 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_EN_i_RNO_0_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_EN_i_RNO_0_LC_7_5_4 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \U400_SDRAM.TA_EN_i_RNO_0_LC_7_5_4  (
            .in0(N__5323),
            .in1(N__5202),
            .in2(N__5183),
            .in3(N__5180),
            .lcout(\U400_SDRAM.N_241_0_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_OUT_LC_7_6_7 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_OUT_LC_7_6_7 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.TA_OUT_LC_7_6_7 .LUT_INIT=16'b0011001110110001;
    LogicCell40 \U400_SDRAM.TA_OUT_LC_7_6_7  (
            .in0(N__5137),
            .in1(N__5648),
            .in2(N__5110),
            .in3(N__5123),
            .lcout(TA_OUT),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5492),
            .ce(),
            .sr(N__6354));
    defparam \U400_BYTE_ENABLE.un1_UUBEn_i_0_LC_7_7_2 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un1_UUBEn_i_0_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un1_UUBEn_i_0_LC_7_7_2 .LUT_INIT=16'b1111101011101010;
    LogicCell40 \U400_BYTE_ENABLE.un1_UUBEn_i_0_LC_7_7_2  (
            .in0(N__5979),
            .in1(N__5919),
            .in2(N__6041),
            .in3(N__6025),
            .lcout(N_53),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_OUT_RNO_0_LC_7_7_6 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_OUT_RNO_0_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_OUT_RNO_0_LC_7_7_6 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \U400_SDRAM.TA_OUT_RNO_0_LC_7_7_6  (
            .in0(N__5552),
            .in1(N__5669),
            .in2(_gnd_net_),
            .in3(N__5382),
            .lcout(\U400_SDRAM.TA_OUT_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_11_LC_7_15_2 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_11_LC_7_15_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_11_LC_7_15_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U400_SDRAM.MA_nesr_11_LC_7_15_2  (
            .in0(N__6612),
            .in1(N__5868),
            .in2(N__5642),
            .in3(N__5763),
            .lcout(MA_c_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_11C_net ),
            .ce(N__6422),
            .sr(N__6362));
    defparam \U400_SDRAM.MA_nesr_9_LC_7_15_6 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_9_LC_7_15_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_9_LC_7_15_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U400_SDRAM.MA_nesr_9_LC_7_15_6  (
            .in0(N__6613),
            .in1(N__5764),
            .in2(N__5878),
            .in3(N__5609),
            .lcout(MA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_11C_net ),
            .ce(N__6422),
            .sr(N__6362));
    defparam \U400_SDRAM.MA_nesr_8_LC_7_15_7 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_8_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_8_LC_7_15_7 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U400_SDRAM.MA_nesr_8_LC_7_15_7  (
            .in0(N__5588),
            .in1(N__6614),
            .in2(N__5576),
            .in3(N__6481),
            .lcout(MA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_11C_net ),
            .ce(N__6422),
            .sr(N__6362));
    defparam \U400_SDRAM.TA_COUNTER_4_LC_8_5_0 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_4_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_4_LC_8_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_4_LC_8_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5510),
            .lcout(\U400_SDRAM.TA_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5495),
            .ce(),
            .sr(N__6358));
    defparam \U400_SDRAM.TA_COUNTER_5_LC_8_5_2 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_5_LC_8_5_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_5_LC_8_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_5_LC_8_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5551),
            .lcout(\U400_SDRAM.TA_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5495),
            .ce(),
            .sr(N__6358));
    defparam \U400_SDRAM.TA_COUNTER_3_LC_8_5_6 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_3_LC_8_5_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_3_LC_8_5_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_3_LC_8_5_6  (
            .in0(_gnd_net_),
            .in1(N__5525),
            .in2(_gnd_net_),
            .in3(N__5383),
            .lcout(\U400_SDRAM.TA_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5495),
            .ce(),
            .sr(N__6358));
    defparam \U400_SDRAM.BURST_LC_8_6_7 .C_ON=1'b0;
    defparam \U400_SDRAM.BURST_LC_8_6_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.BURST_LC_8_6_7 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U400_SDRAM.BURST_LC_8_6_7  (
            .in0(N__6172),
            .in1(N__5384),
            .in2(N__6082),
            .in3(N__5416),
            .lcout(\U400_SDRAM.BURSTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.BURSTC_net ),
            .ce(),
            .sr(N__6356));
    defparam \U400_SDRAM.MA_nesr_10_LC_8_16_2 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_10_LC_8_16_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_10_LC_8_16_2 .LUT_INIT=16'b0100000001000100;
    LogicCell40 \U400_SDRAM.MA_nesr_10_LC_8_16_2  (
            .in0(N__6616),
            .in1(N__5879),
            .in2(N__6299),
            .in3(N__5765),
            .lcout(MA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_10C_net ),
            .ce(N__6419),
            .sr(N__6363));
    defparam \U400_SDRAM.MA_nesr_0_LC_8_16_5 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_0_LC_8_16_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_0_LC_8_16_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \U400_SDRAM.MA_nesr_0_LC_8_16_5  (
            .in0(N__6278),
            .in1(N__6615),
            .in2(N__6266),
            .in3(N__6482),
            .lcout(MA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_10C_net ),
            .ce(N__6419),
            .sr(N__6363));
    defparam \U400_BYTE_ENABLE.un1_UMBEn_i_0_LC_9_3_1 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un1_UMBEn_i_0_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un1_UMBEn_i_0_LC_9_3_1 .LUT_INIT=16'b1111111100101000;
    LogicCell40 \U400_BYTE_ENABLE.un1_UMBEn_i_0_LC_9_3_1  (
            .in0(N__5933),
            .in1(N__6186),
            .in2(N__6113),
            .in3(N__6200),
            .lcout(N_51),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_BYTE_ENABLE.un1_LLBEn_i_0_LC_9_3_3 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un1_LLBEn_i_0_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un1_LLBEn_i_0_LC_9_3_3 .LUT_INIT=16'b1111111100010100;
    LogicCell40 \U400_BYTE_ENABLE.un1_LLBEn_i_0_LC_9_3_3  (
            .in0(N__5932),
            .in1(N__6185),
            .in2(N__6112),
            .in3(N__6199),
            .lcout(N_47),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TAn_obuft_RNO_LC_9_4_3.C_ON=1'b0;
    defparam TAn_obuft_RNO_LC_9_4_3.SEQ_MODE=4'b0000;
    defparam TAn_obuft_RNO_LC_9_4_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 TAn_obuft_RNO_LC_9_4_3 (
            .in0(N__6227),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_542_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_BYTE_ENABLE.un1_LLBEn_i_o3_LC_9_4_5 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un1_LLBEn_i_o3_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un1_LLBEn_i_o3_LC_9_4_5 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \U400_BYTE_ENABLE.un1_LLBEn_i_o3_LC_9_4_5  (
            .in0(N__6173),
            .in1(N__6083),
            .in2(N__5978),
            .in3(N__6026),
            .lcout(\U400_BYTE_ENABLE.N_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_BYTE_ENABLE.un1_LLBEn_i_x2_LC_9_8_6 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un1_LLBEn_i_x2_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un1_LLBEn_i_x2_LC_9_8_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \U400_BYTE_ENABLE.un1_LLBEn_i_x2_LC_9_8_6  (
            .in0(N__6171),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6057),
            .lcout(\U400_BYTE_ENABLE.N_54_i ),
            .ltout(\U400_BYTE_ENABLE.N_54_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_BYTE_ENABLE.un1_LMBEn_i_0_LC_9_8_7 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un1_LMBEn_i_0_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un1_LMBEn_i_0_LC_9_8_7 .LUT_INIT=16'b1110110011111100;
    LogicCell40 \U400_BYTE_ENABLE.un1_LMBEn_i_0_LC_9_8_7  (
            .in0(N__6021),
            .in1(N__5980),
            .in2(N__5936),
            .in3(N__5926),
            .lcout(N_49),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_RNO_0_1_LC_9_15_5 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_RNO_0_1_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.MA_nesr_RNO_0_1_LC_9_15_5 .LUT_INIT=16'b0101111101001110;
    LogicCell40 \U400_SDRAM.MA_nesr_RNO_0_1_LC_9_15_5  (
            .in0(N__6596),
            .in1(N__5867),
            .in2(N__5780),
            .in3(N__5754),
            .lcout(\U400_SDRAM.MA_5_iv_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_1_LC_9_16_4 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_1_LC_9_16_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_1_LC_9_16_4 .LUT_INIT=16'b1011101100110011;
    LogicCell40 \U400_SDRAM.MA_nesr_1_LC_9_16_4  (
            .in0(N__6656),
            .in1(N__6644),
            .in2(_gnd_net_),
            .in3(N__6479),
            .lcout(MA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_1C_net ),
            .ce(N__6420),
            .sr(N__6364));
    defparam \U400_SDRAM.MA_nesr_2_LC_9_16_6 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_2_LC_9_16_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_2_LC_9_16_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \U400_SDRAM.MA_nesr_2_LC_9_16_6  (
            .in0(N__6632),
            .in1(N__6617),
            .in2(N__6491),
            .in3(N__6480),
            .lcout(MA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_1C_net ),
            .ce(N__6420),
            .sr(N__6364));
endmodule // U400_TOP

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 16 2024 18:13:15

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    A : in std_logic_vector(20 downto 0);
    TSn : in std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    LDSn : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    DBRn : in std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RAMENn : out std_logic;
    RASn : out std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__9911\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7827\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7257\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3928\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3873\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3715\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3693\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3669\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3654\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3622\ : std_logic;
signal \N__3619\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3547\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK80_OUT_i_i\ : std_logic;
signal \CLK40_OUT_i_i\ : std_logic;
signal \U712_REG_SM.LDS_OUT_2_0_a2Z0Z_0\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_387_cascade_\ : std_logic;
signal \N_73_i\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_REG_SM.N_301\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \U712_REG_SM.N_281_cascade_\ : std_logic;
signal \U712_REG_SM.N_280_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_308\ : std_logic;
signal \U712_REG_SM.N_288_cascade_\ : std_logic;
signal \U712_REG_SM.N_307\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_2\ : std_logic;
signal \C3_c\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2Z0Z_0\ : std_logic;
signal \N_75_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_395\ : std_logic;
signal \N_74_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_387\ : std_logic;
signal \A_c_1\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_0_0\ : std_logic;
signal \N_76_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_391\ : std_logic;
signal \U712_REG_SM.N_304\ : std_logic;
signal \U712_REG_SM.N_299\ : std_logic;
signal \U712_REG_SM.N_281\ : std_logic;
signal \U712_REG_SM.N_280\ : std_logic;
signal \U712_REG_SM.N_373_cascade_\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_2\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_289\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_6\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_289_cascade_\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_494\ : std_logic;
signal \U712_REG_SM.N_288\ : std_logic;
signal \U712_REG_SM.N_494_cascade_\ : std_logic;
signal \U712_REG_SM.N_424\ : std_logic;
signal \U712_REG_SM.N_369\ : std_logic;
signal \U712_REG_SM.DS_EN_RNOZ0Z_2_cascade_\ : std_logic;
signal \U712_REG_SM.N_123\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \CLK40_OUT_i\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\ : std_logic;
signal \N_886_i\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_2_cascade_\ : std_logic;
signal \A_c_11\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_REG_SM.N_306\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_5\ : std_logic;
signal \U712_REG_SM.N_298\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.UDS_OUTZ0\ : std_logic;
signal \U712_REG_SM_un1_UDSn_i\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.N_305_i_0_en_cascade_\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.N_341_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_1_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\ : std_logic;
signal \U712_BYTE_ENABLE.N_392\ : std_logic;
signal \U712_BYTE_ENABLE.N_388\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \TSn_c\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \U712_CYCLE_TERM.N_305_i_0_en_0\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \A_c_7\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \A_c_9\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \A_c_10\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_1_cascade_\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \U712_CHIP_RAM.N_313\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_3_cascade_\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U712_CHIP_RAM.N_314_cascade_\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_5\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_6_cascade_\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_0\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_3_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_2_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_421_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_293_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_309_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0_a2_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_REG_SM.DS_ENZ0\ : std_logic;
signal \U712_REG_SM.LDS_OUTZ0\ : std_logic;
signal \U712_REG_SM_un1_LDSn_i\ : std_logic;
signal \U712_CHIP_RAM.N_311\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.N_312\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.N_316\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA31_0_i_cascade_\ : std_logic;
signal \A_c_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_4\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U712_CHIP_RAM.N_493_cascade_\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_317\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \A_c_19\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_i_0_8_cascade_\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_285\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_7_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_0_a2_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_427\ : std_logic;
signal \U712_CHIP_RAM.N_421\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_296\ : std_logic;
signal \U712_CHIP_RAM.N_296_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_i_0_a2_0_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_403\ : std_logic;
signal \U712_CHIP_RAM.N_309\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER46_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_420\ : std_logic;
signal \U712_CHIP_RAM.N_282\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_a5_i_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_49\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \N_218\ : std_logic;
signal \RASn_c\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_7_cascade_\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_i_0_8\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.N_318\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_315\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA31_0_i_0\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \RnW_c\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_i_a2_1_0_a2_1_0\ : std_logic;
signal \U712_CHIP_RAM.N_284\ : std_logic;
signal \U712_CHIP_RAM.N_284_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_1_2\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_1_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c6_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_0_3\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.N_274\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U712_CHIP_RAM.N_274_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_337\ : std_logic;
signal \U712_CHIP_RAM.N_337_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_2_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_271\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_5_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER46\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_303\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \WEn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_1\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    CLK_EN <= \CLK_EN_wire\;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    LDSn <= \LDSn_wire\;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_OUT_i\,
            REFERENCECLK => \N__3553\,
            RESETB => \N__8836\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_OUT\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9911\,
            DIN => \N__9910\,
            DOUT => \N__9909\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9911\,
            PADOUT => \N__9910\,
            PADIN => \N__9909\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6190\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9902\,
            DIN => \N__9901\,
            DOUT => \N__9900\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9902\,
            PADOUT => \N__9901\,
            PADIN => \N__9900\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9893\,
            DIN => \N__9892\,
            DOUT => \N__9891\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9893\,
            PADOUT => \N__9892\,
            PADIN => \N__9891\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8461\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9884\,
            DIN => \N__9883\,
            DOUT => \N__9882\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9884\,
            PADOUT => \N__9883\,
            PADIN => \N__9882\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6397\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9875\,
            DIN => \N__9874\,
            DOUT => \N__9873\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9875\,
            PADOUT => \N__9874\,
            PADIN => \N__9873\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9866\,
            DIN => \N__9865\,
            DOUT => \N__9864\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9866\,
            PADOUT => \N__9865\,
            PADIN => \N__9864\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9857\,
            DIN => \N__9856\,
            DOUT => \N__9855\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9857\,
            PADOUT => \N__9856\,
            PADIN => \N__9855\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9848\,
            DIN => \N__9847\,
            DOUT => \N__9846\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9848\,
            PADOUT => \N__9847\,
            PADIN => \N__9846\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9839\,
            DIN => \N__9838\,
            DOUT => \N__9837\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9839\,
            PADOUT => \N__9838\,
            PADIN => \N__9837\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9830\,
            DIN => \N__9829\,
            DOUT => \N__9828\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9830\,
            PADOUT => \N__9829\,
            PADIN => \N__9828\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9821\,
            DIN => \N__9820\,
            DOUT => \N__9819\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9821\,
            PADOUT => \N__9820\,
            PADIN => \N__9819\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7129\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9812\,
            DIN => \N__9811\,
            DOUT => \N__9810\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9812\,
            PADOUT => \N__9811\,
            PADIN => \N__9810\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5166\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9803\,
            DIN => \N__9802\,
            DOUT => \N__9801\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9803\,
            PADOUT => \N__9802\,
            PADIN => \N__9801\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9794\,
            DIN => \N__9793\,
            DOUT => \N__9792\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9794\,
            PADOUT => \N__9793\,
            PADIN => \N__9792\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9785\,
            DIN => \N__9784\,
            DOUT => \N__9783\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9785\,
            PADOUT => \N__9784\,
            PADIN => \N__9783\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3571\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9776\,
            DIN => \N__9775\,
            DOUT => \N__9774\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9776\,
            PADOUT => \N__9775\,
            PADIN => \N__9774\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9767\,
            DIN => \N__9766\,
            DOUT => \N__9765\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9767\,
            PADOUT => \N__9766\,
            PADIN => \N__9765\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9758\,
            DIN => \N__9757\,
            DOUT => \N__9756\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9758\,
            PADOUT => \N__9757\,
            PADIN => \N__9756\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5881\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9749\,
            DIN => \N__9748\,
            DOUT => \N__9747\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9749\,
            PADOUT => \N__9748\,
            PADIN => \N__9747\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9740\,
            DIN => \N__9739\,
            DOUT => \N__9738\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9740\,
            PADOUT => \N__9739\,
            PADIN => \N__9738\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8296\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9731\,
            DIN => \N__9730\,
            DOUT => \N__9729\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9731\,
            PADOUT => \N__9730\,
            PADIN => \N__9729\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9722\,
            DIN => \N__9721\,
            DOUT => \N__9720\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9722\,
            PADOUT => \N__9721\,
            PADIN => \N__9720\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9713\,
            DIN => \N__9712\,
            DOUT => \N__9711\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9713\,
            PADOUT => \N__9712\,
            PADIN => \N__9711\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9704\,
            DIN => \N__9703\,
            DOUT => \N__9702\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9704\,
            PADOUT => \N__9703\,
            PADIN => \N__9702\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9695\,
            DIN => \N__9694\,
            DOUT => \N__9693\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9695\,
            PADOUT => \N__9694\,
            PADIN => \N__9693\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9686\,
            DIN => \N__9685\,
            DOUT => \N__9684\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9686\,
            PADOUT => \N__9685\,
            PADIN => \N__9684\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8829\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9677\,
            DIN => \N__9676\,
            DOUT => \N__9675\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9677\,
            PADOUT => \N__9676\,
            PADIN => \N__9675\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9668\,
            DIN => \N__9667\,
            DOUT => \N__9666\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9668\,
            PADOUT => \N__9667\,
            PADIN => \N__9666\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9659\,
            DIN => \N__9658\,
            DOUT => \N__9657\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9659\,
            PADOUT => \N__9658\,
            PADIN => \N__9657\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9650\,
            DIN => \N__9649\,
            DOUT => \N__9648\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9650\,
            PADOUT => \N__9649\,
            PADIN => \N__9648\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9641\,
            DIN => \N__9640\,
            DOUT => \N__9639\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9641\,
            PADOUT => \N__9640\,
            PADIN => \N__9639\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9632\,
            DIN => \N__9631\,
            DOUT => \N__9630\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9632\,
            PADOUT => \N__9631\,
            PADIN => \N__9630\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6043\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9623\,
            DIN => \N__9622\,
            DOUT => \N__9621\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9623\,
            PADOUT => \N__9622\,
            PADIN => \N__9621\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9614\,
            DIN => \N__9613\,
            DOUT => \N__9612\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9614\,
            PADOUT => \N__9613\,
            PADIN => \N__9612\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9605\,
            DIN => \N__9604\,
            DOUT => \N__9603\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9605\,
            PADOUT => \N__9604\,
            PADIN => \N__9603\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9596\,
            DIN => \N__9595\,
            DOUT => \N__9594\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9596\,
            PADOUT => \N__9595\,
            PADIN => \N__9594\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9587\,
            DIN => \N__9586\,
            DOUT => \N__9585\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9587\,
            PADOUT => \N__9586\,
            PADIN => \N__9585\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3595\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9578\,
            DIN => \N__9577\,
            DOUT => \N__9576\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9578\,
            PADOUT => \N__9577\,
            PADIN => \N__9576\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5908\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9569\,
            DIN => \N__9568\,
            DOUT => \N__9567\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9569\,
            PADOUT => \N__9568\,
            PADIN => \N__9567\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9560\,
            DIN => \N__9559\,
            DOUT => \N__9558\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9560\,
            PADOUT => \N__9559\,
            PADIN => \N__9558\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6382\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9551\,
            DIN => \N__9550\,
            DOUT => \N__9549\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9551\,
            PADOUT => \N__9550\,
            PADIN => \N__9549\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9542\,
            DIN => \N__9541\,
            DOUT => \N__9540\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9542\,
            PADOUT => \N__9541\,
            PADIN => \N__9540\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9533\,
            DIN => \N__9532\,
            DOUT => \N__9531\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9533\,
            PADOUT => \N__9532\,
            PADIN => \N__9531\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3610\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9524\,
            DIN => \N__9523\,
            DOUT => \N__9522\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9524\,
            PADOUT => \N__9523\,
            PADIN => \N__9522\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9515\,
            DIN => \N__9514\,
            DOUT => \N__9513\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9515\,
            PADOUT => \N__9514\,
            PADIN => \N__9513\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3874\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9506\,
            DIN => \N__9505\,
            DOUT => \N__9504\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9506\,
            PADOUT => \N__9505\,
            PADIN => \N__9504\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5659\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9497\,
            DIN => \N__9496\,
            DOUT => \N__9495\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9497\,
            PADOUT => \N__9496\,
            PADIN => \N__9495\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9488\,
            DIN => \N__9487\,
            DOUT => \N__9486\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9488\,
            PADOUT => \N__9487\,
            PADIN => \N__9486\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9479\,
            DIN => \N__9478\,
            DOUT => \N__9477\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9479\,
            PADOUT => \N__9478\,
            PADIN => \N__9477\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9470\,
            DIN => \N__9469\,
            DOUT => \N__9468\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9470\,
            PADOUT => \N__9469\,
            PADIN => \N__9468\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5371\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9461\,
            DIN => \N__9460\,
            DOUT => \N__9459\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9461\,
            PADOUT => \N__9460\,
            PADIN => \N__9459\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9452\,
            DIN => \N__9451\,
            DOUT => \N__9450\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9452\,
            PADOUT => \N__9451\,
            PADIN => \N__9450\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7012\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9443\,
            DIN => \N__9442\,
            DOUT => \N__9441\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9443\,
            PADOUT => \N__9442\,
            PADIN => \N__9441\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7468\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9434\,
            DIN => \N__9433\,
            DOUT => \N__9432\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9434\,
            PADOUT => \N__9433\,
            PADIN => \N__9432\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3715\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9425\,
            DIN => \N__9424\,
            DOUT => \N__9423\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9425\,
            PADOUT => \N__9424\,
            PADIN => \N__9423\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6004\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9416\,
            DIN => \N__9415\,
            DOUT => \N__9414\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9416\,
            PADOUT => \N__9415\,
            PADIN => \N__9414\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3873\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9407\,
            DIN => \N__9406\,
            DOUT => \N__9405\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9407\,
            PADOUT => \N__9406\,
            PADIN => \N__9405\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9398\,
            DIN => \N__9397\,
            DOUT => \N__9396\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9398\,
            PADOUT => \N__9397\,
            PADIN => \N__9396\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9389\,
            DIN => \N__9388\,
            DOUT => \N__9387\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9389\,
            PADOUT => \N__9388\,
            PADIN => \N__9387\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4186\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9380\,
            DIN => \N__9379\,
            DOUT => \N__9378\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9380\,
            PADOUT => \N__9379\,
            PADIN => \N__9378\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8350\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9371\,
            DIN => \N__9370\,
            DOUT => \N__9369\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9371\,
            PADOUT => \N__9370\,
            PADIN => \N__9369\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6436\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9362\,
            DIN => \N__9361\,
            DOUT => \N__9360\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9362\,
            PADOUT => \N__9361\,
            PADIN => \N__9360\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3916\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9353\,
            DIN => \N__9352\,
            DOUT => \N__9351\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9353\,
            PADOUT => \N__9352\,
            PADIN => \N__9351\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9344\,
            DIN => \N__9343\,
            DOUT => \N__9342\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9344\,
            PADOUT => \N__9343\,
            PADIN => \N__9342\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9335\,
            DIN => \N__9334\,
            DOUT => \N__9333\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9335\,
            PADOUT => \N__9334\,
            PADIN => \N__9333\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9326\,
            DIN => \N__9325\,
            DOUT => \N__9324\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9326\,
            PADOUT => \N__9325\,
            PADIN => \N__9324\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9317\,
            DIN => \N__9316\,
            DOUT => \N__9315\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9317\,
            PADOUT => \N__9316\,
            PADIN => \N__9315\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5857\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9308\,
            DIN => \N__9307\,
            DOUT => \N__9306\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9308\,
            PADOUT => \N__9307\,
            PADIN => \N__9306\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9299\,
            DIN => \N__9298\,
            DOUT => \N__9297\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9299\,
            PADOUT => \N__9298\,
            PADIN => \N__9297\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4108\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9290\,
            DIN => \N__9289\,
            DOUT => \N__9288\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9290\,
            PADOUT => \N__9289\,
            PADIN => \N__9288\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4528\,
            DIN0 => OPEN,
            DOUT0 => \N__4246\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9281\,
            DIN => \N__9280\,
            DOUT => \N__9279\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9281\,
            PADOUT => \N__9280\,
            PADIN => \N__9279\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5341\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9272\,
            DIN => \N__9271\,
            DOUT => \N__9270\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9272\,
            PADOUT => \N__9271\,
            PADIN => \N__9270\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9263\,
            DIN => \N__9262\,
            DOUT => \N__9261\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9263\,
            PADOUT => \N__9262\,
            PADIN => \N__9261\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9254\,
            DIN => \N__9253\,
            DOUT => \N__9252\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9254\,
            PADOUT => \N__9253\,
            PADIN => \N__9252\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7156\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9245\,
            DIN => \N__9244\,
            DOUT => \N__9243\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9245\,
            PADOUT => \N__9244\,
            PADIN => \N__9243\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9236\,
            DIN => \N__9235\,
            DOUT => \N__9234\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9236\,
            PADOUT => \N__9235\,
            PADIN => \N__9234\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9227\,
            DIN => \N__9226\,
            DOUT => \N__9225\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9227\,
            PADOUT => \N__9226\,
            PADIN => \N__9225\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9218\,
            DIN => \N__9217\,
            DOUT => \N__9216\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9218\,
            PADOUT => \N__9217\,
            PADIN => \N__9216\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9209\,
            DIN => \N__9208\,
            DOUT => \N__9207\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9209\,
            PADOUT => \N__9208\,
            PADIN => \N__9207\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5833\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9200\,
            DIN => \N__9199\,
            DOUT => \N__9198\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9200\,
            PADOUT => \N__9199\,
            PADIN => \N__9198\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4594\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2181\ : InMux
    port map (
            O => \N__9181\,
            I => \N__9177\
        );

    \I__2180\ : InMux
    port map (
            O => \N__9180\,
            I => \N__9174\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__9177\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__9174\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2177\ : InMux
    port map (
            O => \N__9169\,
            I => \N__9166\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__9166\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\
        );

    \I__2175\ : InMux
    port map (
            O => \N__9163\,
            I => \N__9160\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__9160\,
            I => \N__9136\
        );

    \I__2173\ : ClkMux
    port map (
            O => \N__9159\,
            I => \N__9034\
        );

    \I__2172\ : ClkMux
    port map (
            O => \N__9158\,
            I => \N__9034\
        );

    \I__2171\ : ClkMux
    port map (
            O => \N__9157\,
            I => \N__9034\
        );

    \I__2170\ : ClkMux
    port map (
            O => \N__9156\,
            I => \N__9034\
        );

    \I__2169\ : ClkMux
    port map (
            O => \N__9155\,
            I => \N__9034\
        );

    \I__2168\ : ClkMux
    port map (
            O => \N__9154\,
            I => \N__9034\
        );

    \I__2167\ : ClkMux
    port map (
            O => \N__9153\,
            I => \N__9034\
        );

    \I__2166\ : ClkMux
    port map (
            O => \N__9152\,
            I => \N__9034\
        );

    \I__2165\ : ClkMux
    port map (
            O => \N__9151\,
            I => \N__9034\
        );

    \I__2164\ : ClkMux
    port map (
            O => \N__9150\,
            I => \N__9034\
        );

    \I__2163\ : ClkMux
    port map (
            O => \N__9149\,
            I => \N__9034\
        );

    \I__2162\ : ClkMux
    port map (
            O => \N__9148\,
            I => \N__9034\
        );

    \I__2161\ : ClkMux
    port map (
            O => \N__9147\,
            I => \N__9034\
        );

    \I__2160\ : ClkMux
    port map (
            O => \N__9146\,
            I => \N__9034\
        );

    \I__2159\ : ClkMux
    port map (
            O => \N__9145\,
            I => \N__9034\
        );

    \I__2158\ : ClkMux
    port map (
            O => \N__9144\,
            I => \N__9034\
        );

    \I__2157\ : ClkMux
    port map (
            O => \N__9143\,
            I => \N__9034\
        );

    \I__2156\ : ClkMux
    port map (
            O => \N__9142\,
            I => \N__9034\
        );

    \I__2155\ : ClkMux
    port map (
            O => \N__9141\,
            I => \N__9034\
        );

    \I__2154\ : ClkMux
    port map (
            O => \N__9140\,
            I => \N__9034\
        );

    \I__2153\ : ClkMux
    port map (
            O => \N__9139\,
            I => \N__9034\
        );

    \I__2152\ : Glb2LocalMux
    port map (
            O => \N__9136\,
            I => \N__9034\
        );

    \I__2151\ : ClkMux
    port map (
            O => \N__9135\,
            I => \N__9034\
        );

    \I__2150\ : ClkMux
    port map (
            O => \N__9134\,
            I => \N__9034\
        );

    \I__2149\ : ClkMux
    port map (
            O => \N__9133\,
            I => \N__9034\
        );

    \I__2148\ : ClkMux
    port map (
            O => \N__9132\,
            I => \N__9034\
        );

    \I__2147\ : ClkMux
    port map (
            O => \N__9131\,
            I => \N__9034\
        );

    \I__2146\ : ClkMux
    port map (
            O => \N__9130\,
            I => \N__9034\
        );

    \I__2145\ : ClkMux
    port map (
            O => \N__9129\,
            I => \N__9034\
        );

    \I__2144\ : ClkMux
    port map (
            O => \N__9128\,
            I => \N__9034\
        );

    \I__2143\ : ClkMux
    port map (
            O => \N__9127\,
            I => \N__9034\
        );

    \I__2142\ : ClkMux
    port map (
            O => \N__9126\,
            I => \N__9034\
        );

    \I__2141\ : ClkMux
    port map (
            O => \N__9125\,
            I => \N__9034\
        );

    \I__2140\ : ClkMux
    port map (
            O => \N__9124\,
            I => \N__9034\
        );

    \I__2139\ : ClkMux
    port map (
            O => \N__9123\,
            I => \N__9034\
        );

    \I__2138\ : ClkMux
    port map (
            O => \N__9122\,
            I => \N__9034\
        );

    \I__2137\ : ClkMux
    port map (
            O => \N__9121\,
            I => \N__9034\
        );

    \I__2136\ : ClkMux
    port map (
            O => \N__9120\,
            I => \N__9034\
        );

    \I__2135\ : ClkMux
    port map (
            O => \N__9119\,
            I => \N__9034\
        );

    \I__2134\ : ClkMux
    port map (
            O => \N__9118\,
            I => \N__9034\
        );

    \I__2133\ : ClkMux
    port map (
            O => \N__9117\,
            I => \N__9034\
        );

    \I__2132\ : GlobalMux
    port map (
            O => \N__9034\,
            I => \CLK80_OUT\
        );

    \I__2131\ : CascadeMux
    port map (
            O => \N__9031\,
            I => \N__9024\
        );

    \I__2130\ : InMux
    port map (
            O => \N__9030\,
            I => \N__9013\
        );

    \I__2129\ : InMux
    port map (
            O => \N__9029\,
            I => \N__9013\
        );

    \I__2128\ : InMux
    port map (
            O => \N__9028\,
            I => \N__9010\
        );

    \I__2127\ : InMux
    port map (
            O => \N__9027\,
            I => \N__9005\
        );

    \I__2126\ : InMux
    port map (
            O => \N__9024\,
            I => \N__9005\
        );

    \I__2125\ : InMux
    port map (
            O => \N__9023\,
            I => \N__9002\
        );

    \I__2124\ : InMux
    port map (
            O => \N__9022\,
            I => \N__8997\
        );

    \I__2123\ : InMux
    port map (
            O => \N__9021\,
            I => \N__8997\
        );

    \I__2122\ : InMux
    port map (
            O => \N__9020\,
            I => \N__8994\
        );

    \I__2121\ : InMux
    port map (
            O => \N__9019\,
            I => \N__8991\
        );

    \I__2120\ : InMux
    port map (
            O => \N__9018\,
            I => \N__8988\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__9013\,
            I => \N__8973\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__9010\,
            I => \N__8970\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__9005\,
            I => \N__8962\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__9002\,
            I => \N__8959\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__8997\,
            I => \N__8953\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__8994\,
            I => \N__8948\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__8991\,
            I => \N__8940\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__8988\,
            I => \N__8930\
        );

    \I__2111\ : SRMux
    port map (
            O => \N__8987\,
            I => \N__8842\
        );

    \I__2110\ : SRMux
    port map (
            O => \N__8986\,
            I => \N__8842\
        );

    \I__2109\ : SRMux
    port map (
            O => \N__8985\,
            I => \N__8842\
        );

    \I__2108\ : SRMux
    port map (
            O => \N__8984\,
            I => \N__8842\
        );

    \I__2107\ : SRMux
    port map (
            O => \N__8983\,
            I => \N__8842\
        );

    \I__2106\ : SRMux
    port map (
            O => \N__8982\,
            I => \N__8842\
        );

    \I__2105\ : SRMux
    port map (
            O => \N__8981\,
            I => \N__8842\
        );

    \I__2104\ : SRMux
    port map (
            O => \N__8980\,
            I => \N__8842\
        );

    \I__2103\ : SRMux
    port map (
            O => \N__8979\,
            I => \N__8842\
        );

    \I__2102\ : SRMux
    port map (
            O => \N__8978\,
            I => \N__8842\
        );

    \I__2101\ : SRMux
    port map (
            O => \N__8977\,
            I => \N__8842\
        );

    \I__2100\ : SRMux
    port map (
            O => \N__8976\,
            I => \N__8842\
        );

    \I__2099\ : Glb2LocalMux
    port map (
            O => \N__8973\,
            I => \N__8842\
        );

    \I__2098\ : Glb2LocalMux
    port map (
            O => \N__8970\,
            I => \N__8842\
        );

    \I__2097\ : SRMux
    port map (
            O => \N__8969\,
            I => \N__8842\
        );

    \I__2096\ : SRMux
    port map (
            O => \N__8968\,
            I => \N__8842\
        );

    \I__2095\ : SRMux
    port map (
            O => \N__8967\,
            I => \N__8842\
        );

    \I__2094\ : SRMux
    port map (
            O => \N__8966\,
            I => \N__8842\
        );

    \I__2093\ : SRMux
    port map (
            O => \N__8965\,
            I => \N__8842\
        );

    \I__2092\ : Glb2LocalMux
    port map (
            O => \N__8962\,
            I => \N__8842\
        );

    \I__2091\ : Glb2LocalMux
    port map (
            O => \N__8959\,
            I => \N__8842\
        );

    \I__2090\ : SRMux
    port map (
            O => \N__8958\,
            I => \N__8842\
        );

    \I__2089\ : SRMux
    port map (
            O => \N__8957\,
            I => \N__8842\
        );

    \I__2088\ : SRMux
    port map (
            O => \N__8956\,
            I => \N__8842\
        );

    \I__2087\ : Glb2LocalMux
    port map (
            O => \N__8953\,
            I => \N__8842\
        );

    \I__2086\ : SRMux
    port map (
            O => \N__8952\,
            I => \N__8842\
        );

    \I__2085\ : SRMux
    port map (
            O => \N__8951\,
            I => \N__8842\
        );

    \I__2084\ : Glb2LocalMux
    port map (
            O => \N__8948\,
            I => \N__8842\
        );

    \I__2083\ : SRMux
    port map (
            O => \N__8947\,
            I => \N__8842\
        );

    \I__2082\ : SRMux
    port map (
            O => \N__8946\,
            I => \N__8842\
        );

    \I__2081\ : SRMux
    port map (
            O => \N__8945\,
            I => \N__8842\
        );

    \I__2080\ : SRMux
    port map (
            O => \N__8944\,
            I => \N__8842\
        );

    \I__2079\ : SRMux
    port map (
            O => \N__8943\,
            I => \N__8842\
        );

    \I__2078\ : Glb2LocalMux
    port map (
            O => \N__8940\,
            I => \N__8842\
        );

    \I__2077\ : SRMux
    port map (
            O => \N__8939\,
            I => \N__8842\
        );

    \I__2076\ : SRMux
    port map (
            O => \N__8938\,
            I => \N__8842\
        );

    \I__2075\ : SRMux
    port map (
            O => \N__8937\,
            I => \N__8842\
        );

    \I__2074\ : SRMux
    port map (
            O => \N__8936\,
            I => \N__8842\
        );

    \I__2073\ : SRMux
    port map (
            O => \N__8935\,
            I => \N__8842\
        );

    \I__2072\ : SRMux
    port map (
            O => \N__8934\,
            I => \N__8842\
        );

    \I__2071\ : SRMux
    port map (
            O => \N__8933\,
            I => \N__8842\
        );

    \I__2070\ : Glb2LocalMux
    port map (
            O => \N__8930\,
            I => \N__8842\
        );

    \I__2069\ : SRMux
    port map (
            O => \N__8929\,
            I => \N__8842\
        );

    \I__2068\ : GlobalMux
    port map (
            O => \N__8842\,
            I => \N__8839\
        );

    \I__2067\ : gio2CtrlBuf
    port map (
            O => \N__8839\,
            I => \RESETn_c_i_g\
        );

    \I__2066\ : IoInMux
    port map (
            O => \N__8836\,
            I => \N__8833\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__8833\,
            I => \N__8830\
        );

    \I__2064\ : Span4Mux_s1_v
    port map (
            O => \N__8830\,
            I => \N__8826\
        );

    \I__2063\ : IoInMux
    port map (
            O => \N__8829\,
            I => \N__8823\
        );

    \I__2062\ : Span4Mux_v
    port map (
            O => \N__8826\,
            I => \N__8820\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__8823\,
            I => \N__8817\
        );

    \I__2060\ : Span4Mux_v
    port map (
            O => \N__8820\,
            I => \N__8814\
        );

    \I__2059\ : Span4Mux_s3_h
    port map (
            O => \N__8817\,
            I => \N__8811\
        );

    \I__2058\ : Span4Mux_h
    port map (
            O => \N__8814\,
            I => \N__8808\
        );

    \I__2057\ : Span4Mux_v
    port map (
            O => \N__8811\,
            I => \N__8805\
        );

    \I__2056\ : Odrv4
    port map (
            O => \N__8808\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2055\ : Odrv4
    port map (
            O => \N__8805\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2054\ : InMux
    port map (
            O => \N__8800\,
            I => \N__8797\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__8797\,
            I => \N__8793\
        );

    \I__2052\ : InMux
    port map (
            O => \N__8796\,
            I => \N__8790\
        );

    \I__2051\ : Span4Mux_v
    port map (
            O => \N__8793\,
            I => \N__8787\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__8790\,
            I => \N__8784\
        );

    \I__2049\ : Sp12to4
    port map (
            O => \N__8787\,
            I => \N__8781\
        );

    \I__2048\ : Span12Mux_v
    port map (
            O => \N__8784\,
            I => \N__8778\
        );

    \I__2047\ : Span12Mux_h
    port map (
            O => \N__8781\,
            I => \N__8775\
        );

    \I__2046\ : Span12Mux_h
    port map (
            O => \N__8778\,
            I => \N__8772\
        );

    \I__2045\ : Odrv12
    port map (
            O => \N__8775\,
            I => \DRA_c_7\
        );

    \I__2044\ : Odrv12
    port map (
            O => \N__8772\,
            I => \DRA_c_7\
        );

    \I__2043\ : InMux
    port map (
            O => \N__8767\,
            I => \N__8764\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__8764\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2041\ : InMux
    port map (
            O => \N__8761\,
            I => \N__8758\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__8758\,
            I => \N__8754\
        );

    \I__2039\ : InMux
    port map (
            O => \N__8757\,
            I => \N__8751\
        );

    \I__2038\ : Span4Mux_h
    port map (
            O => \N__8754\,
            I => \N__8746\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__8751\,
            I => \N__8746\
        );

    \I__2036\ : Span4Mux_v
    port map (
            O => \N__8746\,
            I => \N__8743\
        );

    \I__2035\ : Sp12to4
    port map (
            O => \N__8743\,
            I => \N__8740\
        );

    \I__2034\ : Odrv12
    port map (
            O => \N__8740\,
            I => \DRA_c_8\
        );

    \I__2033\ : InMux
    port map (
            O => \N__8737\,
            I => \N__8734\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__8734\,
            I => \N__8731\
        );

    \I__2031\ : Odrv4
    port map (
            O => \N__8731\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__2030\ : CEMux
    port map (
            O => \N__8728\,
            I => \N__8723\
        );

    \I__2029\ : CEMux
    port map (
            O => \N__8727\,
            I => \N__8720\
        );

    \I__2028\ : CEMux
    port map (
            O => \N__8726\,
            I => \N__8717\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__8723\,
            I => \N__8714\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__8720\,
            I => \N__8711\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__8717\,
            I => \N__8708\
        );

    \I__2024\ : Span4Mux_v
    port map (
            O => \N__8714\,
            I => \N__8705\
        );

    \I__2023\ : Span4Mux_h
    port map (
            O => \N__8711\,
            I => \N__8702\
        );

    \I__2022\ : Span4Mux_v
    port map (
            O => \N__8708\,
            I => \N__8699\
        );

    \I__2021\ : Odrv4
    port map (
            O => \N__8705\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__2020\ : Odrv4
    port map (
            O => \N__8702\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__8699\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__2018\ : InMux
    port map (
            O => \N__8692\,
            I => \N__8689\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__8689\,
            I => \N__8685\
        );

    \I__2016\ : InMux
    port map (
            O => \N__8688\,
            I => \N__8682\
        );

    \I__2015\ : Span4Mux_v
    port map (
            O => \N__8685\,
            I => \N__8679\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__8682\,
            I => \N__8676\
        );

    \I__2013\ : Sp12to4
    port map (
            O => \N__8679\,
            I => \N__8673\
        );

    \I__2012\ : Span4Mux_h
    port map (
            O => \N__8676\,
            I => \N__8670\
        );

    \I__2011\ : Span12Mux_h
    port map (
            O => \N__8673\,
            I => \N__8667\
        );

    \I__2010\ : Sp12to4
    port map (
            O => \N__8670\,
            I => \N__8664\
        );

    \I__2009\ : Span12Mux_v
    port map (
            O => \N__8667\,
            I => \N__8661\
        );

    \I__2008\ : Span12Mux_v
    port map (
            O => \N__8664\,
            I => \N__8658\
        );

    \I__2007\ : Odrv12
    port map (
            O => \N__8661\,
            I => \DRA_c_3\
        );

    \I__2006\ : Odrv12
    port map (
            O => \N__8658\,
            I => \DRA_c_3\
        );

    \I__2005\ : InMux
    port map (
            O => \N__8653\,
            I => \N__8650\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__8650\,
            I => \N__8647\
        );

    \I__2003\ : Span4Mux_h
    port map (
            O => \N__8647\,
            I => \N__8644\
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__8644\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__2001\ : CEMux
    port map (
            O => \N__8641\,
            I => \N__8637\
        );

    \I__2000\ : CEMux
    port map (
            O => \N__8640\,
            I => \N__8632\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__8637\,
            I => \N__8629\
        );

    \I__1998\ : CEMux
    port map (
            O => \N__8636\,
            I => \N__8626\
        );

    \I__1997\ : CEMux
    port map (
            O => \N__8635\,
            I => \N__8623\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__8632\,
            I => \N__8619\
        );

    \I__1995\ : Span4Mux_h
    port map (
            O => \N__8629\,
            I => \N__8612\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__8626\,
            I => \N__8612\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__8623\,
            I => \N__8612\
        );

    \I__1992\ : CEMux
    port map (
            O => \N__8622\,
            I => \N__8609\
        );

    \I__1991\ : Span4Mux_h
    port map (
            O => \N__8619\,
            I => \N__8606\
        );

    \I__1990\ : Span4Mux_v
    port map (
            O => \N__8612\,
            I => \N__8603\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__8609\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__1988\ : Odrv4
    port map (
            O => \N__8606\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__1987\ : Odrv4
    port map (
            O => \N__8603\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__1986\ : InMux
    port map (
            O => \N__8596\,
            I => \N__8592\
        );

    \I__1985\ : CascadeMux
    port map (
            O => \N__8595\,
            I => \N__8589\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__8592\,
            I => \N__8580\
        );

    \I__1983\ : InMux
    port map (
            O => \N__8589\,
            I => \N__8577\
        );

    \I__1982\ : CascadeMux
    port map (
            O => \N__8588\,
            I => \N__8572\
        );

    \I__1981\ : CascadeMux
    port map (
            O => \N__8587\,
            I => \N__8569\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__8586\,
            I => \N__8566\
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__8585\,
            I => \N__8563\
        );

    \I__1978\ : InMux
    port map (
            O => \N__8584\,
            I => \N__8556\
        );

    \I__1977\ : InMux
    port map (
            O => \N__8583\,
            I => \N__8556\
        );

    \I__1976\ : Span4Mux_h
    port map (
            O => \N__8580\,
            I => \N__8551\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__8577\,
            I => \N__8551\
        );

    \I__1974\ : InMux
    port map (
            O => \N__8576\,
            I => \N__8546\
        );

    \I__1973\ : InMux
    port map (
            O => \N__8575\,
            I => \N__8546\
        );

    \I__1972\ : InMux
    port map (
            O => \N__8572\,
            I => \N__8543\
        );

    \I__1971\ : InMux
    port map (
            O => \N__8569\,
            I => \N__8540\
        );

    \I__1970\ : InMux
    port map (
            O => \N__8566\,
            I => \N__8534\
        );

    \I__1969\ : InMux
    port map (
            O => \N__8563\,
            I => \N__8531\
        );

    \I__1968\ : CascadeMux
    port map (
            O => \N__8562\,
            I => \N__8528\
        );

    \I__1967\ : CascadeMux
    port map (
            O => \N__8561\,
            I => \N__8525\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__8556\,
            I => \N__8521\
        );

    \I__1965\ : Span4Mux_v
    port map (
            O => \N__8551\,
            I => \N__8518\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__8546\,
            I => \N__8513\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__8543\,
            I => \N__8513\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__8540\,
            I => \N__8510\
        );

    \I__1961\ : InMux
    port map (
            O => \N__8539\,
            I => \N__8503\
        );

    \I__1960\ : InMux
    port map (
            O => \N__8538\,
            I => \N__8503\
        );

    \I__1959\ : InMux
    port map (
            O => \N__8537\,
            I => \N__8503\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__8534\,
            I => \N__8498\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__8531\,
            I => \N__8498\
        );

    \I__1956\ : InMux
    port map (
            O => \N__8528\,
            I => \N__8493\
        );

    \I__1955\ : InMux
    port map (
            O => \N__8525\,
            I => \N__8493\
        );

    \I__1954\ : InMux
    port map (
            O => \N__8524\,
            I => \N__8490\
        );

    \I__1953\ : Span4Mux_v
    port map (
            O => \N__8521\,
            I => \N__8487\
        );

    \I__1952\ : Span4Mux_v
    port map (
            O => \N__8518\,
            I => \N__8484\
        );

    \I__1951\ : Span4Mux_v
    port map (
            O => \N__8513\,
            I => \N__8475\
        );

    \I__1950\ : Span4Mux_h
    port map (
            O => \N__8510\,
            I => \N__8475\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__8503\,
            I => \N__8475\
        );

    \I__1948\ : Span4Mux_h
    port map (
            O => \N__8498\,
            I => \N__8475\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__8493\,
            I => \N__8472\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__8490\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1945\ : Odrv4
    port map (
            O => \N__8487\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1944\ : Odrv4
    port map (
            O => \N__8484\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1943\ : Odrv4
    port map (
            O => \N__8475\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1942\ : Odrv4
    port map (
            O => \N__8472\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1941\ : IoInMux
    port map (
            O => \N__8461\,
            I => \N__8458\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__8458\,
            I => \N__8455\
        );

    \I__1939\ : Span4Mux_s3_v
    port map (
            O => \N__8455\,
            I => \N__8452\
        );

    \I__1938\ : Span4Mux_v
    port map (
            O => \N__8452\,
            I => \N__8449\
        );

    \I__1937\ : Span4Mux_h
    port map (
            O => \N__8449\,
            I => \N__8446\
        );

    \I__1936\ : Odrv4
    port map (
            O => \N__8446\,
            I => \CASn_c\
        );

    \I__1935\ : CascadeMux
    port map (
            O => \N__8443\,
            I => \N__8438\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__8442\,
            I => \N__8432\
        );

    \I__1933\ : InMux
    port map (
            O => \N__8441\,
            I => \N__8427\
        );

    \I__1932\ : InMux
    port map (
            O => \N__8438\,
            I => \N__8420\
        );

    \I__1931\ : InMux
    port map (
            O => \N__8437\,
            I => \N__8420\
        );

    \I__1930\ : CascadeMux
    port map (
            O => \N__8436\,
            I => \N__8416\
        );

    \I__1929\ : InMux
    port map (
            O => \N__8435\,
            I => \N__8413\
        );

    \I__1928\ : InMux
    port map (
            O => \N__8432\,
            I => \N__8410\
        );

    \I__1927\ : InMux
    port map (
            O => \N__8431\,
            I => \N__8405\
        );

    \I__1926\ : InMux
    port map (
            O => \N__8430\,
            I => \N__8405\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__8427\,
            I => \N__8402\
        );

    \I__1924\ : CascadeMux
    port map (
            O => \N__8426\,
            I => \N__8399\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__8425\,
            I => \N__8394\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__8420\,
            I => \N__8391\
        );

    \I__1921\ : InMux
    port map (
            O => \N__8419\,
            I => \N__8386\
        );

    \I__1920\ : InMux
    port map (
            O => \N__8416\,
            I => \N__8386\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__8413\,
            I => \N__8377\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__8410\,
            I => \N__8377\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__8405\,
            I => \N__8377\
        );

    \I__1916\ : Span4Mux_h
    port map (
            O => \N__8402\,
            I => \N__8377\
        );

    \I__1915\ : InMux
    port map (
            O => \N__8399\,
            I => \N__8370\
        );

    \I__1914\ : InMux
    port map (
            O => \N__8398\,
            I => \N__8370\
        );

    \I__1913\ : InMux
    port map (
            O => \N__8397\,
            I => \N__8370\
        );

    \I__1912\ : InMux
    port map (
            O => \N__8394\,
            I => \N__8367\
        );

    \I__1911\ : Span4Mux_v
    port map (
            O => \N__8391\,
            I => \N__8364\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__8386\,
            I => \N__8357\
        );

    \I__1909\ : Sp12to4
    port map (
            O => \N__8377\,
            I => \N__8357\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__8370\,
            I => \N__8357\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__8367\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1906\ : Odrv4
    port map (
            O => \N__8364\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1905\ : Odrv12
    port map (
            O => \N__8357\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1904\ : IoInMux
    port map (
            O => \N__8350\,
            I => \N__8347\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__8347\,
            I => \N__8344\
        );

    \I__1902\ : Span4Mux_s3_h
    port map (
            O => \N__8344\,
            I => \N__8341\
        );

    \I__1901\ : Span4Mux_v
    port map (
            O => \N__8341\,
            I => \N__8338\
        );

    \I__1900\ : Span4Mux_v
    port map (
            O => \N__8338\,
            I => \N__8335\
        );

    \I__1899\ : Span4Mux_h
    port map (
            O => \N__8335\,
            I => \N__8332\
        );

    \I__1898\ : Odrv4
    port map (
            O => \N__8332\,
            I => \WEn_c\
        );

    \I__1897\ : InMux
    port map (
            O => \N__8329\,
            I => \N__8325\
        );

    \I__1896\ : InMux
    port map (
            O => \N__8328\,
            I => \N__8322\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__8325\,
            I => \N__8318\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__8322\,
            I => \N__8315\
        );

    \I__1893\ : InMux
    port map (
            O => \N__8321\,
            I => \N__8312\
        );

    \I__1892\ : Span4Mux_h
    port map (
            O => \N__8318\,
            I => \N__8304\
        );

    \I__1891\ : Span4Mux_h
    port map (
            O => \N__8315\,
            I => \N__8304\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__8312\,
            I => \N__8304\
        );

    \I__1889\ : InMux
    port map (
            O => \N__8311\,
            I => \N__8301\
        );

    \I__1888\ : Odrv4
    port map (
            O => \N__8304\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__8301\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1886\ : IoInMux
    port map (
            O => \N__8296\,
            I => \N__8293\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__8293\,
            I => \N__8290\
        );

    \I__1884\ : Span4Mux_s2_v
    port map (
            O => \N__8290\,
            I => \N__8287\
        );

    \I__1883\ : Span4Mux_v
    port map (
            O => \N__8287\,
            I => \N__8284\
        );

    \I__1882\ : Span4Mux_v
    port map (
            O => \N__8284\,
            I => \N__8281\
        );

    \I__1881\ : Odrv4
    port map (
            O => \N__8281\,
            I => \CRCSn_c\
        );

    \I__1880\ : InMux
    port map (
            O => \N__8278\,
            I => \N__8274\
        );

    \I__1879\ : InMux
    port map (
            O => \N__8277\,
            I => \N__8271\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__8274\,
            I => \N__8268\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__8271\,
            I => \N__8265\
        );

    \I__1876\ : Span4Mux_v
    port map (
            O => \N__8268\,
            I => \N__8262\
        );

    \I__1875\ : Span4Mux_v
    port map (
            O => \N__8265\,
            I => \N__8259\
        );

    \I__1874\ : Sp12to4
    port map (
            O => \N__8262\,
            I => \N__8254\
        );

    \I__1873\ : Sp12to4
    port map (
            O => \N__8259\,
            I => \N__8254\
        );

    \I__1872\ : Span12Mux_h
    port map (
            O => \N__8254\,
            I => \N__8251\
        );

    \I__1871\ : Odrv12
    port map (
            O => \N__8251\,
            I => \RAS0n_c\
        );

    \I__1870\ : InMux
    port map (
            O => \N__8248\,
            I => \N__8245\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__8245\,
            I => \N__8242\
        );

    \I__1868\ : Span12Mux_h
    port map (
            O => \N__8242\,
            I => \N__8239\
        );

    \I__1867\ : Odrv12
    port map (
            O => \N__8239\,
            I => \RAS1n_c\
        );

    \I__1866\ : InMux
    port map (
            O => \N__8236\,
            I => \N__8232\
        );

    \I__1865\ : InMux
    port map (
            O => \N__8235\,
            I => \N__8227\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__8232\,
            I => \N__8221\
        );

    \I__1863\ : InMux
    port map (
            O => \N__8231\,
            I => \N__8218\
        );

    \I__1862\ : InMux
    port map (
            O => \N__8230\,
            I => \N__8215\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__8227\,
            I => \N__8212\
        );

    \I__1860\ : InMux
    port map (
            O => \N__8226\,
            I => \N__8209\
        );

    \I__1859\ : InMux
    port map (
            O => \N__8225\,
            I => \N__8206\
        );

    \I__1858\ : InMux
    port map (
            O => \N__8224\,
            I => \N__8203\
        );

    \I__1857\ : Span4Mux_v
    port map (
            O => \N__8221\,
            I => \N__8198\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__8218\,
            I => \N__8198\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__8215\,
            I => \N__8195\
        );

    \I__1854\ : Span4Mux_v
    port map (
            O => \N__8212\,
            I => \N__8192\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__8209\,
            I => \N__8189\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__8206\,
            I => \N__8184\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__8203\,
            I => \N__8184\
        );

    \I__1850\ : Span4Mux_v
    port map (
            O => \N__8198\,
            I => \N__8179\
        );

    \I__1849\ : Span4Mux_v
    port map (
            O => \N__8195\,
            I => \N__8179\
        );

    \I__1848\ : Span4Mux_h
    port map (
            O => \N__8192\,
            I => \N__8172\
        );

    \I__1847\ : Span4Mux_v
    port map (
            O => \N__8189\,
            I => \N__8172\
        );

    \I__1846\ : Span4Mux_v
    port map (
            O => \N__8184\,
            I => \N__8172\
        );

    \I__1845\ : Sp12to4
    port map (
            O => \N__8179\,
            I => \N__8169\
        );

    \I__1844\ : Sp12to4
    port map (
            O => \N__8172\,
            I => \N__8166\
        );

    \I__1843\ : Span12Mux_h
    port map (
            O => \N__8169\,
            I => \N__8163\
        );

    \I__1842\ : Span12Mux_h
    port map (
            O => \N__8166\,
            I => \N__8160\
        );

    \I__1841\ : Odrv12
    port map (
            O => \N__8163\,
            I => \RESETn_c\
        );

    \I__1840\ : Odrv12
    port map (
            O => \N__8160\,
            I => \RESETn_c\
        );

    \I__1839\ : CascadeMux
    port map (
            O => \N__8155\,
            I => \U712_CHIP_RAM.N_274_cascade_\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__8152\,
            I => \N__8149\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8149\,
            I => \N__8145\
        );

    \I__1836\ : InMux
    port map (
            O => \N__8148\,
            I => \N__8142\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__8145\,
            I => \N__8138\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__8142\,
            I => \N__8135\
        );

    \I__1833\ : InMux
    port map (
            O => \N__8141\,
            I => \N__8132\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__8138\,
            I => \U712_CHIP_RAM.N_337\
        );

    \I__1831\ : Odrv4
    port map (
            O => \N__8135\,
            I => \U712_CHIP_RAM.N_337\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8132\,
            I => \U712_CHIP_RAM.N_337\
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__8125\,
            I => \U712_CHIP_RAM.N_337_cascade_\
        );

    \I__1828\ : InMux
    port map (
            O => \N__8122\,
            I => \N__8119\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8119\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_2_0\
        );

    \I__1826\ : CascadeMux
    port map (
            O => \N__8116\,
            I => \N__8109\
        );

    \I__1825\ : CascadeMux
    port map (
            O => \N__8115\,
            I => \N__8106\
        );

    \I__1824\ : CascadeMux
    port map (
            O => \N__8114\,
            I => \N__8103\
        );

    \I__1823\ : InMux
    port map (
            O => \N__8113\,
            I => \N__8100\
        );

    \I__1822\ : InMux
    port map (
            O => \N__8112\,
            I => \N__8095\
        );

    \I__1821\ : InMux
    port map (
            O => \N__8109\,
            I => \N__8090\
        );

    \I__1820\ : InMux
    port map (
            O => \N__8106\,
            I => \N__8090\
        );

    \I__1819\ : InMux
    port map (
            O => \N__8103\,
            I => \N__8083\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__8100\,
            I => \N__8080\
        );

    \I__1817\ : InMux
    port map (
            O => \N__8099\,
            I => \N__8075\
        );

    \I__1816\ : InMux
    port map (
            O => \N__8098\,
            I => \N__8075\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__8095\,
            I => \N__8072\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__8090\,
            I => \N__8069\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8089\,
            I => \N__8066\
        );

    \I__1812\ : InMux
    port map (
            O => \N__8088\,
            I => \N__8063\
        );

    \I__1811\ : InMux
    port map (
            O => \N__8087\,
            I => \N__8060\
        );

    \I__1810\ : InMux
    port map (
            O => \N__8086\,
            I => \N__8057\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__8083\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1808\ : Odrv4
    port map (
            O => \N__8080\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__8075\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1806\ : Odrv4
    port map (
            O => \N__8072\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1805\ : Odrv4
    port map (
            O => \N__8069\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__8066\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__8063\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__8060\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__8057\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1800\ : InMux
    port map (
            O => \N__8038\,
            I => \N__8031\
        );

    \I__1799\ : InMux
    port map (
            O => \N__8037\,
            I => \N__8028\
        );

    \I__1798\ : InMux
    port map (
            O => \N__8036\,
            I => \N__8021\
        );

    \I__1797\ : InMux
    port map (
            O => \N__8035\,
            I => \N__8021\
        );

    \I__1796\ : InMux
    port map (
            O => \N__8034\,
            I => \N__8021\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__8031\,
            I => \N__8018\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__8028\,
            I => \N__8013\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__8021\,
            I => \N__8008\
        );

    \I__1792\ : Span4Mux_h
    port map (
            O => \N__8018\,
            I => \N__8008\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8017\,
            I => \N__8005\
        );

    \I__1790\ : InMux
    port map (
            O => \N__8016\,
            I => \N__8002\
        );

    \I__1789\ : Odrv4
    port map (
            O => \N__8013\,
            I => \U712_CHIP_RAM.N_271\
        );

    \I__1788\ : Odrv4
    port map (
            O => \N__8008\,
            I => \U712_CHIP_RAM.N_271\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__8005\,
            I => \U712_CHIP_RAM.N_271\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__8002\,
            I => \U712_CHIP_RAM.N_271\
        );

    \I__1785\ : CascadeMux
    port map (
            O => \N__7993\,
            I => \N__7985\
        );

    \I__1784\ : InMux
    port map (
            O => \N__7992\,
            I => \N__7982\
        );

    \I__1783\ : InMux
    port map (
            O => \N__7991\,
            I => \N__7979\
        );

    \I__1782\ : InMux
    port map (
            O => \N__7990\,
            I => \N__7970\
        );

    \I__1781\ : InMux
    port map (
            O => \N__7989\,
            I => \N__7965\
        );

    \I__1780\ : InMux
    port map (
            O => \N__7988\,
            I => \N__7965\
        );

    \I__1779\ : InMux
    port map (
            O => \N__7985\,
            I => \N__7962\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__7982\,
            I => \N__7959\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__7979\,
            I => \N__7956\
        );

    \I__1776\ : InMux
    port map (
            O => \N__7978\,
            I => \N__7951\
        );

    \I__1775\ : InMux
    port map (
            O => \N__7977\,
            I => \N__7951\
        );

    \I__1774\ : InMux
    port map (
            O => \N__7976\,
            I => \N__7948\
        );

    \I__1773\ : InMux
    port map (
            O => \N__7975\,
            I => \N__7945\
        );

    \I__1772\ : InMux
    port map (
            O => \N__7974\,
            I => \N__7940\
        );

    \I__1771\ : InMux
    port map (
            O => \N__7973\,
            I => \N__7940\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__7970\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__7965\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__7962\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1767\ : Odrv12
    port map (
            O => \N__7959\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1766\ : Odrv12
    port map (
            O => \N__7956\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__7951\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__7948\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__7945\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__7940\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1761\ : CascadeMux
    port map (
            O => \N__7921\,
            I => \N__7917\
        );

    \I__1760\ : InMux
    port map (
            O => \N__7920\,
            I => \N__7910\
        );

    \I__1759\ : InMux
    port map (
            O => \N__7917\,
            I => \N__7910\
        );

    \I__1758\ : InMux
    port map (
            O => \N__7916\,
            I => \N__7905\
        );

    \I__1757\ : InMux
    port map (
            O => \N__7915\,
            I => \N__7905\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__7910\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__7905\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1754\ : InMux
    port map (
            O => \N__7900\,
            I => \N__7894\
        );

    \I__1753\ : InMux
    port map (
            O => \N__7899\,
            I => \N__7891\
        );

    \I__1752\ : InMux
    port map (
            O => \N__7898\,
            I => \N__7886\
        );

    \I__1751\ : InMux
    port map (
            O => \N__7897\,
            I => \N__7886\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__7894\,
            I => \N__7883\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__7891\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c3\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__7886\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c3\
        );

    \I__1747\ : Odrv4
    port map (
            O => \N__7883\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c3\
        );

    \I__1746\ : CascadeMux
    port map (
            O => \N__7876\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_5_cascade_\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__7873\,
            I => \N__7870\
        );

    \I__1744\ : InMux
    port map (
            O => \N__7870\,
            I => \N__7866\
        );

    \I__1743\ : InMux
    port map (
            O => \N__7869\,
            I => \N__7863\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__7866\,
            I => \N__7857\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__7863\,
            I => \N__7857\
        );

    \I__1740\ : InMux
    port map (
            O => \N__7862\,
            I => \N__7854\
        );

    \I__1739\ : Odrv4
    port map (
            O => \N__7857\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__7854\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1737\ : CascadeMux
    port map (
            O => \N__7849\,
            I => \N__7843\
        );

    \I__1736\ : CascadeMux
    port map (
            O => \N__7848\,
            I => \N__7840\
        );

    \I__1735\ : InMux
    port map (
            O => \N__7847\,
            I => \N__7833\
        );

    \I__1734\ : InMux
    port map (
            O => \N__7846\,
            I => \N__7833\
        );

    \I__1733\ : InMux
    port map (
            O => \N__7843\,
            I => \N__7828\
        );

    \I__1732\ : InMux
    port map (
            O => \N__7840\,
            I => \N__7828\
        );

    \I__1731\ : CascadeMux
    port map (
            O => \N__7839\,
            I => \N__7824\
        );

    \I__1730\ : CascadeMux
    port map (
            O => \N__7838\,
            I => \N__7820\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__7833\,
            I => \N__7814\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__7828\,
            I => \N__7814\
        );

    \I__1727\ : CascadeMux
    port map (
            O => \N__7827\,
            I => \N__7810\
        );

    \I__1726\ : InMux
    port map (
            O => \N__7824\,
            I => \N__7804\
        );

    \I__1725\ : InMux
    port map (
            O => \N__7823\,
            I => \N__7801\
        );

    \I__1724\ : InMux
    port map (
            O => \N__7820\,
            I => \N__7796\
        );

    \I__1723\ : InMux
    port map (
            O => \N__7819\,
            I => \N__7796\
        );

    \I__1722\ : Span4Mux_h
    port map (
            O => \N__7814\,
            I => \N__7793\
        );

    \I__1721\ : InMux
    port map (
            O => \N__7813\,
            I => \N__7788\
        );

    \I__1720\ : InMux
    port map (
            O => \N__7810\,
            I => \N__7788\
        );

    \I__1719\ : InMux
    port map (
            O => \N__7809\,
            I => \N__7785\
        );

    \I__1718\ : InMux
    port map (
            O => \N__7808\,
            I => \N__7780\
        );

    \I__1717\ : InMux
    port map (
            O => \N__7807\,
            I => \N__7780\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__7804\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__7801\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__7796\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1713\ : Odrv4
    port map (
            O => \N__7793\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__7788\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__7785\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__7780\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1709\ : InMux
    port map (
            O => \N__7765\,
            I => \N__7762\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__7762\,
            I => \N__7758\
        );

    \I__1707\ : InMux
    port map (
            O => \N__7761\,
            I => \N__7754\
        );

    \I__1706\ : Span4Mux_v
    port map (
            O => \N__7758\,
            I => \N__7751\
        );

    \I__1705\ : InMux
    port map (
            O => \N__7757\,
            I => \N__7748\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__7754\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER46\
        );

    \I__1703\ : Odrv4
    port map (
            O => \N__7751\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER46\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__7748\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER46\
        );

    \I__1701\ : CascadeMux
    port map (
            O => \N__7741\,
            I => \N__7736\
        );

    \I__1700\ : CascadeMux
    port map (
            O => \N__7740\,
            I => \N__7727\
        );

    \I__1699\ : InMux
    port map (
            O => \N__7739\,
            I => \N__7723\
        );

    \I__1698\ : InMux
    port map (
            O => \N__7736\,
            I => \N__7717\
        );

    \I__1697\ : CascadeMux
    port map (
            O => \N__7735\,
            I => \N__7713\
        );

    \I__1696\ : InMux
    port map (
            O => \N__7734\,
            I => \N__7710\
        );

    \I__1695\ : InMux
    port map (
            O => \N__7733\,
            I => \N__7703\
        );

    \I__1694\ : InMux
    port map (
            O => \N__7732\,
            I => \N__7703\
        );

    \I__1693\ : InMux
    port map (
            O => \N__7731\,
            I => \N__7703\
        );

    \I__1692\ : CascadeMux
    port map (
            O => \N__7730\,
            I => \N__7691\
        );

    \I__1691\ : InMux
    port map (
            O => \N__7727\,
            I => \N__7688\
        );

    \I__1690\ : InMux
    port map (
            O => \N__7726\,
            I => \N__7685\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__7723\,
            I => \N__7682\
        );

    \I__1688\ : InMux
    port map (
            O => \N__7722\,
            I => \N__7679\
        );

    \I__1687\ : InMux
    port map (
            O => \N__7721\,
            I => \N__7674\
        );

    \I__1686\ : InMux
    port map (
            O => \N__7720\,
            I => \N__7674\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__7717\,
            I => \N__7671\
        );

    \I__1684\ : InMux
    port map (
            O => \N__7716\,
            I => \N__7668\
        );

    \I__1683\ : InMux
    port map (
            O => \N__7713\,
            I => \N__7665\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__7710\,
            I => \N__7662\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__7703\,
            I => \N__7659\
        );

    \I__1680\ : InMux
    port map (
            O => \N__7702\,
            I => \N__7652\
        );

    \I__1679\ : InMux
    port map (
            O => \N__7701\,
            I => \N__7652\
        );

    \I__1678\ : InMux
    port map (
            O => \N__7700\,
            I => \N__7652\
        );

    \I__1677\ : InMux
    port map (
            O => \N__7699\,
            I => \N__7649\
        );

    \I__1676\ : InMux
    port map (
            O => \N__7698\,
            I => \N__7644\
        );

    \I__1675\ : InMux
    port map (
            O => \N__7697\,
            I => \N__7644\
        );

    \I__1674\ : InMux
    port map (
            O => \N__7696\,
            I => \N__7641\
        );

    \I__1673\ : InMux
    port map (
            O => \N__7695\,
            I => \N__7636\
        );

    \I__1672\ : InMux
    port map (
            O => \N__7694\,
            I => \N__7636\
        );

    \I__1671\ : InMux
    port map (
            O => \N__7691\,
            I => \N__7633\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__7688\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__7685\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1668\ : Odrv4
    port map (
            O => \N__7682\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__7679\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__7674\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1665\ : Odrv4
    port map (
            O => \N__7671\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__7668\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__7665\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1662\ : Odrv4
    port map (
            O => \N__7662\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1661\ : Odrv4
    port map (
            O => \N__7659\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__7652\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__7649\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__7644\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__7641\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__7636\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__7633\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1654\ : InMux
    port map (
            O => \N__7600\,
            I => \N__7596\
        );

    \I__1653\ : InMux
    port map (
            O => \N__7599\,
            I => \N__7593\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__7596\,
            I => \N__7590\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__7593\,
            I => \U712_CHIP_RAM.N_303\
        );

    \I__1650\ : Odrv4
    port map (
            O => \N__7590\,
            I => \U712_CHIP_RAM.N_303\
        );

    \I__1649\ : InMux
    port map (
            O => \N__7585\,
            I => \N__7576\
        );

    \I__1648\ : InMux
    port map (
            O => \N__7584\,
            I => \N__7573\
        );

    \I__1647\ : InMux
    port map (
            O => \N__7583\,
            I => \N__7567\
        );

    \I__1646\ : InMux
    port map (
            O => \N__7582\,
            I => \N__7567\
        );

    \I__1645\ : InMux
    port map (
            O => \N__7581\,
            I => \N__7564\
        );

    \I__1644\ : InMux
    port map (
            O => \N__7580\,
            I => \N__7561\
        );

    \I__1643\ : InMux
    port map (
            O => \N__7579\,
            I => \N__7558\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__7576\,
            I => \N__7555\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__7573\,
            I => \N__7552\
        );

    \I__1640\ : InMux
    port map (
            O => \N__7572\,
            I => \N__7549\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__7567\,
            I => \N__7546\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__7564\,
            I => \N__7538\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__7561\,
            I => \N__7538\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__7558\,
            I => \N__7538\
        );

    \I__1635\ : Span4Mux_v
    port map (
            O => \N__7555\,
            I => \N__7531\
        );

    \I__1634\ : Span4Mux_v
    port map (
            O => \N__7552\,
            I => \N__7531\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__7549\,
            I => \N__7531\
        );

    \I__1632\ : Span4Mux_v
    port map (
            O => \N__7546\,
            I => \N__7528\
        );

    \I__1631\ : InMux
    port map (
            O => \N__7545\,
            I => \N__7525\
        );

    \I__1630\ : Span4Mux_v
    port map (
            O => \N__7538\,
            I => \N__7520\
        );

    \I__1629\ : Span4Mux_h
    port map (
            O => \N__7531\,
            I => \N__7520\
        );

    \I__1628\ : Odrv4
    port map (
            O => \N__7528\,
            I => \DMA_CYCLEm\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__7525\,
            I => \DMA_CYCLEm\
        );

    \I__1626\ : Odrv4
    port map (
            O => \N__7520\,
            I => \DMA_CYCLEm\
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__7513\,
            I => \N__7509\
        );

    \I__1624\ : InMux
    port map (
            O => \N__7512\,
            I => \N__7506\
        );

    \I__1623\ : InMux
    port map (
            O => \N__7509\,
            I => \N__7503\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__7506\,
            I => \N__7500\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__7503\,
            I => \N__7497\
        );

    \I__1620\ : Span4Mux_v
    port map (
            O => \N__7500\,
            I => \N__7493\
        );

    \I__1619\ : Span4Mux_v
    port map (
            O => \N__7497\,
            I => \N__7490\
        );

    \I__1618\ : InMux
    port map (
            O => \N__7496\,
            I => \N__7487\
        );

    \I__1617\ : Sp12to4
    port map (
            O => \N__7493\,
            I => \N__7481\
        );

    \I__1616\ : Sp12to4
    port map (
            O => \N__7490\,
            I => \N__7481\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__7487\,
            I => \N__7478\
        );

    \I__1614\ : InMux
    port map (
            O => \N__7486\,
            I => \N__7475\
        );

    \I__1613\ : Odrv12
    port map (
            O => \N__7481\,
            I => \REG_CYCLEm\
        );

    \I__1612\ : Odrv12
    port map (
            O => \N__7478\,
            I => \REG_CYCLEm\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__7475\,
            I => \REG_CYCLEm\
        );

    \I__1610\ : IoInMux
    port map (
            O => \N__7468\,
            I => \N__7465\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__7465\,
            I => \N__7462\
        );

    \I__1608\ : Span12Mux_s4_v
    port map (
            O => \N__7462\,
            I => \N__7459\
        );

    \I__1607\ : Span12Mux_h
    port map (
            O => \N__7459\,
            I => \N__7456\
        );

    \I__1606\ : Odrv12
    port map (
            O => \N__7456\,
            I => \DRDENn_c\
        );

    \I__1605\ : CascadeMux
    port map (
            O => \N__7453\,
            I => \N__7450\
        );

    \I__1604\ : InMux
    port map (
            O => \N__7450\,
            I => \N__7447\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__7447\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__1602\ : CascadeMux
    port map (
            O => \N__7444\,
            I => \U712_CHIP_RAM.N_284_cascade_\
        );

    \I__1601\ : InMux
    port map (
            O => \N__7441\,
            I => \N__7438\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__7438\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_1_2\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7435\,
            I => \N__7432\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__7432\,
            I => \N__7429\
        );

    \I__1597\ : Odrv12
    port map (
            O => \N__7429\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1596\ : CascadeMux
    port map (
            O => \N__7426\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_1_0_cascade_\
        );

    \I__1595\ : InMux
    port map (
            O => \N__7423\,
            I => \N__7420\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__7420\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_0\
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__7417\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c6_cascade_\
        );

    \I__1592\ : InMux
    port map (
            O => \N__7414\,
            I => \N__7400\
        );

    \I__1591\ : InMux
    port map (
            O => \N__7413\,
            I => \N__7400\
        );

    \I__1590\ : InMux
    port map (
            O => \N__7412\,
            I => \N__7400\
        );

    \I__1589\ : InMux
    port map (
            O => \N__7411\,
            I => \N__7393\
        );

    \I__1588\ : InMux
    port map (
            O => \N__7410\,
            I => \N__7393\
        );

    \I__1587\ : InMux
    port map (
            O => \N__7409\,
            I => \N__7393\
        );

    \I__1586\ : InMux
    port map (
            O => \N__7408\,
            I => \N__7390\
        );

    \I__1585\ : CascadeMux
    port map (
            O => \N__7407\,
            I => \N__7385\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__7400\,
            I => \N__7378\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__7393\,
            I => \N__7375\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__7390\,
            I => \N__7367\
        );

    \I__1581\ : InMux
    port map (
            O => \N__7389\,
            I => \N__7362\
        );

    \I__1580\ : InMux
    port map (
            O => \N__7388\,
            I => \N__7362\
        );

    \I__1579\ : InMux
    port map (
            O => \N__7385\,
            I => \N__7355\
        );

    \I__1578\ : InMux
    port map (
            O => \N__7384\,
            I => \N__7352\
        );

    \I__1577\ : InMux
    port map (
            O => \N__7383\,
            I => \N__7345\
        );

    \I__1576\ : InMux
    port map (
            O => \N__7382\,
            I => \N__7345\
        );

    \I__1575\ : InMux
    port map (
            O => \N__7381\,
            I => \N__7345\
        );

    \I__1574\ : Span4Mux_h
    port map (
            O => \N__7378\,
            I => \N__7342\
        );

    \I__1573\ : Span4Mux_h
    port map (
            O => \N__7375\,
            I => \N__7339\
        );

    \I__1572\ : InMux
    port map (
            O => \N__7374\,
            I => \N__7330\
        );

    \I__1571\ : InMux
    port map (
            O => \N__7373\,
            I => \N__7330\
        );

    \I__1570\ : InMux
    port map (
            O => \N__7372\,
            I => \N__7330\
        );

    \I__1569\ : InMux
    port map (
            O => \N__7371\,
            I => \N__7330\
        );

    \I__1568\ : InMux
    port map (
            O => \N__7370\,
            I => \N__7327\
        );

    \I__1567\ : Span4Mux_h
    port map (
            O => \N__7367\,
            I => \N__7322\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__7362\,
            I => \N__7322\
        );

    \I__1565\ : InMux
    port map (
            O => \N__7361\,
            I => \N__7317\
        );

    \I__1564\ : InMux
    port map (
            O => \N__7360\,
            I => \N__7317\
        );

    \I__1563\ : InMux
    port map (
            O => \N__7359\,
            I => \N__7314\
        );

    \I__1562\ : InMux
    port map (
            O => \N__7358\,
            I => \N__7311\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__7355\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__7352\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__7345\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1558\ : Odrv4
    port map (
            O => \N__7342\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1557\ : Odrv4
    port map (
            O => \N__7339\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__7330\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__7327\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1554\ : Odrv4
    port map (
            O => \N__7322\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__7317\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__7314\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__7311\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1550\ : InMux
    port map (
            O => \N__7288\,
            I => \N__7285\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__7285\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_0_3\
        );

    \I__1548\ : CascadeMux
    port map (
            O => \N__7282\,
            I => \N__7279\
        );

    \I__1547\ : InMux
    port map (
            O => \N__7279\,
            I => \N__7276\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__7276\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c6\
        );

    \I__1545\ : InMux
    port map (
            O => \N__7273\,
            I => \N__7268\
        );

    \I__1544\ : InMux
    port map (
            O => \N__7272\,
            I => \N__7263\
        );

    \I__1543\ : InMux
    port map (
            O => \N__7271\,
            I => \N__7263\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__7268\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__7263\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1540\ : CascadeMux
    port map (
            O => \N__7258\,
            I => \N__7254\
        );

    \I__1539\ : InMux
    port map (
            O => \N__7257\,
            I => \N__7249\
        );

    \I__1538\ : InMux
    port map (
            O => \N__7254\,
            I => \N__7249\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__7249\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1536\ : InMux
    port map (
            O => \N__7246\,
            I => \N__7241\
        );

    \I__1535\ : InMux
    port map (
            O => \N__7245\,
            I => \N__7231\
        );

    \I__1534\ : InMux
    port map (
            O => \N__7244\,
            I => \N__7231\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__7241\,
            I => \N__7228\
        );

    \I__1532\ : InMux
    port map (
            O => \N__7240\,
            I => \N__7225\
        );

    \I__1531\ : CascadeMux
    port map (
            O => \N__7239\,
            I => \N__7222\
        );

    \I__1530\ : InMux
    port map (
            O => \N__7238\,
            I => \N__7218\
        );

    \I__1529\ : InMux
    port map (
            O => \N__7237\,
            I => \N__7215\
        );

    \I__1528\ : InMux
    port map (
            O => \N__7236\,
            I => \N__7212\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7231\,
            I => \N__7209\
        );

    \I__1526\ : Span4Mux_v
    port map (
            O => \N__7228\,
            I => \N__7204\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__7225\,
            I => \N__7204\
        );

    \I__1524\ : InMux
    port map (
            O => \N__7222\,
            I => \N__7201\
        );

    \I__1523\ : InMux
    port map (
            O => \N__7221\,
            I => \N__7198\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__7218\,
            I => \U712_CHIP_RAM.N_274\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__7215\,
            I => \U712_CHIP_RAM.N_274\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__7212\,
            I => \U712_CHIP_RAM.N_274\
        );

    \I__1519\ : Odrv4
    port map (
            O => \N__7209\,
            I => \U712_CHIP_RAM.N_274\
        );

    \I__1518\ : Odrv4
    port map (
            O => \N__7204\,
            I => \U712_CHIP_RAM.N_274\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__7201\,
            I => \U712_CHIP_RAM.N_274\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__7198\,
            I => \U712_CHIP_RAM.N_274\
        );

    \I__1515\ : InMux
    port map (
            O => \N__7183\,
            I => \N__7180\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__7180\,
            I => \N__7177\
        );

    \I__1513\ : Sp12to4
    port map (
            O => \N__7177\,
            I => \N__7174\
        );

    \I__1512\ : Span12Mux_v
    port map (
            O => \N__7174\,
            I => \N__7171\
        );

    \I__1511\ : Span12Mux_h
    port map (
            O => \N__7171\,
            I => \N__7168\
        );

    \I__1510\ : Odrv12
    port map (
            O => \N__7168\,
            I => \A_c_17\
        );

    \I__1509\ : InMux
    port map (
            O => \N__7165\,
            I => \N__7162\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__7162\,
            I => \N__7159\
        );

    \I__1507\ : Odrv4
    port map (
            O => \N__7159\,
            I => \U712_CHIP_RAM.CMA_5_i_0_8\
        );

    \I__1506\ : IoInMux
    port map (
            O => \N__7156\,
            I => \N__7153\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__7153\,
            I => \N__7150\
        );

    \I__1504\ : IoSpan4Mux
    port map (
            O => \N__7150\,
            I => \N__7147\
        );

    \I__1503\ : Span4Mux_s0_h
    port map (
            O => \N__7147\,
            I => \N__7144\
        );

    \I__1502\ : Sp12to4
    port map (
            O => \N__7144\,
            I => \N__7141\
        );

    \I__1501\ : Span12Mux_h
    port map (
            O => \N__7141\,
            I => \N__7138\
        );

    \I__1500\ : Odrv12
    port map (
            O => \N__7138\,
            I => \CMA_c_8\
        );

    \I__1499\ : InMux
    port map (
            O => \N__7135\,
            I => \N__7132\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__7132\,
            I => \U712_CHIP_RAM.N_318\
        );

    \I__1497\ : IoInMux
    port map (
            O => \N__7129\,
            I => \N__7126\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__7126\,
            I => \N__7123\
        );

    \I__1495\ : Span4Mux_s2_h
    port map (
            O => \N__7123\,
            I => \N__7120\
        );

    \I__1494\ : Span4Mux_v
    port map (
            O => \N__7120\,
            I => \N__7117\
        );

    \I__1493\ : Sp12to4
    port map (
            O => \N__7117\,
            I => \N__7114\
        );

    \I__1492\ : Span12Mux_h
    port map (
            O => \N__7114\,
            I => \N__7111\
        );

    \I__1491\ : Odrv12
    port map (
            O => \N__7111\,
            I => \CMA_c_7\
        );

    \I__1490\ : CascadeMux
    port map (
            O => \N__7108\,
            I => \N__7104\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7107\,
            I => \N__7096\
        );

    \I__1488\ : InMux
    port map (
            O => \N__7104\,
            I => \N__7089\
        );

    \I__1487\ : InMux
    port map (
            O => \N__7103\,
            I => \N__7089\
        );

    \I__1486\ : InMux
    port map (
            O => \N__7102\,
            I => \N__7084\
        );

    \I__1485\ : InMux
    port map (
            O => \N__7101\,
            I => \N__7084\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7100\,
            I => \N__7081\
        );

    \I__1483\ : InMux
    port map (
            O => \N__7099\,
            I => \N__7078\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__7096\,
            I => \N__7070\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7095\,
            I => \N__7065\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7094\,
            I => \N__7065\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__7089\,
            I => \N__7060\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__7084\,
            I => \N__7060\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__7081\,
            I => \N__7055\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__7078\,
            I => \N__7055\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7077\,
            I => \N__7052\
        );

    \I__1474\ : InMux
    port map (
            O => \N__7076\,
            I => \N__7045\
        );

    \I__1473\ : InMux
    port map (
            O => \N__7075\,
            I => \N__7045\
        );

    \I__1472\ : InMux
    port map (
            O => \N__7074\,
            I => \N__7045\
        );

    \I__1471\ : InMux
    port map (
            O => \N__7073\,
            I => \N__7042\
        );

    \I__1470\ : Span4Mux_v
    port map (
            O => \N__7070\,
            I => \N__7039\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__7065\,
            I => \N__7028\
        );

    \I__1468\ : Span4Mux_h
    port map (
            O => \N__7060\,
            I => \N__7028\
        );

    \I__1467\ : Span4Mux_v
    port map (
            O => \N__7055\,
            I => \N__7028\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7052\,
            I => \N__7028\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__7045\,
            I => \N__7028\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__7042\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1463\ : Odrv4
    port map (
            O => \N__7039\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1462\ : Odrv4
    port map (
            O => \N__7028\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1461\ : InMux
    port map (
            O => \N__7021\,
            I => \N__7018\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__7018\,
            I => \N__7015\
        );

    \I__1459\ : Odrv4
    port map (
            O => \N__7015\,
            I => \U712_CHIP_RAM.N_315\
        );

    \I__1458\ : IoInMux
    port map (
            O => \N__7012\,
            I => \N__7009\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__7009\,
            I => \N__7006\
        );

    \I__1456\ : Span4Mux_s3_h
    port map (
            O => \N__7006\,
            I => \N__7003\
        );

    \I__1455\ : Sp12to4
    port map (
            O => \N__7003\,
            I => \N__7000\
        );

    \I__1454\ : Span12Mux_s10_v
    port map (
            O => \N__7000\,
            I => \N__6997\
        );

    \I__1453\ : Odrv12
    port map (
            O => \N__6997\,
            I => \CMA_c_4\
        );

    \I__1452\ : CEMux
    port map (
            O => \N__6994\,
            I => \N__6990\
        );

    \I__1451\ : CEMux
    port map (
            O => \N__6993\,
            I => \N__6986\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__6990\,
            I => \N__6982\
        );

    \I__1449\ : CEMux
    port map (
            O => \N__6989\,
            I => \N__6979\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__6986\,
            I => \N__6975\
        );

    \I__1447\ : CEMux
    port map (
            O => \N__6985\,
            I => \N__6972\
        );

    \I__1446\ : Span4Mux_v
    port map (
            O => \N__6982\,
            I => \N__6968\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__6979\,
            I => \N__6965\
        );

    \I__1444\ : CEMux
    port map (
            O => \N__6978\,
            I => \N__6962\
        );

    \I__1443\ : Span4Mux_v
    port map (
            O => \N__6975\,
            I => \N__6957\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__6972\,
            I => \N__6957\
        );

    \I__1441\ : CEMux
    port map (
            O => \N__6971\,
            I => \N__6954\
        );

    \I__1440\ : Span4Mux_h
    port map (
            O => \N__6968\,
            I => \N__6951\
        );

    \I__1439\ : Span4Mux_v
    port map (
            O => \N__6965\,
            I => \N__6948\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__6962\,
            I => \N__6945\
        );

    \I__1437\ : Span4Mux_v
    port map (
            O => \N__6957\,
            I => \N__6942\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__6954\,
            I => \N__6939\
        );

    \I__1435\ : Odrv4
    port map (
            O => \N__6951\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1434\ : Odrv4
    port map (
            O => \N__6948\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1433\ : Odrv4
    port map (
            O => \N__6945\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1432\ : Odrv4
    port map (
            O => \N__6942\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1431\ : Odrv4
    port map (
            O => \N__6939\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1430\ : InMux
    port map (
            O => \N__6928\,
            I => \N__6924\
        );

    \I__1429\ : InMux
    port map (
            O => \N__6927\,
            I => \N__6921\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__6924\,
            I => \N__6918\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__6921\,
            I => \N__6915\
        );

    \I__1426\ : Span4Mux_v
    port map (
            O => \N__6918\,
            I => \N__6912\
        );

    \I__1425\ : Sp12to4
    port map (
            O => \N__6915\,
            I => \N__6909\
        );

    \I__1424\ : Sp12to4
    port map (
            O => \N__6912\,
            I => \N__6906\
        );

    \I__1423\ : Span12Mux_v
    port map (
            O => \N__6909\,
            I => \N__6903\
        );

    \I__1422\ : Span12Mux_h
    port map (
            O => \N__6906\,
            I => \N__6900\
        );

    \I__1421\ : Span12Mux_h
    port map (
            O => \N__6903\,
            I => \N__6897\
        );

    \I__1420\ : Span12Mux_v
    port map (
            O => \N__6900\,
            I => \N__6894\
        );

    \I__1419\ : Odrv12
    port map (
            O => \N__6897\,
            I => \AWEn_c\
        );

    \I__1418\ : Odrv12
    port map (
            O => \N__6894\,
            I => \AWEn_c\
        );

    \I__1417\ : CascadeMux
    port map (
            O => \N__6889\,
            I => \N__6886\
        );

    \I__1416\ : InMux
    port map (
            O => \N__6886\,
            I => \N__6883\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__6883\,
            I => \N__6880\
        );

    \I__1414\ : Span4Mux_v
    port map (
            O => \N__6880\,
            I => \N__6875\
        );

    \I__1413\ : InMux
    port map (
            O => \N__6879\,
            I => \N__6871\
        );

    \I__1412\ : InMux
    port map (
            O => \N__6878\,
            I => \N__6868\
        );

    \I__1411\ : Span4Mux_v
    port map (
            O => \N__6875\,
            I => \N__6865\
        );

    \I__1410\ : InMux
    port map (
            O => \N__6874\,
            I => \N__6862\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__6871\,
            I => \N__6859\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__6868\,
            I => \N__6856\
        );

    \I__1407\ : Span4Mux_h
    port map (
            O => \N__6865\,
            I => \N__6853\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__6862\,
            I => \N__6850\
        );

    \I__1405\ : Span4Mux_v
    port map (
            O => \N__6859\,
            I => \N__6847\
        );

    \I__1404\ : Span4Mux_v
    port map (
            O => \N__6856\,
            I => \N__6844\
        );

    \I__1403\ : Sp12to4
    port map (
            O => \N__6853\,
            I => \N__6835\
        );

    \I__1402\ : Span12Mux_h
    port map (
            O => \N__6850\,
            I => \N__6835\
        );

    \I__1401\ : Sp12to4
    port map (
            O => \N__6847\,
            I => \N__6835\
        );

    \I__1400\ : Sp12to4
    port map (
            O => \N__6844\,
            I => \N__6835\
        );

    \I__1399\ : Span12Mux_h
    port map (
            O => \N__6835\,
            I => \N__6832\
        );

    \I__1398\ : Span12Mux_v
    port map (
            O => \N__6832\,
            I => \N__6829\
        );

    \I__1397\ : Odrv12
    port map (
            O => \N__6829\,
            I => \RnW_c\
        );

    \I__1396\ : InMux
    port map (
            O => \N__6826\,
            I => \N__6817\
        );

    \I__1395\ : InMux
    port map (
            O => \N__6825\,
            I => \N__6806\
        );

    \I__1394\ : InMux
    port map (
            O => \N__6824\,
            I => \N__6801\
        );

    \I__1393\ : InMux
    port map (
            O => \N__6823\,
            I => \N__6801\
        );

    \I__1392\ : InMux
    port map (
            O => \N__6822\,
            I => \N__6798\
        );

    \I__1391\ : InMux
    port map (
            O => \N__6821\,
            I => \N__6793\
        );

    \I__1390\ : InMux
    port map (
            O => \N__6820\,
            I => \N__6793\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__6817\,
            I => \N__6787\
        );

    \I__1388\ : InMux
    port map (
            O => \N__6816\,
            I => \N__6782\
        );

    \I__1387\ : InMux
    port map (
            O => \N__6815\,
            I => \N__6782\
        );

    \I__1386\ : CascadeMux
    port map (
            O => \N__6814\,
            I => \N__6777\
        );

    \I__1385\ : InMux
    port map (
            O => \N__6813\,
            I => \N__6770\
        );

    \I__1384\ : InMux
    port map (
            O => \N__6812\,
            I => \N__6767\
        );

    \I__1383\ : InMux
    port map (
            O => \N__6811\,
            I => \N__6764\
        );

    \I__1382\ : InMux
    port map (
            O => \N__6810\,
            I => \N__6759\
        );

    \I__1381\ : InMux
    port map (
            O => \N__6809\,
            I => \N__6759\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__6806\,
            I => \N__6754\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__6801\,
            I => \N__6754\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__6798\,
            I => \N__6749\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__6793\,
            I => \N__6749\
        );

    \I__1376\ : InMux
    port map (
            O => \N__6792\,
            I => \N__6744\
        );

    \I__1375\ : InMux
    port map (
            O => \N__6791\,
            I => \N__6740\
        );

    \I__1374\ : InMux
    port map (
            O => \N__6790\,
            I => \N__6737\
        );

    \I__1373\ : Span4Mux_h
    port map (
            O => \N__6787\,
            I => \N__6732\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__6782\,
            I => \N__6732\
        );

    \I__1371\ : InMux
    port map (
            O => \N__6781\,
            I => \N__6723\
        );

    \I__1370\ : InMux
    port map (
            O => \N__6780\,
            I => \N__6723\
        );

    \I__1369\ : InMux
    port map (
            O => \N__6777\,
            I => \N__6723\
        );

    \I__1368\ : InMux
    port map (
            O => \N__6776\,
            I => \N__6723\
        );

    \I__1367\ : CascadeMux
    port map (
            O => \N__6775\,
            I => \N__6720\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__6774\,
            I => \N__6717\
        );

    \I__1365\ : CascadeMux
    port map (
            O => \N__6773\,
            I => \N__6714\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__6770\,
            I => \N__6711\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__6767\,
            I => \N__6706\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__6764\,
            I => \N__6706\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__6759\,
            I => \N__6701\
        );

    \I__1360\ : Span4Mux_h
    port map (
            O => \N__6754\,
            I => \N__6701\
        );

    \I__1359\ : Span4Mux_v
    port map (
            O => \N__6749\,
            I => \N__6698\
        );

    \I__1358\ : InMux
    port map (
            O => \N__6748\,
            I => \N__6695\
        );

    \I__1357\ : InMux
    port map (
            O => \N__6747\,
            I => \N__6692\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__6744\,
            I => \N__6689\
        );

    \I__1355\ : InMux
    port map (
            O => \N__6743\,
            I => \N__6686\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__6740\,
            I => \N__6683\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__6737\,
            I => \N__6676\
        );

    \I__1352\ : Sp12to4
    port map (
            O => \N__6732\,
            I => \N__6676\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__6723\,
            I => \N__6676\
        );

    \I__1350\ : InMux
    port map (
            O => \N__6720\,
            I => \N__6669\
        );

    \I__1349\ : InMux
    port map (
            O => \N__6717\,
            I => \N__6669\
        );

    \I__1348\ : InMux
    port map (
            O => \N__6714\,
            I => \N__6669\
        );

    \I__1347\ : Span4Mux_v
    port map (
            O => \N__6711\,
            I => \N__6662\
        );

    \I__1346\ : Span4Mux_v
    port map (
            O => \N__6706\,
            I => \N__6662\
        );

    \I__1345\ : Span4Mux_v
    port map (
            O => \N__6701\,
            I => \N__6662\
        );

    \I__1344\ : Odrv4
    port map (
            O => \N__6698\,
            I => \CPU_CYCLEm\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__6695\,
            I => \CPU_CYCLEm\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__6692\,
            I => \CPU_CYCLEm\
        );

    \I__1341\ : Odrv4
    port map (
            O => \N__6689\,
            I => \CPU_CYCLEm\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__6686\,
            I => \CPU_CYCLEm\
        );

    \I__1339\ : Odrv4
    port map (
            O => \N__6683\,
            I => \CPU_CYCLEm\
        );

    \I__1338\ : Odrv12
    port map (
            O => \N__6676\,
            I => \CPU_CYCLEm\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__6669\,
            I => \CPU_CYCLEm\
        );

    \I__1336\ : Odrv4
    port map (
            O => \N__6662\,
            I => \CPU_CYCLEm\
        );

    \I__1335\ : CEMux
    port map (
            O => \N__6643\,
            I => \N__6640\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__6640\,
            I => \N__6637\
        );

    \I__1333\ : Odrv4
    port map (
            O => \N__6637\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_0\
        );

    \I__1332\ : InMux
    port map (
            O => \N__6634\,
            I => \N__6631\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__6631\,
            I => \N__6626\
        );

    \I__1330\ : CascadeMux
    port map (
            O => \N__6630\,
            I => \N__6621\
        );

    \I__1329\ : InMux
    port map (
            O => \N__6629\,
            I => \N__6616\
        );

    \I__1328\ : Span4Mux_v
    port map (
            O => \N__6626\,
            I => \N__6613\
        );

    \I__1327\ : InMux
    port map (
            O => \N__6625\,
            I => \N__6608\
        );

    \I__1326\ : InMux
    port map (
            O => \N__6624\,
            I => \N__6608\
        );

    \I__1325\ : InMux
    port map (
            O => \N__6621\,
            I => \N__6601\
        );

    \I__1324\ : InMux
    port map (
            O => \N__6620\,
            I => \N__6601\
        );

    \I__1323\ : InMux
    port map (
            O => \N__6619\,
            I => \N__6601\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__6616\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1321\ : Odrv4
    port map (
            O => \N__6613\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__6608\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__6601\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1318\ : CEMux
    port map (
            O => \N__6592\,
            I => \N__6589\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__6589\,
            I => \N__6586\
        );

    \I__1316\ : Span4Mux_v
    port map (
            O => \N__6586\,
            I => \N__6583\
        );

    \I__1315\ : Span4Mux_h
    port map (
            O => \N__6583\,
            I => \N__6580\
        );

    \I__1314\ : Odrv4
    port map (
            O => \N__6580\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_0\
        );

    \I__1313\ : CEMux
    port map (
            O => \N__6577\,
            I => \N__6574\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__6574\,
            I => \N__6571\
        );

    \I__1311\ : Span4Mux_v
    port map (
            O => \N__6571\,
            I => \N__6568\
        );

    \I__1310\ : Span4Mux_h
    port map (
            O => \N__6568\,
            I => \N__6565\
        );

    \I__1309\ : Odrv4
    port map (
            O => \N__6565\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0\
        );

    \I__1308\ : InMux
    port map (
            O => \N__6562\,
            I => \N__6559\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__6559\,
            I => \N__6556\
        );

    \I__1306\ : Odrv4
    port map (
            O => \N__6556\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_i_a2_1_0_a2_1_0\
        );

    \I__1305\ : InMux
    port map (
            O => \N__6553\,
            I => \N__6550\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__6550\,
            I => \U712_CHIP_RAM.N_284\
        );

    \I__1303\ : InMux
    port map (
            O => \N__6547\,
            I => \N__6542\
        );

    \I__1302\ : InMux
    port map (
            O => \N__6546\,
            I => \N__6539\
        );

    \I__1301\ : InMux
    port map (
            O => \N__6545\,
            I => \N__6536\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__6542\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__6539\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__6536\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__1297\ : InMux
    port map (
            O => \N__6529\,
            I => \N__6525\
        );

    \I__1296\ : InMux
    port map (
            O => \N__6528\,
            I => \N__6522\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__6525\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__6522\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\
        );

    \I__1293\ : CascadeMux
    port map (
            O => \N__6517\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER46_cascade_\
        );

    \I__1292\ : CascadeMux
    port map (
            O => \N__6514\,
            I => \N__6511\
        );

    \I__1291\ : InMux
    port map (
            O => \N__6511\,
            I => \N__6507\
        );

    \I__1290\ : InMux
    port map (
            O => \N__6510\,
            I => \N__6504\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__6507\,
            I => \N__6501\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__6504\,
            I => \U712_CHIP_RAM.N_420\
        );

    \I__1287\ : Odrv4
    port map (
            O => \N__6501\,
            I => \U712_CHIP_RAM.N_420\
        );

    \I__1286\ : InMux
    port map (
            O => \N__6496\,
            I => \N__6488\
        );

    \I__1285\ : InMux
    port map (
            O => \N__6495\,
            I => \N__6479\
        );

    \I__1284\ : InMux
    port map (
            O => \N__6494\,
            I => \N__6479\
        );

    \I__1283\ : InMux
    port map (
            O => \N__6493\,
            I => \N__6479\
        );

    \I__1282\ : InMux
    port map (
            O => \N__6492\,
            I => \N__6475\
        );

    \I__1281\ : InMux
    port map (
            O => \N__6491\,
            I => \N__6472\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__6488\,
            I => \N__6469\
        );

    \I__1279\ : InMux
    port map (
            O => \N__6487\,
            I => \N__6464\
        );

    \I__1278\ : InMux
    port map (
            O => \N__6486\,
            I => \N__6464\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__6479\,
            I => \N__6461\
        );

    \I__1276\ : InMux
    port map (
            O => \N__6478\,
            I => \N__6458\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__6475\,
            I => \U712_CHIP_RAM.N_282\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__6472\,
            I => \U712_CHIP_RAM.N_282\
        );

    \I__1273\ : Odrv12
    port map (
            O => \N__6469\,
            I => \U712_CHIP_RAM.N_282\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__6464\,
            I => \U712_CHIP_RAM.N_282\
        );

    \I__1271\ : Odrv4
    port map (
            O => \N__6461\,
            I => \U712_CHIP_RAM.N_282\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__6458\,
            I => \U712_CHIP_RAM.N_282\
        );

    \I__1269\ : CascadeMux
    port map (
            O => \N__6445\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_a5_i_0_cascade_\
        );

    \I__1268\ : InMux
    port map (
            O => \N__6442\,
            I => \N__6439\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__6439\,
            I => \U712_CHIP_RAM.N_49\
        );

    \I__1266\ : IoInMux
    port map (
            O => \N__6436\,
            I => \N__6433\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__6433\,
            I => \N__6430\
        );

    \I__1264\ : IoSpan4Mux
    port map (
            O => \N__6430\,
            I => \N__6427\
        );

    \I__1263\ : IoSpan4Mux
    port map (
            O => \N__6427\,
            I => \N__6423\
        );

    \I__1262\ : InMux
    port map (
            O => \N__6426\,
            I => \N__6420\
        );

    \I__1261\ : Sp12to4
    port map (
            O => \N__6423\,
            I => \N__6417\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__6420\,
            I => \N__6414\
        );

    \I__1259\ : Span12Mux_s9_v
    port map (
            O => \N__6417\,
            I => \N__6410\
        );

    \I__1258\ : Span4Mux_v
    port map (
            O => \N__6414\,
            I => \N__6407\
        );

    \I__1257\ : InMux
    port map (
            O => \N__6413\,
            I => \N__6404\
        );

    \I__1256\ : Odrv12
    port map (
            O => \N__6410\,
            I => \DBDIR_c\
        );

    \I__1255\ : Odrv4
    port map (
            O => \N__6407\,
            I => \DBDIR_c\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__6404\,
            I => \DBDIR_c\
        );

    \I__1253\ : IoInMux
    port map (
            O => \N__6397\,
            I => \N__6394\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__6394\,
            I => \N__6391\
        );

    \I__1251\ : Span12Mux_s8_h
    port map (
            O => \N__6391\,
            I => \N__6388\
        );

    \I__1250\ : Span12Mux_v
    port map (
            O => \N__6388\,
            I => \N__6385\
        );

    \I__1249\ : Odrv12
    port map (
            O => \N__6385\,
            I => \N_218\
        );

    \I__1248\ : IoInMux
    port map (
            O => \N__6382\,
            I => \N__6379\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__6379\,
            I => \N__6376\
        );

    \I__1246\ : Span4Mux_s0_v
    port map (
            O => \N__6376\,
            I => \N__6373\
        );

    \I__1245\ : Span4Mux_v
    port map (
            O => \N__6373\,
            I => \N__6370\
        );

    \I__1244\ : Span4Mux_v
    port map (
            O => \N__6370\,
            I => \N__6367\
        );

    \I__1243\ : Span4Mux_h
    port map (
            O => \N__6367\,
            I => \N__6364\
        );

    \I__1242\ : Odrv4
    port map (
            O => \N__6364\,
            I => \RASn_c\
        );

    \I__1241\ : InMux
    port map (
            O => \N__6361\,
            I => \N__6358\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__6358\,
            I => \N__6355\
        );

    \I__1239\ : Span4Mux_v
    port map (
            O => \N__6355\,
            I => \N__6352\
        );

    \I__1238\ : Span4Mux_v
    port map (
            O => \N__6352\,
            I => \N__6349\
        );

    \I__1237\ : Sp12to4
    port map (
            O => \N__6349\,
            I => \N__6346\
        );

    \I__1236\ : Span12Mux_h
    port map (
            O => \N__6346\,
            I => \N__6343\
        );

    \I__1235\ : Odrv12
    port map (
            O => \N__6343\,
            I => \A_c_18\
        );

    \I__1234\ : CascadeMux
    port map (
            O => \N__6340\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_7_cascade_\
        );

    \I__1233\ : InMux
    port map (
            O => \N__6337\,
            I => \N__6334\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__6334\,
            I => \N__6331\
        );

    \I__1231\ : Span4Mux_v
    port map (
            O => \N__6331\,
            I => \N__6328\
        );

    \I__1230\ : Span4Mux_v
    port map (
            O => \N__6328\,
            I => \N__6325\
        );

    \I__1229\ : Sp12to4
    port map (
            O => \N__6325\,
            I => \N__6322\
        );

    \I__1228\ : Span12Mux_h
    port map (
            O => \N__6322\,
            I => \N__6319\
        );

    \I__1227\ : Odrv12
    port map (
            O => \N__6319\,
            I => \A_c_16\
        );

    \I__1226\ : CascadeMux
    port map (
            O => \N__6316\,
            I => \U712_CHIP_RAM.N_296_cascade_\
        );

    \I__1225\ : InMux
    port map (
            O => \N__6313\,
            I => \N__6310\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__6310\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_i_0_a2_0_0_0\
        );

    \I__1223\ : InMux
    port map (
            O => \N__6307\,
            I => \N__6304\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__6304\,
            I => \N__6301\
        );

    \I__1221\ : Odrv12
    port map (
            O => \N__6301\,
            I => \U712_CHIP_RAM.N_403\
        );

    \I__1220\ : InMux
    port map (
            O => \N__6298\,
            I => \N__6289\
        );

    \I__1219\ : InMux
    port map (
            O => \N__6297\,
            I => \N__6289\
        );

    \I__1218\ : InMux
    port map (
            O => \N__6296\,
            I => \N__6289\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__6289\,
            I => \U712_CHIP_RAM.N_309\
        );

    \I__1216\ : CascadeMux
    port map (
            O => \N__6286\,
            I => \N__6281\
        );

    \I__1215\ : InMux
    port map (
            O => \N__6285\,
            I => \N__6278\
        );

    \I__1214\ : InMux
    port map (
            O => \N__6284\,
            I => \N__6273\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6281\,
            I => \N__6273\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__6278\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__6273\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\
        );

    \I__1210\ : InMux
    port map (
            O => \N__6268\,
            I => \N__6265\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__6265\,
            I => \N__6262\
        );

    \I__1208\ : Span4Mux_v
    port map (
            O => \N__6262\,
            I => \N__6259\
        );

    \I__1207\ : Odrv4
    port map (
            O => \N__6259\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1206\ : CascadeMux
    port map (
            O => \N__6256\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_1_cascade_\
        );

    \I__1205\ : InMux
    port map (
            O => \N__6253\,
            I => \N__6250\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__6250\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0\
        );

    \I__1203\ : InMux
    port map (
            O => \N__6247\,
            I => \N__6242\
        );

    \I__1202\ : InMux
    port map (
            O => \N__6246\,
            I => \N__6237\
        );

    \I__1201\ : InMux
    port map (
            O => \N__6245\,
            I => \N__6237\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__6242\,
            I => \U712_CHIP_RAM.N_285\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__6237\,
            I => \U712_CHIP_RAM.N_285\
        );

    \I__1198\ : CascadeMux
    port map (
            O => \N__6232\,
            I => \N__6228\
        );

    \I__1197\ : InMux
    port map (
            O => \N__6231\,
            I => \N__6225\
        );

    \I__1196\ : InMux
    port map (
            O => \N__6228\,
            I => \N__6222\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__6225\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__6222\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\
        );

    \I__1193\ : InMux
    port map (
            O => \N__6217\,
            I => \N__6214\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__6214\,
            I => \N__6211\
        );

    \I__1191\ : Span4Mux_h
    port map (
            O => \N__6211\,
            I => \N__6208\
        );

    \I__1190\ : Odrv4
    port map (
            O => \N__6208\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__1189\ : CascadeMux
    port map (
            O => \N__6205\,
            I => \U712_CHIP_RAM.DMA_CYCLE_7_cascade_\
        );

    \I__1188\ : InMux
    port map (
            O => \N__6202\,
            I => \N__6198\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6201\,
            I => \N__6195\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__6198\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__6195\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0\
        );

    \I__1184\ : IoInMux
    port map (
            O => \N__6190\,
            I => \N__6187\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__6187\,
            I => \N__6184\
        );

    \I__1182\ : IoSpan4Mux
    port map (
            O => \N__6184\,
            I => \N__6181\
        );

    \I__1181\ : Span4Mux_s3_v
    port map (
            O => \N__6181\,
            I => \N__6174\
        );

    \I__1180\ : InMux
    port map (
            O => \N__6180\,
            I => \N__6171\
        );

    \I__1179\ : InMux
    port map (
            O => \N__6179\,
            I => \N__6168\
        );

    \I__1178\ : InMux
    port map (
            O => \N__6178\,
            I => \N__6163\
        );

    \I__1177\ : InMux
    port map (
            O => \N__6177\,
            I => \N__6163\
        );

    \I__1176\ : Sp12to4
    port map (
            O => \N__6174\,
            I => \N__6160\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6171\,
            I => \N__6155\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__6168\,
            I => \N__6155\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__6163\,
            I => \N__6152\
        );

    \I__1172\ : Span12Mux_v
    port map (
            O => \N__6160\,
            I => \N__6148\
        );

    \I__1171\ : Span4Mux_v
    port map (
            O => \N__6155\,
            I => \N__6145\
        );

    \I__1170\ : Span4Mux_v
    port map (
            O => \N__6152\,
            I => \N__6142\
        );

    \I__1169\ : InMux
    port map (
            O => \N__6151\,
            I => \N__6139\
        );

    \I__1168\ : Odrv12
    port map (
            O => \N__6148\,
            I => \DBENn_c\
        );

    \I__1167\ : Odrv4
    port map (
            O => \N__6145\,
            I => \DBENn_c\
        );

    \I__1166\ : Odrv4
    port map (
            O => \N__6142\,
            I => \DBENn_c\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__6139\,
            I => \DBENn_c\
        );

    \I__1164\ : InMux
    port map (
            O => \N__6130\,
            I => \N__6127\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__6127\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_0_a2_0_0\
        );

    \I__1162\ : InMux
    port map (
            O => \N__6124\,
            I => \N__6121\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__6121\,
            I => \N__6118\
        );

    \I__1160\ : Odrv4
    port map (
            O => \N__6118\,
            I => \U712_CHIP_RAM.N_427\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6115\,
            I => \N__6112\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__6112\,
            I => \U712_CHIP_RAM.N_421\
        );

    \I__1157\ : InMux
    port map (
            O => \N__6109\,
            I => \N__6106\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__6106\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__6103\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_cascade_\
        );

    \I__1154\ : InMux
    port map (
            O => \N__6100\,
            I => \N__6096\
        );

    \I__1153\ : CascadeMux
    port map (
            O => \N__6099\,
            I => \N__6093\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__6096\,
            I => \N__6090\
        );

    \I__1151\ : InMux
    port map (
            O => \N__6093\,
            I => \N__6087\
        );

    \I__1150\ : Odrv4
    port map (
            O => \N__6090\,
            I => \U712_CHIP_RAM.N_296\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__6087\,
            I => \U712_CHIP_RAM.N_296\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6082\,
            I => \N__6079\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__6079\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_4\
        );

    \I__1146\ : CascadeMux
    port map (
            O => \N__6076\,
            I => \N__6073\
        );

    \I__1145\ : InMux
    port map (
            O => \N__6073\,
            I => \N__6070\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__6070\,
            I => \N__6067\
        );

    \I__1143\ : Span4Mux_v
    port map (
            O => \N__6067\,
            I => \N__6064\
        );

    \I__1142\ : Sp12to4
    port map (
            O => \N__6064\,
            I => \N__6061\
        );

    \I__1141\ : Span12Mux_h
    port map (
            O => \N__6061\,
            I => \N__6058\
        );

    \I__1140\ : Odrv12
    port map (
            O => \N__6058\,
            I => \A_c_13\
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__6055\,
            I => \U712_CHIP_RAM.N_493_cascade_\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__6052\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_cascade_\
        );

    \I__1137\ : InMux
    port map (
            O => \N__6049\,
            I => \N__6046\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__6046\,
            I => \U712_CHIP_RAM.N_317\
        );

    \I__1135\ : IoInMux
    port map (
            O => \N__6043\,
            I => \N__6040\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__6040\,
            I => \N__6037\
        );

    \I__1133\ : Span12Mux_s2_h
    port map (
            O => \N__6037\,
            I => \N__6034\
        );

    \I__1132\ : Span12Mux_h
    port map (
            O => \N__6034\,
            I => \N__6031\
        );

    \I__1131\ : Odrv12
    port map (
            O => \N__6031\,
            I => \CMA_c_6\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6028\,
            I => \N__6025\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6025\,
            I => \N__6022\
        );

    \I__1128\ : Span4Mux_v
    port map (
            O => \N__6022\,
            I => \N__6019\
        );

    \I__1127\ : Sp12to4
    port map (
            O => \N__6019\,
            I => \N__6016\
        );

    \I__1126\ : Span12Mux_h
    port map (
            O => \N__6016\,
            I => \N__6013\
        );

    \I__1125\ : Span12Mux_v
    port map (
            O => \N__6013\,
            I => \N__6010\
        );

    \I__1124\ : Odrv12
    port map (
            O => \N__6010\,
            I => \A_c_19\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__6007\,
            I => \U712_CHIP_RAM.CMA_5_i_0_8_cascade_\
        );

    \I__1122\ : IoInMux
    port map (
            O => \N__6004\,
            I => \N__6001\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__6001\,
            I => \N__5998\
        );

    \I__1120\ : IoSpan4Mux
    port map (
            O => \N__5998\,
            I => \N__5995\
        );

    \I__1119\ : Span4Mux_s3_h
    port map (
            O => \N__5995\,
            I => \N__5992\
        );

    \I__1118\ : Sp12to4
    port map (
            O => \N__5992\,
            I => \N__5989\
        );

    \I__1117\ : Span12Mux_h
    port map (
            O => \N__5989\,
            I => \N__5986\
        );

    \I__1116\ : Odrv12
    port map (
            O => \N__5986\,
            I => \CMA_c_9\
        );

    \I__1115\ : SRMux
    port map (
            O => \N__5983\,
            I => \N__5980\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__5980\,
            I => \N__5976\
        );

    \I__1113\ : InMux
    port map (
            O => \N__5979\,
            I => \N__5973\
        );

    \I__1112\ : Span4Mux_v
    port map (
            O => \N__5976\,
            I => \N__5970\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__5973\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__1110\ : Odrv4
    port map (
            O => \N__5970\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__1109\ : CascadeMux
    port map (
            O => \N__5965\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_cascade_\
        );

    \I__1108\ : InMux
    port map (
            O => \N__5962\,
            I => \N__5959\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__5959\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0\
        );

    \I__1106\ : InMux
    port map (
            O => \N__5956\,
            I => \N__5952\
        );

    \I__1105\ : InMux
    port map (
            O => \N__5955\,
            I => \N__5949\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__5952\,
            I => \CPU_TACKm\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__5949\,
            I => \CPU_TACKm\
        );

    \I__1102\ : InMux
    port map (
            O => \N__5944\,
            I => \N__5941\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__5941\,
            I => \N__5936\
        );

    \I__1100\ : InMux
    port map (
            O => \N__5940\,
            I => \N__5933\
        );

    \I__1099\ : InMux
    port map (
            O => \N__5939\,
            I => \N__5930\
        );

    \I__1098\ : Odrv12
    port map (
            O => \N__5936\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__5933\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__5930\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__1095\ : InMux
    port map (
            O => \N__5923\,
            I => \N__5920\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__5920\,
            I => \N__5916\
        );

    \I__1093\ : InMux
    port map (
            O => \N__5919\,
            I => \N__5913\
        );

    \I__1092\ : Odrv12
    port map (
            O => \N__5916\,
            I => \U712_REG_SM.LDS_OUTZ0\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__5913\,
            I => \U712_REG_SM.LDS_OUTZ0\
        );

    \I__1090\ : IoInMux
    port map (
            O => \N__5908\,
            I => \N__5905\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__5905\,
            I => \N__5902\
        );

    \I__1088\ : IoSpan4Mux
    port map (
            O => \N__5902\,
            I => \N__5899\
        );

    \I__1087\ : Span4Mux_s2_v
    port map (
            O => \N__5899\,
            I => \N__5896\
        );

    \I__1086\ : Sp12to4
    port map (
            O => \N__5896\,
            I => \N__5893\
        );

    \I__1085\ : Span12Mux_v
    port map (
            O => \N__5893\,
            I => \N__5890\
        );

    \I__1084\ : Odrv12
    port map (
            O => \N__5890\,
            I => \U712_REG_SM_un1_LDSn_i\
        );

    \I__1083\ : InMux
    port map (
            O => \N__5887\,
            I => \N__5884\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__5884\,
            I => \U712_CHIP_RAM.N_311\
        );

    \I__1081\ : IoInMux
    port map (
            O => \N__5881\,
            I => \N__5878\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__5878\,
            I => \N__5875\
        );

    \I__1079\ : Span4Mux_s1_v
    port map (
            O => \N__5875\,
            I => \N__5872\
        );

    \I__1078\ : Span4Mux_v
    port map (
            O => \N__5872\,
            I => \N__5869\
        );

    \I__1077\ : Span4Mux_v
    port map (
            O => \N__5869\,
            I => \N__5866\
        );

    \I__1076\ : Odrv4
    port map (
            O => \N__5866\,
            I => \CMA_c_0\
        );

    \I__1075\ : InMux
    port map (
            O => \N__5863\,
            I => \N__5860\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__5860\,
            I => \U712_CHIP_RAM.N_312\
        );

    \I__1073\ : IoInMux
    port map (
            O => \N__5857\,
            I => \N__5854\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__5854\,
            I => \N__5851\
        );

    \I__1071\ : Span4Mux_s2_v
    port map (
            O => \N__5851\,
            I => \N__5848\
        );

    \I__1070\ : Span4Mux_v
    port map (
            O => \N__5848\,
            I => \N__5845\
        );

    \I__1069\ : Span4Mux_v
    port map (
            O => \N__5845\,
            I => \N__5842\
        );

    \I__1068\ : Odrv4
    port map (
            O => \N__5842\,
            I => \CMA_c_1\
        );

    \I__1067\ : InMux
    port map (
            O => \N__5839\,
            I => \N__5836\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__5836\,
            I => \U712_CHIP_RAM.N_316\
        );

    \I__1065\ : IoInMux
    port map (
            O => \N__5833\,
            I => \N__5830\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__5830\,
            I => \N__5827\
        );

    \I__1063\ : Span4Mux_s2_h
    port map (
            O => \N__5827\,
            I => \N__5824\
        );

    \I__1062\ : Span4Mux_v
    port map (
            O => \N__5824\,
            I => \N__5821\
        );

    \I__1061\ : Sp12to4
    port map (
            O => \N__5821\,
            I => \N__5818\
        );

    \I__1060\ : Span12Mux_h
    port map (
            O => \N__5818\,
            I => \N__5815\
        );

    \I__1059\ : Odrv12
    port map (
            O => \N__5815\,
            I => \CMA_c_5\
        );

    \I__1058\ : CascadeMux
    port map (
            O => \N__5812\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_cascade_\
        );

    \I__1057\ : InMux
    port map (
            O => \N__5809\,
            I => \N__5806\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__5806\,
            I => \N__5803\
        );

    \I__1055\ : Span12Mux_v
    port map (
            O => \N__5803\,
            I => \N__5800\
        );

    \I__1054\ : Span12Mux_h
    port map (
            O => \N__5800\,
            I => \N__5797\
        );

    \I__1053\ : Odrv12
    port map (
            O => \N__5797\,
            I => \A_c_6\
        );

    \I__1052\ : InMux
    port map (
            O => \N__5794\,
            I => \N__5790\
        );

    \I__1051\ : InMux
    port map (
            O => \N__5793\,
            I => \N__5787\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__5790\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__5787\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1048\ : CascadeMux
    port map (
            O => \N__5782\,
            I => \N__5779\
        );

    \I__1047\ : InMux
    port map (
            O => \N__5779\,
            I => \N__5776\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__5776\,
            I => \N__5772\
        );

    \I__1045\ : InMux
    port map (
            O => \N__5775\,
            I => \N__5768\
        );

    \I__1044\ : Span4Mux_v
    port map (
            O => \N__5772\,
            I => \N__5765\
        );

    \I__1043\ : InMux
    port map (
            O => \N__5771\,
            I => \N__5762\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__5768\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__1041\ : Odrv4
    port map (
            O => \N__5765\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__5762\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__1039\ : InMux
    port map (
            O => \N__5755\,
            I => \N__5752\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__5752\,
            I => \N__5749\
        );

    \I__1037\ : Span4Mux_h
    port map (
            O => \N__5749\,
            I => \N__5745\
        );

    \I__1036\ : InMux
    port map (
            O => \N__5748\,
            I => \N__5742\
        );

    \I__1035\ : Odrv4
    port map (
            O => \N__5745\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__5742\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__1033\ : InMux
    port map (
            O => \N__5737\,
            I => \N__5734\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__5734\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_3_1\
        );

    \I__1031\ : CascadeMux
    port map (
            O => \N__5731\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_2_1_cascade_\
        );

    \I__1030\ : CascadeMux
    port map (
            O => \N__5728\,
            I => \U712_CHIP_RAM.N_421_cascade_\
        );

    \I__1029\ : CascadeMux
    port map (
            O => \N__5725\,
            I => \U712_CHIP_RAM.N_293_cascade_\
        );

    \I__1028\ : CascadeMux
    port map (
            O => \N__5722\,
            I => \U712_CHIP_RAM.N_309_cascade_\
        );

    \I__1027\ : InMux
    port map (
            O => \N__5719\,
            I => \N__5716\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__5716\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0_a2_0_a2_0\
        );

    \I__1025\ : InMux
    port map (
            O => \N__5713\,
            I => \N__5710\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__5710\,
            I => \N__5707\
        );

    \I__1023\ : Span4Mux_v
    port map (
            O => \N__5707\,
            I => \N__5704\
        );

    \I__1022\ : Sp12to4
    port map (
            O => \N__5704\,
            I => \N__5701\
        );

    \I__1021\ : Span12Mux_v
    port map (
            O => \N__5701\,
            I => \N__5698\
        );

    \I__1020\ : Span12Mux_h
    port map (
            O => \N__5698\,
            I => \N__5695\
        );

    \I__1019\ : Odrv12
    port map (
            O => \N__5695\,
            I => \DBRn_c\
        );

    \I__1018\ : CascadeMux
    port map (
            O => \N__5692\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_0_cascade_\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__5689\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_2_cascade_\
        );

    \I__1016\ : InMux
    port map (
            O => \N__5686\,
            I => \N__5680\
        );

    \I__1015\ : InMux
    port map (
            O => \N__5685\,
            I => \N__5680\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__5680\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1013\ : InMux
    port map (
            O => \N__5677\,
            I => \N__5672\
        );

    \I__1012\ : InMux
    port map (
            O => \N__5676\,
            I => \N__5667\
        );

    \I__1011\ : InMux
    port map (
            O => \N__5675\,
            I => \N__5667\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__5672\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__5667\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1008\ : CascadeMux
    port map (
            O => \N__5662\,
            I => \U712_CHIP_RAM.N_314_cascade_\
        );

    \I__1007\ : IoInMux
    port map (
            O => \N__5659\,
            I => \N__5656\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__5656\,
            I => \N__5653\
        );

    \I__1005\ : IoSpan4Mux
    port map (
            O => \N__5653\,
            I => \N__5650\
        );

    \I__1004\ : Span4Mux_s1_h
    port map (
            O => \N__5650\,
            I => \N__5647\
        );

    \I__1003\ : Sp12to4
    port map (
            O => \N__5647\,
            I => \N__5644\
        );

    \I__1002\ : Span12Mux_h
    port map (
            O => \N__5644\,
            I => \N__5641\
        );

    \I__1001\ : Odrv12
    port map (
            O => \N__5641\,
            I => \CMA_c_3\
        );

    \I__1000\ : InMux
    port map (
            O => \N__5638\,
            I => \N__5635\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__5635\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__998\ : InMux
    port map (
            O => \N__5632\,
            I => \N__5629\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__5629\,
            I => \N__5626\
        );

    \I__996\ : Odrv4
    port map (
            O => \N__5626\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_5\
        );

    \I__995\ : InMux
    port map (
            O => \N__5623\,
            I => \N__5619\
        );

    \I__994\ : InMux
    port map (
            O => \N__5622\,
            I => \N__5616\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__5619\,
            I => \N__5611\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__5616\,
            I => \N__5611\
        );

    \I__991\ : Span4Mux_v
    port map (
            O => \N__5611\,
            I => \N__5608\
        );

    \I__990\ : Span4Mux_v
    port map (
            O => \N__5608\,
            I => \N__5605\
        );

    \I__989\ : Sp12to4
    port map (
            O => \N__5605\,
            I => \N__5602\
        );

    \I__988\ : Span12Mux_h
    port map (
            O => \N__5602\,
            I => \N__5599\
        );

    \I__987\ : Odrv12
    port map (
            O => \N__5599\,
            I => \DRA_c_6\
        );

    \I__986\ : InMux
    port map (
            O => \N__5596\,
            I => \N__5593\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__5593\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__984\ : InMux
    port map (
            O => \N__5590\,
            I => \N__5587\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__5587\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__982\ : InMux
    port map (
            O => \N__5584\,
            I => \N__5581\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__5581\,
            I => \N__5577\
        );

    \I__980\ : InMux
    port map (
            O => \N__5580\,
            I => \N__5574\
        );

    \I__979\ : Span4Mux_v
    port map (
            O => \N__5577\,
            I => \N__5571\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__5574\,
            I => \N__5568\
        );

    \I__977\ : Span4Mux_v
    port map (
            O => \N__5571\,
            I => \N__5565\
        );

    \I__976\ : Sp12to4
    port map (
            O => \N__5568\,
            I => \N__5562\
        );

    \I__975\ : Sp12to4
    port map (
            O => \N__5565\,
            I => \N__5557\
        );

    \I__974\ : Span12Mux_v
    port map (
            O => \N__5562\,
            I => \N__5557\
        );

    \I__973\ : Span12Mux_h
    port map (
            O => \N__5557\,
            I => \N__5554\
        );

    \I__972\ : Odrv12
    port map (
            O => \N__5554\,
            I => \DRA_c_5\
        );

    \I__971\ : InMux
    port map (
            O => \N__5551\,
            I => \N__5548\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__5548\,
            I => \N__5545\
        );

    \I__969\ : Odrv4
    port map (
            O => \N__5545\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__968\ : InMux
    port map (
            O => \N__5542\,
            I => \N__5539\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__5539\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__966\ : InMux
    port map (
            O => \N__5536\,
            I => \N__5533\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__5533\,
            I => \N__5530\
        );

    \I__964\ : Sp12to4
    port map (
            O => \N__5530\,
            I => \N__5527\
        );

    \I__963\ : Span12Mux_v
    port map (
            O => \N__5527\,
            I => \N__5524\
        );

    \I__962\ : Span12Mux_h
    port map (
            O => \N__5524\,
            I => \N__5521\
        );

    \I__961\ : Odrv12
    port map (
            O => \N__5521\,
            I => \A_c_8\
        );

    \I__960\ : CascadeMux
    port map (
            O => \N__5518\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_6_cascade_\
        );

    \I__959\ : InMux
    port map (
            O => \N__5515\,
            I => \N__5512\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__5512\,
            I => \N__5509\
        );

    \I__957\ : Span4Mux_v
    port map (
            O => \N__5509\,
            I => \N__5506\
        );

    \I__956\ : Span4Mux_v
    port map (
            O => \N__5506\,
            I => \N__5503\
        );

    \I__955\ : Sp12to4
    port map (
            O => \N__5503\,
            I => \N__5500\
        );

    \I__954\ : Span12Mux_h
    port map (
            O => \N__5500\,
            I => \N__5497\
        );

    \I__953\ : Odrv12
    port map (
            O => \N__5497\,
            I => \A_c_15\
        );

    \I__952\ : InMux
    port map (
            O => \N__5494\,
            I => \N__5491\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__5491\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__950\ : InMux
    port map (
            O => \N__5488\,
            I => \N__5485\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__5485\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__948\ : InMux
    port map (
            O => \N__5482\,
            I => \N__5479\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__5479\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__946\ : InMux
    port map (
            O => \N__5476\,
            I => \N__5473\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__5473\,
            I => \N__5470\
        );

    \I__944\ : Span4Mux_v
    port map (
            O => \N__5470\,
            I => \N__5467\
        );

    \I__943\ : Span4Mux_v
    port map (
            O => \N__5467\,
            I => \N__5464\
        );

    \I__942\ : Sp12to4
    port map (
            O => \N__5464\,
            I => \N__5461\
        );

    \I__941\ : Span12Mux_h
    port map (
            O => \N__5461\,
            I => \N__5458\
        );

    \I__940\ : Odrv12
    port map (
            O => \N__5458\,
            I => \A_c_9\
        );

    \I__939\ : InMux
    port map (
            O => \N__5455\,
            I => \N__5452\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__5452\,
            I => \N__5449\
        );

    \I__937\ : Span4Mux_h
    port map (
            O => \N__5449\,
            I => \N__5446\
        );

    \I__936\ : Span4Mux_v
    port map (
            O => \N__5446\,
            I => \N__5443\
        );

    \I__935\ : Sp12to4
    port map (
            O => \N__5443\,
            I => \N__5440\
        );

    \I__934\ : Span12Mux_h
    port map (
            O => \N__5440\,
            I => \N__5437\
        );

    \I__933\ : Span12Mux_v
    port map (
            O => \N__5437\,
            I => \N__5434\
        );

    \I__932\ : Odrv12
    port map (
            O => \N__5434\,
            I => \A_c_2\
        );

    \I__931\ : CascadeMux
    port map (
            O => \N__5431\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_0_cascade_\
        );

    \I__930\ : InMux
    port map (
            O => \N__5428\,
            I => \N__5425\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__5425\,
            I => \N__5422\
        );

    \I__928\ : Odrv4
    port map (
            O => \N__5422\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__927\ : InMux
    port map (
            O => \N__5419\,
            I => \N__5416\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__5416\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__925\ : InMux
    port map (
            O => \N__5413\,
            I => \N__5410\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__5410\,
            I => \N__5407\
        );

    \I__923\ : Span4Mux_v
    port map (
            O => \N__5407\,
            I => \N__5404\
        );

    \I__922\ : Sp12to4
    port map (
            O => \N__5404\,
            I => \N__5401\
        );

    \I__921\ : Span12Mux_h
    port map (
            O => \N__5401\,
            I => \N__5398\
        );

    \I__920\ : Odrv12
    port map (
            O => \N__5398\,
            I => \A_c_10\
        );

    \I__919\ : InMux
    port map (
            O => \N__5395\,
            I => \N__5392\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__5392\,
            I => \N__5389\
        );

    \I__917\ : Span4Mux_v
    port map (
            O => \N__5389\,
            I => \N__5386\
        );

    \I__916\ : Sp12to4
    port map (
            O => \N__5386\,
            I => \N__5383\
        );

    \I__915\ : Span12Mux_h
    port map (
            O => \N__5383\,
            I => \N__5380\
        );

    \I__914\ : Span12Mux_v
    port map (
            O => \N__5380\,
            I => \N__5377\
        );

    \I__913\ : Odrv12
    port map (
            O => \N__5377\,
            I => \A_c_3\
        );

    \I__912\ : CascadeMux
    port map (
            O => \N__5374\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_1_cascade_\
        );

    \I__911\ : IoInMux
    port map (
            O => \N__5371\,
            I => \N__5368\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__5368\,
            I => \N__5365\
        );

    \I__909\ : Span4Mux_s2_v
    port map (
            O => \N__5365\,
            I => \N__5362\
        );

    \I__908\ : Span4Mux_v
    port map (
            O => \N__5362\,
            I => \N__5359\
        );

    \I__907\ : Span4Mux_v
    port map (
            O => \N__5359\,
            I => \N__5356\
        );

    \I__906\ : Span4Mux_h
    port map (
            O => \N__5356\,
            I => \N__5353\
        );

    \I__905\ : Odrv4
    port map (
            O => \N__5353\,
            I => \CMA_c_10\
        );

    \I__904\ : InMux
    port map (
            O => \N__5350\,
            I => \N__5347\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5347\,
            I => \N__5344\
        );

    \I__902\ : Odrv4
    port map (
            O => \N__5344\,
            I => \U712_CHIP_RAM.N_313\
        );

    \I__901\ : IoInMux
    port map (
            O => \N__5341\,
            I => \N__5338\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__5338\,
            I => \N__5335\
        );

    \I__899\ : IoSpan4Mux
    port map (
            O => \N__5335\,
            I => \N__5332\
        );

    \I__898\ : Span4Mux_s3_v
    port map (
            O => \N__5332\,
            I => \N__5329\
        );

    \I__897\ : Span4Mux_v
    port map (
            O => \N__5329\,
            I => \N__5326\
        );

    \I__896\ : Odrv4
    port map (
            O => \N__5326\,
            I => \CMA_c_2\
        );

    \I__895\ : InMux
    port map (
            O => \N__5323\,
            I => \N__5320\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__5320\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__893\ : InMux
    port map (
            O => \N__5317\,
            I => \N__5314\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__5314\,
            I => \N__5311\
        );

    \I__891\ : Span4Mux_v
    port map (
            O => \N__5311\,
            I => \N__5308\
        );

    \I__890\ : Sp12to4
    port map (
            O => \N__5308\,
            I => \N__5305\
        );

    \I__889\ : Span12Mux_h
    port map (
            O => \N__5305\,
            I => \N__5302\
        );

    \I__888\ : Span12Mux_v
    port map (
            O => \N__5302\,
            I => \N__5299\
        );

    \I__887\ : Odrv12
    port map (
            O => \N__5299\,
            I => \A_c_5\
        );

    \I__886\ : CascadeMux
    port map (
            O => \N__5296\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_3_cascade_\
        );

    \I__885\ : InMux
    port map (
            O => \N__5293\,
            I => \N__5290\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__5290\,
            I => \N__5287\
        );

    \I__883\ : Span4Mux_v
    port map (
            O => \N__5287\,
            I => \N__5284\
        );

    \I__882\ : Sp12to4
    port map (
            O => \N__5284\,
            I => \N__5281\
        );

    \I__881\ : Span12Mux_h
    port map (
            O => \N__5281\,
            I => \N__5278\
        );

    \I__880\ : Odrv12
    port map (
            O => \N__5278\,
            I => \A_c_12\
        );

    \I__879\ : CascadeMux
    port map (
            O => \N__5275\,
            I => \N__5272\
        );

    \I__878\ : InMux
    port map (
            O => \N__5272\,
            I => \N__5269\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__5269\,
            I => \N__5266\
        );

    \I__876\ : Span4Mux_v
    port map (
            O => \N__5266\,
            I => \N__5263\
        );

    \I__875\ : Odrv4
    port map (
            O => \N__5263\,
            I => \U712_BYTE_ENABLE.N_392\
        );

    \I__874\ : InMux
    port map (
            O => \N__5260\,
            I => \N__5257\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__5257\,
            I => \N__5254\
        );

    \I__872\ : Span4Mux_v
    port map (
            O => \N__5254\,
            I => \N__5251\
        );

    \I__871\ : Odrv4
    port map (
            O => \N__5251\,
            I => \U712_BYTE_ENABLE.N_388\
        );

    \I__870\ : InMux
    port map (
            O => \N__5248\,
            I => \N__5243\
        );

    \I__869\ : InMux
    port map (
            O => \N__5247\,
            I => \N__5240\
        );

    \I__868\ : InMux
    port map (
            O => \N__5246\,
            I => \N__5237\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__5243\,
            I => \N__5234\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__5240\,
            I => \N__5229\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__5237\,
            I => \N__5229\
        );

    \I__864\ : Span4Mux_v
    port map (
            O => \N__5234\,
            I => \N__5226\
        );

    \I__863\ : Span12Mux_v
    port map (
            O => \N__5229\,
            I => \N__5223\
        );

    \I__862\ : Sp12to4
    port map (
            O => \N__5226\,
            I => \N__5220\
        );

    \I__861\ : Span12Mux_h
    port map (
            O => \N__5223\,
            I => \N__5217\
        );

    \I__860\ : Span12Mux_h
    port map (
            O => \N__5220\,
            I => \N__5214\
        );

    \I__859\ : Span12Mux_v
    port map (
            O => \N__5217\,
            I => \N__5211\
        );

    \I__858\ : Span12Mux_v
    port map (
            O => \N__5214\,
            I => \N__5208\
        );

    \I__857\ : Odrv12
    port map (
            O => \N__5211\,
            I => \CASLn_c\
        );

    \I__856\ : Odrv12
    port map (
            O => \N__5208\,
            I => \CASLn_c\
        );

    \I__855\ : CascadeMux
    port map (
            O => \N__5203\,
            I => \N__5199\
        );

    \I__854\ : InMux
    port map (
            O => \N__5202\,
            I => \N__5191\
        );

    \I__853\ : InMux
    port map (
            O => \N__5199\,
            I => \N__5191\
        );

    \I__852\ : InMux
    port map (
            O => \N__5198\,
            I => \N__5191\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__5191\,
            I => \N__5188\
        );

    \I__850\ : Span12Mux_v
    port map (
            O => \N__5188\,
            I => \N__5185\
        );

    \I__849\ : Span12Mux_h
    port map (
            O => \N__5185\,
            I => \N__5182\
        );

    \I__848\ : Span12Mux_v
    port map (
            O => \N__5182\,
            I => \N__5179\
        );

    \I__847\ : Odrv12
    port map (
            O => \N__5179\,
            I => \CASUn_c\
        );

    \I__846\ : InMux
    port map (
            O => \N__5176\,
            I => \N__5173\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__5173\,
            I => \N__5170\
        );

    \I__844\ : Span4Mux_v
    port map (
            O => \N__5170\,
            I => \N__5167\
        );

    \I__843\ : Sp12to4
    port map (
            O => \N__5167\,
            I => \N__5163\
        );

    \I__842\ : IoInMux
    port map (
            O => \N__5166\,
            I => \N__5160\
        );

    \I__841\ : Span12Mux_h
    port map (
            O => \N__5163\,
            I => \N__5157\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__5160\,
            I => \N__5154\
        );

    \I__839\ : Span12Mux_v
    port map (
            O => \N__5157\,
            I => \N__5151\
        );

    \I__838\ : IoSpan4Mux
    port map (
            O => \N__5154\,
            I => \N__5148\
        );

    \I__837\ : Odrv12
    port map (
            O => \N__5151\,
            I => \RAMENn_c\
        );

    \I__836\ : Odrv4
    port map (
            O => \N__5148\,
            I => \RAMENn_c\
        );

    \I__835\ : CascadeMux
    port map (
            O => \N__5143\,
            I => \N__5140\
        );

    \I__834\ : InMux
    port map (
            O => \N__5140\,
            I => \N__5136\
        );

    \I__833\ : InMux
    port map (
            O => \N__5139\,
            I => \N__5133\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__5136\,
            I => \N__5130\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__5133\,
            I => \N__5127\
        );

    \I__830\ : Span4Mux_v
    port map (
            O => \N__5130\,
            I => \N__5124\
        );

    \I__829\ : Span4Mux_v
    port map (
            O => \N__5127\,
            I => \N__5121\
        );

    \I__828\ : Sp12to4
    port map (
            O => \N__5124\,
            I => \N__5116\
        );

    \I__827\ : Sp12to4
    port map (
            O => \N__5121\,
            I => \N__5116\
        );

    \I__826\ : Span12Mux_h
    port map (
            O => \N__5116\,
            I => \N__5113\
        );

    \I__825\ : Span12Mux_v
    port map (
            O => \N__5113\,
            I => \N__5110\
        );

    \I__824\ : Odrv12
    port map (
            O => \N__5110\,
            I => \TSn_c\
        );

    \I__823\ : InMux
    port map (
            O => \N__5107\,
            I => \N__5103\
        );

    \I__822\ : InMux
    port map (
            O => \N__5106\,
            I => \N__5100\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__5103\,
            I => \REG_TACK\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__5100\,
            I => \REG_TACK\
        );

    \I__819\ : CascadeMux
    port map (
            O => \N__5095\,
            I => \N__5091\
        );

    \I__818\ : InMux
    port map (
            O => \N__5094\,
            I => \N__5088\
        );

    \I__817\ : InMux
    port map (
            O => \N__5091\,
            I => \N__5084\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__5088\,
            I => \N__5081\
        );

    \I__815\ : InMux
    port map (
            O => \N__5087\,
            I => \N__5078\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__5084\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__813\ : Odrv4
    port map (
            O => \N__5081\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5078\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__811\ : InMux
    port map (
            O => \N__5071\,
            I => \N__5065\
        );

    \I__810\ : InMux
    port map (
            O => \N__5070\,
            I => \N__5065\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__5065\,
            I => \N__5061\
        );

    \I__808\ : InMux
    port map (
            O => \N__5064\,
            I => \N__5057\
        );

    \I__807\ : Span4Mux_v
    port map (
            O => \N__5061\,
            I => \N__5054\
        );

    \I__806\ : InMux
    port map (
            O => \N__5060\,
            I => \N__5051\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__5057\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__804\ : Odrv4
    port map (
            O => \N__5054\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__5051\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__802\ : InMux
    port map (
            O => \N__5044\,
            I => \N__5041\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__5041\,
            I => \N__5038\
        );

    \I__800\ : Span4Mux_v
    port map (
            O => \N__5038\,
            I => \N__5035\
        );

    \I__799\ : Span4Mux_v
    port map (
            O => \N__5035\,
            I => \N__5032\
        );

    \I__798\ : Odrv4
    port map (
            O => \N__5032\,
            I => \TACK_EN_i_ess\
        );

    \I__797\ : CEMux
    port map (
            O => \N__5029\,
            I => \N__5026\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__5026\,
            I => \U712_CYCLE_TERM.N_305_i_0_en_0\
        );

    \I__795\ : IoInMux
    port map (
            O => \N__5023\,
            I => \N__5020\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__5020\,
            I => \N__5017\
        );

    \I__793\ : Odrv12
    port map (
            O => \N__5017\,
            I => \RESETn_c_i\
        );

    \I__792\ : InMux
    port map (
            O => \N__5014\,
            I => \N__5011\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__5011\,
            I => \N__5008\
        );

    \I__790\ : Span4Mux_v
    port map (
            O => \N__5008\,
            I => \N__5005\
        );

    \I__789\ : Sp12to4
    port map (
            O => \N__5005\,
            I => \N__5002\
        );

    \I__788\ : Span12Mux_h
    port map (
            O => \N__5002\,
            I => \N__4999\
        );

    \I__787\ : Span12Mux_v
    port map (
            O => \N__4999\,
            I => \N__4996\
        );

    \I__786\ : Odrv12
    port map (
            O => \N__4996\,
            I => \A_c_7\
        );

    \I__785\ : CascadeMux
    port map (
            O => \N__4993\,
            I => \N__4990\
        );

    \I__784\ : InMux
    port map (
            O => \N__4990\,
            I => \N__4987\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__4987\,
            I => \N__4984\
        );

    \I__782\ : Span4Mux_v
    port map (
            O => \N__4984\,
            I => \N__4981\
        );

    \I__781\ : Sp12to4
    port map (
            O => \N__4981\,
            I => \N__4978\
        );

    \I__780\ : Span12Mux_h
    port map (
            O => \N__4978\,
            I => \N__4975\
        );

    \I__779\ : Odrv12
    port map (
            O => \N__4975\,
            I => \A_c_14\
        );

    \I__778\ : InMux
    port map (
            O => \N__4972\,
            I => \N__4968\
        );

    \I__777\ : InMux
    port map (
            O => \N__4971\,
            I => \N__4965\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__4968\,
            I => \N__4962\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__4965\,
            I => \N__4959\
        );

    \I__774\ : Span4Mux_v
    port map (
            O => \N__4962\,
            I => \N__4954\
        );

    \I__773\ : Span4Mux_v
    port map (
            O => \N__4959\,
            I => \N__4954\
        );

    \I__772\ : Sp12to4
    port map (
            O => \N__4954\,
            I => \N__4951\
        );

    \I__771\ : Span12Mux_h
    port map (
            O => \N__4951\,
            I => \N__4948\
        );

    \I__770\ : Span12Mux_v
    port map (
            O => \N__4948\,
            I => \N__4945\
        );

    \I__769\ : Odrv12
    port map (
            O => \N__4945\,
            I => \DRA_c_2\
        );

    \I__768\ : InMux
    port map (
            O => \N__4942\,
            I => \N__4939\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__4939\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__766\ : InMux
    port map (
            O => \N__4936\,
            I => \N__4932\
        );

    \I__765\ : InMux
    port map (
            O => \N__4935\,
            I => \N__4929\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__4932\,
            I => \N__4924\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__4929\,
            I => \N__4924\
        );

    \I__762\ : Span12Mux_v
    port map (
            O => \N__4924\,
            I => \N__4921\
        );

    \I__761\ : Span12Mux_h
    port map (
            O => \N__4921\,
            I => \N__4918\
        );

    \I__760\ : Odrv12
    port map (
            O => \N__4918\,
            I => \DRA_c_4\
        );

    \I__759\ : CascadeMux
    port map (
            O => \N__4915\,
            I => \U712_CHIP_RAM.N_341_cascade_\
        );

    \I__758\ : CascadeMux
    port map (
            O => \N__4912\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_1_1_cascade_\
        );

    \I__757\ : InMux
    port map (
            O => \N__4909\,
            I => \N__4905\
        );

    \I__756\ : InMux
    port map (
            O => \N__4908\,
            I => \N__4902\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__4905\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__4902\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__753\ : InMux
    port map (
            O => \N__4897\,
            I => \N__4893\
        );

    \I__752\ : InMux
    port map (
            O => \N__4896\,
            I => \N__4890\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__4893\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__4890\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__749\ : CascadeMux
    port map (
            O => \N__4885\,
            I => \N__4881\
        );

    \I__748\ : InMux
    port map (
            O => \N__4884\,
            I => \N__4878\
        );

    \I__747\ : InMux
    port map (
            O => \N__4881\,
            I => \N__4875\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__4878\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__4875\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__744\ : InMux
    port map (
            O => \N__4870\,
            I => \N__4866\
        );

    \I__743\ : InMux
    port map (
            O => \N__4869\,
            I => \N__4863\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__4866\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__4863\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__740\ : InMux
    port map (
            O => \N__4858\,
            I => \N__4854\
        );

    \I__739\ : InMux
    port map (
            O => \N__4857\,
            I => \N__4851\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__4854\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__4851\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__736\ : InMux
    port map (
            O => \N__4846\,
            I => \N__4842\
        );

    \I__735\ : InMux
    port map (
            O => \N__4845\,
            I => \N__4839\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__4842\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__4839\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__732\ : CascadeMux
    port map (
            O => \N__4834\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0_cascade_\
        );

    \I__731\ : InMux
    port map (
            O => \N__4831\,
            I => \N__4828\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__4828\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\
        );

    \I__729\ : CascadeMux
    port map (
            O => \N__4825\,
            I => \N__4821\
        );

    \I__728\ : CascadeMux
    port map (
            O => \N__4824\,
            I => \N__4818\
        );

    \I__727\ : InMux
    port map (
            O => \N__4821\,
            I => \N__4815\
        );

    \I__726\ : InMux
    port map (
            O => \N__4818\,
            I => \N__4812\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__4815\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__4812\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__723\ : CascadeMux
    port map (
            O => \N__4807\,
            I => \U712_CYCLE_TERM.N_305_i_0_en_cascade_\
        );

    \I__722\ : InMux
    port map (
            O => \N__4804\,
            I => \N__4800\
        );

    \I__721\ : InMux
    port map (
            O => \N__4803\,
            I => \N__4797\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__4800\,
            I => \N__4792\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__4797\,
            I => \N__4792\
        );

    \I__718\ : Span12Mux_v
    port map (
            O => \N__4792\,
            I => \N__4789\
        );

    \I__717\ : Span12Mux_v
    port map (
            O => \N__4789\,
            I => \N__4786\
        );

    \I__716\ : Span12Mux_h
    port map (
            O => \N__4786\,
            I => \N__4783\
        );

    \I__715\ : Odrv12
    port map (
            O => \N__4783\,
            I => \DRA_c_0\
        );

    \I__714\ : InMux
    port map (
            O => \N__4780\,
            I => \N__4777\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__4777\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__712\ : InMux
    port map (
            O => \N__4774\,
            I => \N__4771\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__4771\,
            I => \N__4767\
        );

    \I__710\ : InMux
    port map (
            O => \N__4770\,
            I => \N__4764\
        );

    \I__709\ : Span4Mux_v
    port map (
            O => \N__4767\,
            I => \N__4761\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__4764\,
            I => \N__4758\
        );

    \I__707\ : Span4Mux_h
    port map (
            O => \N__4761\,
            I => \N__4753\
        );

    \I__706\ : Span4Mux_v
    port map (
            O => \N__4758\,
            I => \N__4753\
        );

    \I__705\ : Sp12to4
    port map (
            O => \N__4753\,
            I => \N__4750\
        );

    \I__704\ : Span12Mux_h
    port map (
            O => \N__4750\,
            I => \N__4747\
        );

    \I__703\ : Span12Mux_v
    port map (
            O => \N__4747\,
            I => \N__4744\
        );

    \I__702\ : Odrv12
    port map (
            O => \N__4744\,
            I => \DRA_c_1\
        );

    \I__701\ : InMux
    port map (
            O => \N__4741\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__700\ : InMux
    port map (
            O => \N__4738\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__699\ : InMux
    port map (
            O => \N__4735\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__698\ : InMux
    port map (
            O => \N__4732\,
            I => \N__4728\
        );

    \I__697\ : InMux
    port map (
            O => \N__4731\,
            I => \N__4725\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__4728\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__4725\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__694\ : InMux
    port map (
            O => \N__4720\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__693\ : InMux
    port map (
            O => \N__4717\,
            I => \N__4713\
        );

    \I__692\ : InMux
    port map (
            O => \N__4716\,
            I => \N__4710\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__4713\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__4710\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__689\ : InMux
    port map (
            O => \N__4705\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__688\ : InMux
    port map (
            O => \N__4702\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__687\ : ClkMux
    port map (
            O => \N__4699\,
            I => \N__4696\
        );

    \I__686\ : GlobalMux
    port map (
            O => \N__4696\,
            I => \N__4693\
        );

    \I__685\ : gio2CtrlBuf
    port map (
            O => \N__4693\,
            I => \C1_c_g\
        );

    \I__684\ : InMux
    port map (
            O => \N__4690\,
            I => \N__4686\
        );

    \I__683\ : InMux
    port map (
            O => \N__4689\,
            I => \N__4683\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__4686\,
            I => \U712_REG_SM.N_306\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__4683\,
            I => \U712_REG_SM.N_306\
        );

    \I__680\ : CascadeMux
    port map (
            O => \N__4678\,
            I => \N__4675\
        );

    \I__679\ : InMux
    port map (
            O => \N__4675\,
            I => \N__4669\
        );

    \I__678\ : InMux
    port map (
            O => \N__4674\,
            I => \N__4666\
        );

    \I__677\ : InMux
    port map (
            O => \N__4673\,
            I => \N__4661\
        );

    \I__676\ : InMux
    port map (
            O => \N__4672\,
            I => \N__4661\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__4669\,
            I => \N__4658\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__4666\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__4661\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__672\ : Odrv4
    port map (
            O => \N__4658\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__671\ : InMux
    port map (
            O => \N__4651\,
            I => \N__4646\
        );

    \I__670\ : InMux
    port map (
            O => \N__4650\,
            I => \N__4641\
        );

    \I__669\ : InMux
    port map (
            O => \N__4649\,
            I => \N__4641\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__4646\,
            I => \U712_REG_SM.N_298\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__4641\,
            I => \U712_REG_SM.N_298\
        );

    \I__666\ : CascadeMux
    port map (
            O => \N__4636\,
            I => \N__4633\
        );

    \I__665\ : InMux
    port map (
            O => \N__4633\,
            I => \N__4629\
        );

    \I__664\ : InMux
    port map (
            O => \N__4632\,
            I => \N__4625\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__4629\,
            I => \N__4622\
        );

    \I__662\ : InMux
    port map (
            O => \N__4628\,
            I => \N__4619\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__4625\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__660\ : Odrv4
    port map (
            O => \N__4622\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__4619\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__658\ : InMux
    port map (
            O => \N__4612\,
            I => \N__4608\
        );

    \I__657\ : CascadeMux
    port map (
            O => \N__4611\,
            I => \N__4605\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__4608\,
            I => \N__4602\
        );

    \I__655\ : InMux
    port map (
            O => \N__4605\,
            I => \N__4599\
        );

    \I__654\ : Odrv4
    port map (
            O => \N__4602\,
            I => \U712_REG_SM.UDS_OUTZ0\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__4599\,
            I => \U712_REG_SM.UDS_OUTZ0\
        );

    \I__652\ : IoInMux
    port map (
            O => \N__4594\,
            I => \N__4591\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__4591\,
            I => \N__4588\
        );

    \I__650\ : Span12Mux_s4_v
    port map (
            O => \N__4588\,
            I => \N__4585\
        );

    \I__649\ : Span12Mux_h
    port map (
            O => \N__4585\,
            I => \N__4582\
        );

    \I__648\ : Odrv12
    port map (
            O => \N__4582\,
            I => \U712_REG_SM_un1_UDSn_i\
        );

    \I__647\ : InMux
    port map (
            O => \N__4579\,
            I => \N__4567\
        );

    \I__646\ : InMux
    port map (
            O => \N__4578\,
            I => \N__4567\
        );

    \I__645\ : InMux
    port map (
            O => \N__4577\,
            I => \N__4567\
        );

    \I__644\ : InMux
    port map (
            O => \N__4576\,
            I => \N__4567\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__4567\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__642\ : CascadeMux
    port map (
            O => \N__4564\,
            I => \N__4560\
        );

    \I__641\ : InMux
    port map (
            O => \N__4563\,
            I => \N__4554\
        );

    \I__640\ : InMux
    port map (
            O => \N__4560\,
            I => \N__4554\
        );

    \I__639\ : InMux
    port map (
            O => \N__4559\,
            I => \N__4551\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__4554\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__4551\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__636\ : InMux
    port map (
            O => \N__4546\,
            I => \N__4542\
        );

    \I__635\ : InMux
    port map (
            O => \N__4545\,
            I => \N__4539\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__4542\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__4539\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__632\ : InMux
    port map (
            O => \N__4534\,
            I => \N__4531\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__4531\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\
        );

    \I__630\ : IoInMux
    port map (
            O => \N__4528\,
            I => \N__4525\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__4525\,
            I => \N__4522\
        );

    \I__628\ : IoSpan4Mux
    port map (
            O => \N__4522\,
            I => \N__4519\
        );

    \I__627\ : Span4Mux_s3_h
    port map (
            O => \N__4519\,
            I => \N__4516\
        );

    \I__626\ : Span4Mux_h
    port map (
            O => \N__4516\,
            I => \N__4513\
        );

    \I__625\ : Span4Mux_h
    port map (
            O => \N__4513\,
            I => \N__4510\
        );

    \I__624\ : Odrv4
    port map (
            O => \N__4510\,
            I => \N_886_i\
        );

    \I__623\ : InMux
    port map (
            O => \N__4507\,
            I => \N__4504\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__4504\,
            I => \N__4501\
        );

    \I__621\ : Span4Mux_v
    port map (
            O => \N__4501\,
            I => \N__4498\
        );

    \I__620\ : Sp12to4
    port map (
            O => \N__4498\,
            I => \N__4495\
        );

    \I__619\ : Span12Mux_h
    port map (
            O => \N__4495\,
            I => \N__4492\
        );

    \I__618\ : Span12Mux_v
    port map (
            O => \N__4492\,
            I => \N__4489\
        );

    \I__617\ : Odrv12
    port map (
            O => \N__4489\,
            I => \A_c_4\
        );

    \I__616\ : CascadeMux
    port map (
            O => \N__4486\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_2_cascade_\
        );

    \I__615\ : InMux
    port map (
            O => \N__4483\,
            I => \N__4480\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__4480\,
            I => \N__4477\
        );

    \I__613\ : Span12Mux_h
    port map (
            O => \N__4477\,
            I => \N__4474\
        );

    \I__612\ : Odrv12
    port map (
            O => \N__4474\,
            I => \A_c_11\
        );

    \I__611\ : InMux
    port map (
            O => \N__4471\,
            I => \bfn_11_9_0_\
        );

    \I__610\ : InMux
    port map (
            O => \N__4468\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__609\ : InMux
    port map (
            O => \N__4465\,
            I => \N__4462\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__4462\,
            I => \N__4456\
        );

    \I__607\ : InMux
    port map (
            O => \N__4461\,
            I => \N__4453\
        );

    \I__606\ : InMux
    port map (
            O => \N__4460\,
            I => \N__4448\
        );

    \I__605\ : InMux
    port map (
            O => \N__4459\,
            I => \N__4448\
        );

    \I__604\ : Odrv4
    port map (
            O => \N__4456\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__4453\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__4448\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__601\ : InMux
    port map (
            O => \N__4441\,
            I => \N__4437\
        );

    \I__600\ : InMux
    port map (
            O => \N__4440\,
            I => \N__4431\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__4437\,
            I => \N__4428\
        );

    \I__598\ : InMux
    port map (
            O => \N__4436\,
            I => \N__4425\
        );

    \I__597\ : InMux
    port map (
            O => \N__4435\,
            I => \N__4420\
        );

    \I__596\ : InMux
    port map (
            O => \N__4434\,
            I => \N__4420\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__4431\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__594\ : Odrv4
    port map (
            O => \N__4428\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__4425\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__4420\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__591\ : CascadeMux
    port map (
            O => \N__4411\,
            I => \N__4407\
        );

    \I__590\ : CascadeMux
    port map (
            O => \N__4410\,
            I => \N__4404\
        );

    \I__589\ : InMux
    port map (
            O => \N__4407\,
            I => \N__4399\
        );

    \I__588\ : InMux
    port map (
            O => \N__4404\,
            I => \N__4399\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__4399\,
            I => \U712_REG_SM.N_289\
        );

    \I__586\ : InMux
    port map (
            O => \N__4396\,
            I => \N__4392\
        );

    \I__585\ : InMux
    port map (
            O => \N__4395\,
            I => \N__4389\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__4392\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__4389\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__582\ : InMux
    port map (
            O => \N__4384\,
            I => \N__4375\
        );

    \I__581\ : InMux
    port map (
            O => \N__4383\,
            I => \N__4368\
        );

    \I__580\ : InMux
    port map (
            O => \N__4382\,
            I => \N__4368\
        );

    \I__579\ : InMux
    port map (
            O => \N__4381\,
            I => \N__4368\
        );

    \I__578\ : InMux
    port map (
            O => \N__4380\,
            I => \N__4361\
        );

    \I__577\ : InMux
    port map (
            O => \N__4379\,
            I => \N__4361\
        );

    \I__576\ : InMux
    port map (
            O => \N__4378\,
            I => \N__4361\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__4375\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__4368\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__4361\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__572\ : CascadeMux
    port map (
            O => \N__4354\,
            I => \U712_REG_SM.N_289_cascade_\
        );

    \I__571\ : InMux
    port map (
            O => \N__4351\,
            I => \N__4341\
        );

    \I__570\ : InMux
    port map (
            O => \N__4350\,
            I => \N__4341\
        );

    \I__569\ : InMux
    port map (
            O => \N__4349\,
            I => \N__4336\
        );

    \I__568\ : InMux
    port map (
            O => \N__4348\,
            I => \N__4331\
        );

    \I__567\ : InMux
    port map (
            O => \N__4347\,
            I => \N__4331\
        );

    \I__566\ : InMux
    port map (
            O => \N__4346\,
            I => \N__4328\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__4341\,
            I => \N__4325\
        );

    \I__564\ : InMux
    port map (
            O => \N__4340\,
            I => \N__4320\
        );

    \I__563\ : InMux
    port map (
            O => \N__4339\,
            I => \N__4320\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__4336\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__4331\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__4328\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__559\ : Odrv4
    port map (
            O => \N__4325\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__4320\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__557\ : InMux
    port map (
            O => \N__4309\,
            I => \N__4303\
        );

    \I__556\ : InMux
    port map (
            O => \N__4308\,
            I => \N__4303\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__4303\,
            I => \U712_REG_SM.N_494\
        );

    \I__554\ : CascadeMux
    port map (
            O => \N__4300\,
            I => \N__4296\
        );

    \I__553\ : InMux
    port map (
            O => \N__4299\,
            I => \N__4288\
        );

    \I__552\ : InMux
    port map (
            O => \N__4296\,
            I => \N__4288\
        );

    \I__551\ : InMux
    port map (
            O => \N__4295\,
            I => \N__4281\
        );

    \I__550\ : InMux
    port map (
            O => \N__4294\,
            I => \N__4281\
        );

    \I__549\ : InMux
    port map (
            O => \N__4293\,
            I => \N__4281\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__4288\,
            I => \U712_REG_SM.N_288\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4281\,
            I => \U712_REG_SM.N_288\
        );

    \I__546\ : CascadeMux
    port map (
            O => \N__4276\,
            I => \U712_REG_SM.N_494_cascade_\
        );

    \I__545\ : InMux
    port map (
            O => \N__4273\,
            I => \N__4269\
        );

    \I__544\ : InMux
    port map (
            O => \N__4272\,
            I => \N__4266\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__4269\,
            I => \U712_REG_SM.N_424\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__4266\,
            I => \U712_REG_SM.N_424\
        );

    \I__541\ : InMux
    port map (
            O => \N__4261\,
            I => \N__4258\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__4258\,
            I => \U712_REG_SM.N_369\
        );

    \I__539\ : CascadeMux
    port map (
            O => \N__4255\,
            I => \U712_REG_SM.DS_EN_RNOZ0Z_2_cascade_\
        );

    \I__538\ : InMux
    port map (
            O => \N__4252\,
            I => \N__4249\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__4249\,
            I => \U712_REG_SM.N_123\
        );

    \I__536\ : IoInMux
    port map (
            O => \N__4246\,
            I => \N__4243\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__4243\,
            I => \N__4240\
        );

    \I__534\ : Span12Mux_s1_h
    port map (
            O => \N__4240\,
            I => \N__4237\
        );

    \I__533\ : Span12Mux_h
    port map (
            O => \N__4237\,
            I => \N__4233\
        );

    \I__532\ : InMux
    port map (
            O => \N__4236\,
            I => \N__4230\
        );

    \I__531\ : Odrv12
    port map (
            O => \N__4233\,
            I => \TACK_OUTn\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__4230\,
            I => \TACK_OUTn\
        );

    \I__529\ : InMux
    port map (
            O => \N__4225\,
            I => \N__4222\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__4222\,
            I => \N__4216\
        );

    \I__527\ : InMux
    port map (
            O => \N__4221\,
            I => \N__4209\
        );

    \I__526\ : InMux
    port map (
            O => \N__4220\,
            I => \N__4209\
        );

    \I__525\ : InMux
    port map (
            O => \N__4219\,
            I => \N__4209\
        );

    \I__524\ : Span4Mux_v
    port map (
            O => \N__4216\,
            I => \N__4204\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__4209\,
            I => \N__4204\
        );

    \I__522\ : Span4Mux_h
    port map (
            O => \N__4204\,
            I => \N__4201\
        );

    \I__521\ : Sp12to4
    port map (
            O => \N__4201\,
            I => \N__4198\
        );

    \I__520\ : Span12Mux_v
    port map (
            O => \N__4198\,
            I => \N__4195\
        );

    \I__519\ : Odrv12
    port map (
            O => \N__4195\,
            I => \CLK40_OUT_i\
        );

    \I__518\ : InMux
    port map (
            O => \N__4192\,
            I => \N__4189\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__4189\,
            I => \U712_BYTE_ENABLE.N_395\
        );

    \I__516\ : IoInMux
    port map (
            O => \N__4186\,
            I => \N__4183\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__4183\,
            I => \N__4180\
        );

    \I__514\ : IoSpan4Mux
    port map (
            O => \N__4180\,
            I => \N__4177\
        );

    \I__513\ : Span4Mux_s3_h
    port map (
            O => \N__4177\,
            I => \N__4174\
        );

    \I__512\ : Sp12to4
    port map (
            O => \N__4174\,
            I => \N__4171\
        );

    \I__511\ : Span12Mux_s8_h
    port map (
            O => \N__4171\,
            I => \N__4168\
        );

    \I__510\ : Span12Mux_v
    port map (
            O => \N__4168\,
            I => \N__4165\
        );

    \I__509\ : Odrv12
    port map (
            O => \N__4165\,
            I => \N_74_i\
        );

    \I__508\ : InMux
    port map (
            O => \N__4162\,
            I => \N__4153\
        );

    \I__507\ : InMux
    port map (
            O => \N__4161\,
            I => \N__4153\
        );

    \I__506\ : InMux
    port map (
            O => \N__4160\,
            I => \N__4153\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4153\,
            I => \U712_BYTE_ENABLE.N_387\
        );

    \I__504\ : InMux
    port map (
            O => \N__4150\,
            I => \N__4140\
        );

    \I__503\ : InMux
    port map (
            O => \N__4149\,
            I => \N__4140\
        );

    \I__502\ : InMux
    port map (
            O => \N__4148\,
            I => \N__4140\
        );

    \I__501\ : InMux
    port map (
            O => \N__4147\,
            I => \N__4137\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4140\,
            I => \N__4132\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__4137\,
            I => \N__4132\
        );

    \I__498\ : Span4Mux_h
    port map (
            O => \N__4132\,
            I => \N__4129\
        );

    \I__497\ : Sp12to4
    port map (
            O => \N__4129\,
            I => \N__4126\
        );

    \I__496\ : Span12Mux_v
    port map (
            O => \N__4126\,
            I => \N__4123\
        );

    \I__495\ : Odrv12
    port map (
            O => \N__4123\,
            I => \A_c_1\
        );

    \I__494\ : CascadeMux
    port map (
            O => \N__4120\,
            I => \N__4117\
        );

    \I__493\ : InMux
    port map (
            O => \N__4117\,
            I => \N__4111\
        );

    \I__492\ : InMux
    port map (
            O => \N__4116\,
            I => \N__4111\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__4111\,
            I => \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_0_0\
        );

    \I__490\ : IoInMux
    port map (
            O => \N__4108\,
            I => \N__4105\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__4105\,
            I => \N__4102\
        );

    \I__488\ : Span12Mux_s6_h
    port map (
            O => \N__4102\,
            I => \N__4099\
        );

    \I__487\ : Span12Mux_h
    port map (
            O => \N__4099\,
            I => \N__4096\
        );

    \I__486\ : Odrv12
    port map (
            O => \N__4096\,
            I => \N_76_i\
        );

    \I__485\ : CascadeMux
    port map (
            O => \N__4093\,
            I => \N__4090\
        );

    \I__484\ : InMux
    port map (
            O => \N__4090\,
            I => \N__4087\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__4087\,
            I => \U712_BYTE_ENABLE.N_391\
        );

    \I__482\ : InMux
    port map (
            O => \N__4084\,
            I => \N__4080\
        );

    \I__481\ : InMux
    port map (
            O => \N__4083\,
            I => \N__4077\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__4080\,
            I => \U712_REG_SM.N_304\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4077\,
            I => \U712_REG_SM.N_304\
        );

    \I__478\ : CascadeMux
    port map (
            O => \N__4072\,
            I => \N__4068\
        );

    \I__477\ : InMux
    port map (
            O => \N__4071\,
            I => \N__4060\
        );

    \I__476\ : InMux
    port map (
            O => \N__4068\,
            I => \N__4060\
        );

    \I__475\ : InMux
    port map (
            O => \N__4067\,
            I => \N__4060\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__4060\,
            I => \U712_REG_SM.N_299\
        );

    \I__473\ : InMux
    port map (
            O => \N__4057\,
            I => \N__4048\
        );

    \I__472\ : InMux
    port map (
            O => \N__4056\,
            I => \N__4048\
        );

    \I__471\ : InMux
    port map (
            O => \N__4055\,
            I => \N__4048\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__4048\,
            I => \U712_REG_SM.N_281\
        );

    \I__469\ : InMux
    port map (
            O => \N__4045\,
            I => \N__4040\
        );

    \I__468\ : InMux
    port map (
            O => \N__4044\,
            I => \N__4037\
        );

    \I__467\ : InMux
    port map (
            O => \N__4043\,
            I => \N__4034\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__4040\,
            I => \U712_REG_SM.N_280\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__4037\,
            I => \U712_REG_SM.N_280\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__4034\,
            I => \U712_REG_SM.N_280\
        );

    \I__463\ : CascadeMux
    port map (
            O => \N__4027\,
            I => \U712_REG_SM.N_373_cascade_\
        );

    \I__462\ : CascadeMux
    port map (
            O => \N__4024\,
            I => \U712_REG_SM.N_288_cascade_\
        );

    \I__461\ : InMux
    port map (
            O => \N__4021\,
            I => \N__4014\
        );

    \I__460\ : InMux
    port map (
            O => \N__4020\,
            I => \N__4014\
        );

    \I__459\ : InMux
    port map (
            O => \N__4019\,
            I => \N__4011\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__4014\,
            I => \U712_REG_SM.N_307\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__4011\,
            I => \U712_REG_SM.N_307\
        );

    \I__456\ : CascadeMux
    port map (
            O => \N__4006\,
            I => \N__4003\
        );

    \I__455\ : InMux
    port map (
            O => \N__4003\,
            I => \N__3999\
        );

    \I__454\ : InMux
    port map (
            O => \N__4002\,
            I => \N__3996\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__3999\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__3996\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__451\ : InMux
    port map (
            O => \N__3991\,
            I => \N__3988\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__3988\,
            I => \N__3985\
        );

    \I__449\ : Span4Mux_v
    port map (
            O => \N__3985\,
            I => \N__3982\
        );

    \I__448\ : Sp12to4
    port map (
            O => \N__3982\,
            I => \N__3979\
        );

    \I__447\ : Span12Mux_h
    port map (
            O => \N__3979\,
            I => \N__3976\
        );

    \I__446\ : Odrv12
    port map (
            O => \N__3976\,
            I => \C3_c\
        );

    \I__445\ : IoInMux
    port map (
            O => \N__3973\,
            I => \N__3969\
        );

    \I__444\ : InMux
    port map (
            O => \N__3972\,
            I => \N__3966\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__3969\,
            I => \N__3963\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__3966\,
            I => \N__3960\
        );

    \I__441\ : Span4Mux_s3_h
    port map (
            O => \N__3963\,
            I => \N__3957\
        );

    \I__440\ : Span12Mux_h
    port map (
            O => \N__3960\,
            I => \N__3952\
        );

    \I__439\ : Sp12to4
    port map (
            O => \N__3957\,
            I => \N__3952\
        );

    \I__438\ : Span12Mux_v
    port map (
            O => \N__3952\,
            I => \N__3949\
        );

    \I__437\ : Odrv12
    port map (
            O => \N__3949\,
            I => \C1_c\
        );

    \I__436\ : InMux
    port map (
            O => \N__3946\,
            I => \N__3940\
        );

    \I__435\ : InMux
    port map (
            O => \N__3945\,
            I => \N__3933\
        );

    \I__434\ : InMux
    port map (
            O => \N__3944\,
            I => \N__3933\
        );

    \I__433\ : InMux
    port map (
            O => \N__3943\,
            I => \N__3933\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__3940\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__3933\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__430\ : InMux
    port map (
            O => \N__3928\,
            I => \N__3924\
        );

    \I__429\ : InMux
    port map (
            O => \N__3927\,
            I => \N__3921\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__3924\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2Z0Z_0\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__3921\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2Z0Z_0\
        );

    \I__426\ : IoInMux
    port map (
            O => \N__3916\,
            I => \N__3913\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__3913\,
            I => \N__3910\
        );

    \I__424\ : Span4Mux_s2_h
    port map (
            O => \N__3910\,
            I => \N__3907\
        );

    \I__423\ : Span4Mux_h
    port map (
            O => \N__3907\,
            I => \N__3904\
        );

    \I__422\ : Sp12to4
    port map (
            O => \N__3904\,
            I => \N__3901\
        );

    \I__421\ : Span12Mux_s11_v
    port map (
            O => \N__3901\,
            I => \N__3898\
        );

    \I__420\ : Span12Mux_h
    port map (
            O => \N__3898\,
            I => \N__3895\
        );

    \I__419\ : Odrv12
    port map (
            O => \N__3895\,
            I => \N_75_i\
        );

    \I__418\ : InMux
    port map (
            O => \N__3892\,
            I => \N__3886\
        );

    \I__417\ : InMux
    port map (
            O => \N__3891\,
            I => \N__3886\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__3886\,
            I => \U712_REG_SM.N_301\
        );

    \I__415\ : InMux
    port map (
            O => \N__3883\,
            I => \N__3877\
        );

    \I__414\ : InMux
    port map (
            O => \N__3882\,
            I => \N__3877\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__3877\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__412\ : IoInMux
    port map (
            O => \N__3874\,
            I => \N__3870\
        );

    \I__411\ : IoInMux
    port map (
            O => \N__3873\,
            I => \N__3867\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__3870\,
            I => \N__3864\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__3867\,
            I => \N__3861\
        );

    \I__408\ : IoSpan4Mux
    port map (
            O => \N__3864\,
            I => \N__3858\
        );

    \I__407\ : IoSpan4Mux
    port map (
            O => \N__3861\,
            I => \N__3855\
        );

    \I__406\ : Span4Mux_s3_v
    port map (
            O => \N__3858\,
            I => \N__3852\
        );

    \I__405\ : Span4Mux_s3_v
    port map (
            O => \N__3855\,
            I => \N__3849\
        );

    \I__404\ : Sp12to4
    port map (
            O => \N__3852\,
            I => \N__3846\
        );

    \I__403\ : Sp12to4
    port map (
            O => \N__3849\,
            I => \N__3843\
        );

    \I__402\ : Span12Mux_s9_h
    port map (
            O => \N__3846\,
            I => \N__3839\
        );

    \I__401\ : Span12Mux_s10_h
    port map (
            O => \N__3843\,
            I => \N__3836\
        );

    \I__400\ : CascadeMux
    port map (
            O => \N__3842\,
            I => \N__3833\
        );

    \I__399\ : Span12Mux_v
    port map (
            O => \N__3839\,
            I => \N__3828\
        );

    \I__398\ : Span12Mux_v
    port map (
            O => \N__3836\,
            I => \N__3828\
        );

    \I__397\ : InMux
    port map (
            O => \N__3833\,
            I => \N__3825\
        );

    \I__396\ : Odrv12
    port map (
            O => \N__3828\,
            I => \ASn_c\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__3825\,
            I => \ASn_c\
        );

    \I__394\ : InMux
    port map (
            O => \N__3820\,
            I => \N__3815\
        );

    \I__393\ : InMux
    port map (
            O => \N__3819\,
            I => \N__3810\
        );

    \I__392\ : InMux
    port map (
            O => \N__3818\,
            I => \N__3810\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__3815\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__3810\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__389\ : CascadeMux
    port map (
            O => \N__3805\,
            I => \N__3802\
        );

    \I__388\ : InMux
    port map (
            O => \N__3802\,
            I => \N__3795\
        );

    \I__387\ : InMux
    port map (
            O => \N__3801\,
            I => \N__3795\
        );

    \I__386\ : InMux
    port map (
            O => \N__3800\,
            I => \N__3792\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__3795\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__3792\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__383\ : CascadeMux
    port map (
            O => \N__3787\,
            I => \U712_REG_SM.N_281_cascade_\
        );

    \I__382\ : CascadeMux
    port map (
            O => \N__3784\,
            I => \U712_REG_SM.N_280_cascade_\
        );

    \I__381\ : CascadeMux
    port map (
            O => \N__3781\,
            I => \N__3777\
        );

    \I__380\ : CascadeMux
    port map (
            O => \N__3780\,
            I => \N__3774\
        );

    \I__379\ : InMux
    port map (
            O => \N__3777\,
            I => \N__3769\
        );

    \I__378\ : InMux
    port map (
            O => \N__3774\,
            I => \N__3766\
        );

    \I__377\ : InMux
    port map (
            O => \N__3773\,
            I => \N__3761\
        );

    \I__376\ : InMux
    port map (
            O => \N__3772\,
            I => \N__3761\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__3769\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__3766\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__3761\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__372\ : InMux
    port map (
            O => \N__3754\,
            I => \N__3748\
        );

    \I__371\ : InMux
    port map (
            O => \N__3753\,
            I => \N__3748\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__3748\,
            I => \U712_REG_SM.N_308\
        );

    \I__369\ : InMux
    port map (
            O => \N__3745\,
            I => \N__3742\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__3742\,
            I => \N__3739\
        );

    \I__367\ : Span4Mux_v
    port map (
            O => \N__3739\,
            I => \N__3735\
        );

    \I__366\ : InMux
    port map (
            O => \N__3738\,
            I => \N__3732\
        );

    \I__365\ : Sp12to4
    port map (
            O => \N__3735\,
            I => \N__3727\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__3732\,
            I => \N__3727\
        );

    \I__363\ : Span12Mux_h
    port map (
            O => \N__3727\,
            I => \N__3724\
        );

    \I__362\ : Span12Mux_v
    port map (
            O => \N__3724\,
            I => \N__3721\
        );

    \I__361\ : Odrv12
    port map (
            O => \N__3721\,
            I => \SIZ_c_0\
        );

    \I__360\ : CascadeMux
    port map (
            O => \N__3718\,
            I => \U712_BYTE_ENABLE.N_387_cascade_\
        );

    \I__359\ : IoInMux
    port map (
            O => \N__3715\,
            I => \N__3712\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__3712\,
            I => \N__3709\
        );

    \I__357\ : Span4Mux_s2_v
    port map (
            O => \N__3709\,
            I => \N__3706\
        );

    \I__356\ : Span4Mux_v
    port map (
            O => \N__3706\,
            I => \N__3703\
        );

    \I__355\ : Span4Mux_v
    port map (
            O => \N__3703\,
            I => \N__3700\
        );

    \I__354\ : Span4Mux_v
    port map (
            O => \N__3700\,
            I => \N__3697\
        );

    \I__353\ : Odrv4
    port map (
            O => \N__3697\,
            I => \N_73_i\
        );

    \I__352\ : InMux
    port map (
            O => \N__3694\,
            I => \N__3690\
        );

    \I__351\ : InMux
    port map (
            O => \N__3693\,
            I => \N__3687\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__3690\,
            I => \N__3682\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__3687\,
            I => \N__3682\
        );

    \I__348\ : Span4Mux_v
    port map (
            O => \N__3682\,
            I => \N__3677\
        );

    \I__347\ : InMux
    port map (
            O => \N__3681\,
            I => \N__3672\
        );

    \I__346\ : InMux
    port map (
            O => \N__3680\,
            I => \N__3672\
        );

    \I__345\ : Span4Mux_v
    port map (
            O => \N__3677\,
            I => \N__3669\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__3672\,
            I => \N__3666\
        );

    \I__343\ : Sp12to4
    port map (
            O => \N__3669\,
            I => \N__3661\
        );

    \I__342\ : Span12Mux_v
    port map (
            O => \N__3666\,
            I => \N__3661\
        );

    \I__341\ : Odrv12
    port map (
            O => \N__3661\,
            I => \A_c_0\
        );

    \I__340\ : InMux
    port map (
            O => \N__3658\,
            I => \N__3655\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__3655\,
            I => \N__3651\
        );

    \I__338\ : InMux
    port map (
            O => \N__3654\,
            I => \N__3648\
        );

    \I__337\ : Span4Mux_v
    port map (
            O => \N__3651\,
            I => \N__3643\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__3648\,
            I => \N__3643\
        );

    \I__335\ : Span4Mux_h
    port map (
            O => \N__3643\,
            I => \N__3640\
        );

    \I__334\ : Sp12to4
    port map (
            O => \N__3640\,
            I => \N__3637\
        );

    \I__333\ : Span12Mux_v
    port map (
            O => \N__3637\,
            I => \N__3634\
        );

    \I__332\ : Odrv12
    port map (
            O => \N__3634\,
            I => \SIZ_c_1\
        );

    \I__331\ : InMux
    port map (
            O => \N__3631\,
            I => \N__3628\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__3628\,
            I => \N__3625\
        );

    \I__329\ : Span4Mux_v
    port map (
            O => \N__3625\,
            I => \N__3622\
        );

    \I__328\ : Sp12to4
    port map (
            O => \N__3622\,
            I => \N__3619\
        );

    \I__327\ : Span12Mux_h
    port map (
            O => \N__3619\,
            I => \N__3616\
        );

    \I__326\ : Span12Mux_v
    port map (
            O => \N__3616\,
            I => \N__3613\
        );

    \I__325\ : Odrv12
    port map (
            O => \N__3613\,
            I => \REGSPACEn_c\
        );

    \I__324\ : IoInMux
    port map (
            O => \N__3610\,
            I => \N__3607\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__3607\,
            I => \N__3604\
        );

    \I__322\ : Span4Mux_s3_v
    port map (
            O => \N__3604\,
            I => \N__3601\
        );

    \I__321\ : Span4Mux_h
    port map (
            O => \N__3601\,
            I => \N__3598\
        );

    \I__320\ : Odrv4
    port map (
            O => \N__3598\,
            I => \CLK80_OUT_i_i\
        );

    \I__319\ : IoInMux
    port map (
            O => \N__3595\,
            I => \N__3592\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__3592\,
            I => \N__3589\
        );

    \I__317\ : Span12Mux_s6_h
    port map (
            O => \N__3589\,
            I => \N__3586\
        );

    \I__316\ : Odrv12
    port map (
            O => \N__3586\,
            I => \CLK40_OUT_i_i\
        );

    \I__315\ : CascadeMux
    port map (
            O => \N__3583\,
            I => \N__3579\
        );

    \I__314\ : InMux
    port map (
            O => \N__3582\,
            I => \N__3574\
        );

    \I__313\ : InMux
    port map (
            O => \N__3579\,
            I => \N__3574\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__3574\,
            I => \U712_REG_SM.LDS_OUT_2_0_a2Z0Z_0\
        );

    \I__311\ : IoInMux
    port map (
            O => \N__3571\,
            I => \N__3568\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__3568\,
            I => \N__3565\
        );

    \I__309\ : Span4Mux_s1_v
    port map (
            O => \N__3565\,
            I => \N__3562\
        );

    \I__308\ : Span4Mux_v
    port map (
            O => \N__3562\,
            I => \N__3559\
        );

    \I__307\ : Span4Mux_v
    port map (
            O => \N__3559\,
            I => \N__3556\
        );

    \I__306\ : Odrv4
    port map (
            O => \N__3556\,
            I => \VBENn_c\
        );

    \I__305\ : IoInMux
    port map (
            O => \N__3553\,
            I => \N__3550\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__3550\,
            I => \N__3547\
        );

    \I__303\ : IoSpan4Mux
    port map (
            O => \N__3547\,
            I => \N__3544\
        );

    \I__302\ : Span4Mux_s2_v
    port map (
            O => \N__3544\,
            I => \N__3541\
        );

    \I__301\ : Sp12to4
    port map (
            O => \N__3541\,
            I => \N__3538\
        );

    \I__300\ : Span12Mux_v
    port map (
            O => \N__3538\,
            I => \N__3535\
        );

    \I__299\ : Odrv12
    port map (
            O => \N__3535\,
            I => \CLK40_IN_c\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_9_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5023\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3973\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_3_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9163\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK80_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDS_OUT_2_0_a2_0_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6878\,
            in2 => \_gnd_net_\,
            in3 => \N__3738\,
            lcout => \U712_REG_SM.LDS_OUT_2_0_a2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK40C_obuf_RNO_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4225\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDS_OUT_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000111110101"
        )
    port map (
            in0 => \N__3754\,
            in1 => \N__3681\,
            in2 => \N__4611\,
            in3 => \N__3582\,
            lcout => \U712_REG_SM.UDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9158\,
            ce => 'H',
            sr => \N__8944\
        );

    \U712_REG_SM.LDS_OUT_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101111"
        )
    port map (
            in0 => \N__3680\,
            in1 => \N__5919\,
            in2 => \N__3583\,
            in3 => \N__3753\,
            lcout => \U712_REG_SM.LDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9158\,
            ce => 'H',
            sr => \N__8944\
        );

    \U712_BUFFERS.un1_VBENn_0_a2_0_a2_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6826\,
            in2 => \_gnd_net_\,
            in3 => \N__7496\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_1_0_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6820\,
            in2 => \_gnd_net_\,
            in3 => \N__3694\,
            lcout => \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001000100"
        )
    port map (
            in0 => \N__3658\,
            in1 => \N__6821\,
            in2 => \_gnd_net_\,
            in3 => \N__3745\,
            lcout => \U712_BYTE_ENABLE.N_387\,
            ltout => \U712_BYTE_ENABLE.N_387_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_73_i_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__4192\,
            in1 => \N__4147\,
            in2 => \N__3718\,
            in3 => \N__3927\,
            lcout => \N_73_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_0_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__6822\,
            in1 => \N__3693\,
            in2 => \_gnd_net_\,
            in3 => \N__3654\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_srsts_0_i_o3_0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__5139\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3631\,
            lcout => \U712_REG_SM.N_301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010011000100"
        )
    port map (
            in0 => \N__3892\,
            in1 => \N__3882\,
            in2 => \N__3780\,
            in3 => \N__4020\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9155\,
            ce => 'H',
            sr => \N__8945\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000000000"
        )
    port map (
            in0 => \N__4021\,
            in1 => \N__3801\,
            in2 => \N__3781\,
            in3 => \N__4084\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9155\,
            ce => 'H',
            sr => \N__8945\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111000000000"
        )
    port map (
            in0 => \N__3819\,
            in1 => \N__4632\,
            in2 => \N__4072\,
            in3 => \N__4651\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9155\,
            ce => 'H',
            sr => \N__8945\
        );

    \U712_REG_SM.REG_CYCLE_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001110"
        )
    port map (
            in0 => \N__7486\,
            in1 => \N__3818\,
            in2 => \N__4678\,
            in3 => \N__4071\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9155\,
            ce => 'H',
            sr => \N__8945\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010111000001100"
        )
    port map (
            in0 => \N__3891\,
            in1 => \N__4309\,
            in2 => \N__4300\,
            in3 => \N__3883\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9155\,
            ce => 'H',
            sr => \N__8945\
        );

    \U712_REG_SM.REGENn_1_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000010111010"
        )
    port map (
            in0 => \N__4308\,
            in1 => \N__4273\,
            in2 => \N__3842\,
            in3 => \N__4299\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9155\,
            ce => 'H',
            sr => \N__8945\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101000100000"
        )
    port map (
            in0 => \N__4067\,
            in1 => \N__4083\,
            in2 => \N__3805\,
            in3 => \N__3820\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9155\,
            ce => 'H',
            sr => \N__8945\
        );

    \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__4339\,
            in1 => \N__3944\,
            in2 => \N__4006\,
            in3 => \N__4379\,
            lcout => \U712_REG_SM.N_281\,
            ltout => \U712_REG_SM.N_281_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_1_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__3800\,
            in1 => \N__4460\,
            in2 => \N__3787\,
            in3 => \N__4435\,
            lcout => \U712_REG_SM.N_369\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_0_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__6879\,
            in1 => \N__3945\,
            in2 => \_gnd_net_\,
            in3 => \N__4351\,
            lcout => \U712_REG_SM.N_123\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI90BP_0_2_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4459\,
            in2 => \_gnd_net_\,
            in3 => \N__4434\,
            lcout => \U712_REG_SM.N_280\,
            ltout => \U712_REG_SM.N_280_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNINB3L1_1_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__3772\,
            in1 => \N__4350\,
            in2 => \N__3784\,
            in3 => \N__4380\,
            lcout => \U712_REG_SM.N_424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3773\,
            in2 => \_gnd_net_\,
            in3 => \N__4019\,
            lcout => \U712_REG_SM.N_308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3943\,
            in2 => \_gnd_net_\,
            in3 => \N__4002\,
            lcout => \U712_REG_SM.N_288\,
            ltout => \U712_REG_SM.N_288_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4378\,
            in1 => \N__4340\,
            in2 => \N__4024\,
            in3 => \N__4043\,
            lcout => \U712_REG_SM.N_307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_2_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4384\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9159\,
            ce => 'H',
            sr => \N__8935\
        );

    \U712_REG_SM.C3_SYNC_0_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3991\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9159\,
            ce => 'H',
            sr => \N__8935\
        );

    \U712_REG_SM.C1_SYNC_0_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__3972\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9159\,
            ce => 'H',
            sr => \N__8935\
        );

    \U712_REG_SM.C1_SYNC_1_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4349\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9159\,
            ce => 'H',
            sr => \N__8935\
        );

    \U712_REG_SM.C3_SYNC_1_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3946\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9159\,
            ce => 'H',
            sr => \N__8935\
        );

    \U712_REG_SM.C3_SYNC_2_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4440\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9159\,
            ce => 'H',
            sr => \N__8935\
        );

    \U712_BYTE_ENABLE.N_75_i_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000101"
        )
    port map (
            in0 => \N__4161\,
            in1 => \N__4149\,
            in2 => \N__4093\,
            in3 => \N__3928\,
            lcout => \N_75_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7584\,
            in1 => \N__5247\,
            in2 => \_gnd_net_\,
            in3 => \N__6179\,
            lcout => \U712_BYTE_ENABLE.N_395\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_74_i_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__4148\,
            in1 => \N__4160\,
            in2 => \N__5275\,
            in3 => \N__4116\,
            lcout => \N_74_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_76_i_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__4162\,
            in1 => \N__4150\,
            in2 => \N__4120\,
            in3 => \N__5260\,
            lcout => \N_76_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__5246\,
            in1 => \N__7585\,
            in2 => \_gnd_net_\,
            in3 => \N__6180\,
            lcout => \U712_BYTE_ENABLE.N_391\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4056\,
            in1 => \N__4465\,
            in2 => \_gnd_net_\,
            in3 => \N__4441\,
            lcout => \U712_REG_SM.N_304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__4057\,
            in1 => \N__4045\,
            in2 => \N__5782\,
            in3 => \N__5755\,
            lcout => \U712_REG_SM.N_299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI0ULC2_4_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__4628\,
            in1 => \N__4055\,
            in2 => \_gnd_net_\,
            in3 => \N__4044\,
            lcout => \U712_REG_SM.N_298\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__4348\,
            in1 => \N__4383\,
            in2 => \N__4411\,
            in3 => \N__4295\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_373_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_6_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001110"
        )
    port map (
            in0 => \N__4396\,
            in1 => \N__4674\,
            in2 => \N__4027\,
            in3 => \N__4689\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9156\,
            ce => 'H',
            sr => \N__8936\
        );

    \U712_REG_SM.C1_SYNC_RNIIDN62_0_1_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4347\,
            in1 => \N__4382\,
            in2 => \N__4410\,
            in3 => \N__4293\,
            lcout => \U712_REG_SM.N_306\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4461\,
            in2 => \_gnd_net_\,
            in3 => \N__4436\,
            lcout => \U712_REG_SM.N_289\,
            ltout => \U712_REG_SM.N_289_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4395\,
            in1 => \N__4381\,
            in2 => \N__4354\,
            in3 => \N__4346\,
            lcout => \U712_REG_SM.N_494\,
            ltout => \U712_REG_SM.N_494_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_2_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010000"
        )
    port map (
            in0 => \N__4294\,
            in1 => \_gnd_net_\,
            in2 => \N__4276\,
            in3 => \N__4272\,
            lcout => OPEN,
            ltout => \U712_REG_SM.DS_EN_RNOZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__5939\,
            in1 => \N__4261\,
            in2 => \N__4255\,
            in3 => \N__4252\,
            lcout => \U712_REG_SM.DS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9156\,
            ce => 'H',
            sr => \N__8936\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110011110100"
        )
    port map (
            in0 => \N__4578\,
            in1 => \N__4236\,
            in2 => \N__4564\,
            in3 => \N__4219\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9157\,
            ce => 'H',
            sr => \N__8933\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100011111000"
        )
    port map (
            in0 => \N__4220\,
            in1 => \N__4579\,
            in2 => \N__5095\,
            in3 => \N__5071\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9157\,
            ce => 'H',
            sr => \N__8933\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__4577\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4221\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9157\,
            ce => 'H',
            sr => \N__8933\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4563\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9157\,
            ce => 'H',
            sr => \N__8933\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001000110000"
        )
    port map (
            in0 => \N__4534\,
            in1 => \N__4576\,
            in2 => \N__4825\,
            in3 => \N__5070\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9157\,
            ce => 'H',
            sr => \N__8933\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4546\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9157\,
            ce => 'H',
            sr => \N__8933\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4559\,
            in2 => \_gnd_net_\,
            in3 => \N__4545\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_obuft_RNO_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5044\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_886_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__4780\,
            in1 => \N__6809\,
            in2 => \N__8587\,
            in3 => \N__4942\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__6810\,
            in1 => \N__4507\,
            in2 => \N__4486\,
            in3 => \N__4483\,
            lcout => \U712_CHIP_RAM.N_313\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4716\,
            in2 => \_gnd_net_\,
            in3 => \N__4731\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4870\,
            in2 => \_gnd_net_\,
            in3 => \N__4471\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__4699\,
            ce => 'H',
            sr => \N__5983\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4897\,
            in2 => \_gnd_net_\,
            in3 => \N__4468\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__4699\,
            ce => 'H',
            sr => \N__5983\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4909\,
            in2 => \_gnd_net_\,
            in3 => \N__4741\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__4699\,
            ce => 'H',
            sr => \N__5983\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4846\,
            in2 => \_gnd_net_\,
            in3 => \N__4738\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__4699\,
            ce => 'H',
            sr => \N__5983\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4884\,
            in2 => \_gnd_net_\,
            in3 => \N__4735\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__4699\,
            ce => 'H',
            sr => \N__5983\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4732\,
            in2 => \_gnd_net_\,
            in3 => \N__4720\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__4699\,
            ce => 'H',
            sr => \N__5983\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4717\,
            in2 => \_gnd_net_\,
            in3 => \N__4705\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__4699\,
            ce => 'H',
            sr => \N__5983\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4858\,
            in2 => \_gnd_net_\,
            in3 => \N__4702\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4699\,
            ce => 'H',
            sr => \N__5983\
        );

    \U712_REG_SM.STATE_COUNT_5_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__4650\,
            in1 => \N__4673\,
            in2 => \_gnd_net_\,
            in3 => \N__4690\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9148\,
            ce => 'H',
            sr => \N__8937\
        );

    \U712_REG_SM.REG_TACK_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__4672\,
            in1 => \N__4649\,
            in2 => \N__4636\,
            in3 => \N__5107\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9148\,
            ce => 'H',
            sr => \N__8937\
        );

    \U712_REG_SM.UDS_OUT_RNIUP9B_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__5940\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4612\,
            lcout => \U712_REG_SM_un1_UDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__8235\,
            in1 => \N__5087\,
            in2 => \N__4824\,
            in3 => \N__5060\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_305_i_0_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9018\,
            in1 => \_gnd_net_\,
            in2 => \N__4807\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.N_305_i_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4804\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9117\,
            ce => \N__8636\,
            sr => \N__8965\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4803\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9118\,
            ce => \N__8727\,
            sr => \N__8956\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4774\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9118\,
            ce => \N__8727\,
            sr => \N__8956\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4972\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9118\,
            ce => \N__8727\,
            sr => \N__8956\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8692\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9118\,
            ce => \N__8727\,
            sr => \N__8956\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4936\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9118\,
            ce => \N__8727\,
            sr => \N__8956\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4770\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9122\,
            ce => \N__8635\,
            sr => \N__8951\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5584\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9122\,
            ce => \N__8635\,
            sr => \N__8951\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4971\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9122\,
            ce => \N__8635\,
            sr => \N__8951\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5623\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9122\,
            ce => \N__8635\,
            sr => \N__8951\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4935\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9126\,
            ce => \N__8641\,
            sr => \N__8943\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111101110"
        )
    port map (
            in0 => \N__8112\,
            in1 => \N__7991\,
            in2 => \N__7848\,
            in3 => \N__7731\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_341_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__7846\,
            in1 => \N__7765\,
            in2 => \N__4915\,
            in3 => \N__7382\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111001"
        )
    port map (
            in0 => \N__7383\,
            in1 => \N__7733\,
            in2 => \N__4912\,
            in3 => \N__7847\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__4908\,
            in1 => \N__4896\,
            in2 => \N__4885\,
            in3 => \N__4869\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111011111111"
        )
    port map (
            in0 => \N__4857\,
            in1 => \N__4845\,
            in2 => \N__4834\,
            in3 => \N__4831\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9130\,
            ce => 'H',
            sr => \N__8939\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010100000"
        )
    port map (
            in0 => \N__7381\,
            in1 => \_gnd_net_\,
            in2 => \N__7849\,
            in3 => \N__7732\,
            lcout => \U712_CHIP_RAM.N_403\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7582\,
            in1 => \N__5198\,
            in2 => \_gnd_net_\,
            in3 => \N__6177\,
            lcout => \U712_BYTE_ENABLE.N_392\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_0_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__6178\,
            in1 => \_gnd_net_\,
            in2 => \N__5203\,
            in3 => \N__7583\,
            lcout => \U712_BYTE_ENABLE.N_388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5248\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5202\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9135\,
            ce => 'H',
            sr => \N__8934\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011100000011"
        )
    port map (
            in0 => \N__6813\,
            in1 => \N__5176\,
            in2 => \N__5143\,
            in3 => \N__5794\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9135\,
            ce => 'H',
            sr => \N__8934\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5106\,
            in2 => \_gnd_net_\,
            in3 => \N__5955\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__8231\,
            in1 => \N__5094\,
            in2 => \_gnd_net_\,
            in3 => \N__5064\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9152\,
            ce => \N__5029\,
            sr => \N__8929\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8236\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_13_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__5014\,
            in1 => \N__5632\,
            in2 => \N__4993\,
            in3 => \N__6825\,
            lcout => \U712_CHIP_RAM.N_316\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101011011"
        )
    port map (
            in0 => \N__6776\,
            in1 => \N__5488\,
            in2 => \N__8588\,
            in3 => \N__5482\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__5476\,
            in1 => \N__5455\,
            in2 => \N__5431\,
            in3 => \N__6780\,
            lcout => \U712_CHIP_RAM.N_311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111110011"
        )
    port map (
            in0 => \N__5428\,
            in1 => \N__5419\,
            in2 => \N__6814\,
            in3 => \N__8575\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__5413\,
            in1 => \N__5395\,
            in2 => \N__5374\,
            in3 => \N__6781\,
            lcout => \U712_CHIP_RAM.N_312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__8576\,
            in1 => \N__7099\,
            in2 => \N__8442\,
            in3 => \N__8328\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9119\,
            ce => \N__6989\,
            sr => \N__8968\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__7094\,
            in1 => \N__5350\,
            in2 => \_gnd_net_\,
            in3 => \N__8431\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9123\,
            ce => \N__6971\,
            sr => \N__8966\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__5323\,
            in1 => \N__6815\,
            in2 => \N__8586\,
            in3 => \N__8653\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__6816\,
            in1 => \N__5317\,
            in2 => \N__5296\,
            in3 => \N__5293\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_314_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__8430\,
            in1 => \_gnd_net_\,
            in2 => \N__5662\,
            in3 => \N__7095\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9123\,
            ce => \N__6971\,
            sr => \N__8966\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111101"
        )
    port map (
            in0 => \N__5596\,
            in1 => \N__8537\,
            in2 => \N__6773\,
            in3 => \N__5638\,
            lcout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5622\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9127\,
            ce => \N__8726\,
            sr => \N__8957\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111101"
        )
    port map (
            in0 => \N__5551\,
            in1 => \N__8538\,
            in2 => \N__6774\,
            in3 => \N__5590\,
            lcout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5580\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9127\,
            ce => \N__8726\,
            sr => \N__8957\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111101"
        )
    port map (
            in0 => \N__5494\,
            in1 => \N__8539\,
            in2 => \N__6775\,
            in3 => \N__5542\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__6743\,
            in1 => \N__5536\,
            in2 => \N__5518\,
            in3 => \N__5515\,
            lcout => \U712_CHIP_RAM.N_317\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8800\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9127\,
            ce => \N__8726\,
            sr => \N__8957\
        );

    \U712_CHIP_RAM.DBDIR_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__6928\,
            in1 => \N__6413\,
            in2 => \_gnd_net_\,
            in3 => \N__6231\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9131\,
            ce => 'H',
            sr => \N__8952\
        );

    \U712_CHIP_RAM.DBR_SYNC_0_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5713\,
            lcout => \U712_REG_SM_DBR_SYNC_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9131\,
            ce => 'H',
            sr => \N__8952\
        );

    \U712_REG_SM.DBR_SYNC_1_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5775\,
            lcout => \U712_REG_SM_DBR_SYNC_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9131\,
            ce => 'H',
            sr => \N__8952\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011100000010"
        )
    port map (
            in0 => \N__6202\,
            in1 => \N__6629\,
            in2 => \N__7740\,
            in3 => \N__6747\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9131\,
            ce => 'H',
            sr => \N__8952\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNI32IV_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8230\,
            in2 => \_gnd_net_\,
            in3 => \N__6619\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIT6BC2_2_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__7370\,
            in1 => \N__7696\,
            in2 => \N__5692\,
            in3 => \N__8088\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIFP3R8_2_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__6245\,
            in1 => \N__6486\,
            in2 => \N__5689\,
            in3 => \N__6253\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111010"
        )
    port map (
            in0 => \N__5686\,
            in1 => \N__7572\,
            in2 => \N__6630\,
            in3 => \N__5677\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9139\,
            ce => 'H',
            sr => \N__8946\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__6246\,
            in1 => \N__6620\,
            in2 => \_gnd_net_\,
            in3 => \N__6487\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_0_i_0_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5676\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9139\,
            ce => 'H',
            sr => \N__8946\
        );

    \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__9020\,
            in1 => \N__5685\,
            in2 => \_gnd_net_\,
            in3 => \N__5675\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIKEL61_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__5793\,
            in1 => \N__5771\,
            in2 => \_gnd_net_\,
            in3 => \N__5748\,
            lcout => \U712_CHIP_RAM.N_285\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__8148\,
            in1 => \N__7373\,
            in2 => \_gnd_net_\,
            in3 => \N__6492\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000110010"
        )
    port map (
            in0 => \N__5737\,
            in1 => \N__6285\,
            in2 => \N__5731\,
            in3 => \N__8524\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9144\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_2_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__7976\,
            in1 => \N__8089\,
            in2 => \N__7827\,
            in3 => \N__7371\,
            lcout => \U712_CHIP_RAM.N_421\,
            ltout => \U712_CHIP_RAM.N_421_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIMMGI5_2_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__6124\,
            in1 => \_gnd_net_\,
            in2 => \N__5728\,
            in3 => \N__6510\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_293_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIJ42D8_0_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__7720\,
            in1 => \N__9019\,
            in2 => \N__5725\,
            in3 => \N__7245\,
            lcout => \U712_CHIP_RAM.N_309\,
            ltout => \U712_CHIP_RAM.N_309_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__7374\,
            in1 => \_gnd_net_\,
            in2 => \N__5722\,
            in3 => \N__7721\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9144\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__5719\,
            in1 => \N__8037\,
            in2 => \_gnd_net_\,
            in3 => \N__7244\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_RNO_1_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000100000000"
        )
    port map (
            in0 => \N__7372\,
            in1 => \N__7757\,
            in2 => \N__7735\,
            in3 => \N__7813\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0_a2_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__6100\,
            in1 => \N__5962\,
            in2 => \_gnd_net_\,
            in3 => \N__6547\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9149\,
            ce => 'H',
            sr => \N__8938\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110001000"
        )
    port map (
            in0 => \N__5956\,
            in1 => \N__6442\,
            in2 => \N__7407\,
            in3 => \N__6790\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9149\,
            ce => 'H',
            sr => \N__8938\
        );

    \U712_REG_SM.LDS_OUT_RNIL31J_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110111"
        )
    port map (
            in0 => \N__5944\,
            in1 => \N__5923\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM_un1_LDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__5887\,
            in1 => \N__7100\,
            in2 => \_gnd_net_\,
            in3 => \N__8435\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9120\,
            ce => \N__6978\,
            sr => \N__8980\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100011"
        )
    port map (
            in0 => \N__5863\,
            in1 => \N__8584\,
            in2 => \N__7108\,
            in3 => \N__8419\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9124\,
            ce => \N__6985\,
            sr => \N__8976\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100000001"
        )
    port map (
            in0 => \N__8583\,
            in1 => \N__7103\,
            in2 => \N__8436\,
            in3 => \N__5839\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9124\,
            ce => \N__6985\,
            sr => \N__8976\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI9T531_3_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__7077\,
            in1 => \N__8321\,
            in2 => \N__8585\,
            in3 => \N__5979\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_CMA31_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIV62J1_3_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9029\,
            in1 => \_gnd_net_\,
            in2 => \N__5812\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_CMA31_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__5809\,
            in1 => \N__6082\,
            in2 => \N__6076\,
            in3 => \N__6791\,
            lcout => \U712_CHIP_RAM.N_315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_2_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__6496\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7408\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_493_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_1_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__7246\,
            in1 => \N__7734\,
            in2 => \N__6055\,
            in3 => \N__8038\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9030\,
            in1 => \_gnd_net_\,
            in2 => \N__6052\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__6049\,
            in1 => \_gnd_net_\,
            in2 => \N__8426\,
            in3 => \N__7076\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9132\,
            ce => \N__6993\,
            sr => \N__8967\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101011111"
        )
    port map (
            in0 => \N__8398\,
            in1 => \_gnd_net_\,
            in2 => \N__8562\,
            in3 => \N__7075\,
            lcout => \U712_CHIP_RAM.CMA_5_i_0_8\,
            ltout => \U712_CHIP_RAM.CMA_5_i_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__8278\,
            in1 => \N__6028\,
            in2 => \N__6007\,
            in3 => \N__6748\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9132\,
            ce => \N__6993\,
            sr => \N__8967\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_RNITDMK_3_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__8397\,
            in1 => \N__8311\,
            in2 => \N__8561\,
            in3 => \N__7074\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_3_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__6130\,
            in1 => \N__7240\,
            in2 => \N__6232\,
            in3 => \N__7978\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9023\,
            in1 => \_gnd_net_\,
            in2 => \N__5965\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNI7Q5U5_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__6493\,
            in1 => \N__6247\,
            in2 => \N__6099\,
            in3 => \N__6624\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIAEJU_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__6625\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7722\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.DMA_CYCLE_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101111111001100"
        )
    port map (
            in0 => \N__6217\,
            in1 => \N__6151\,
            in2 => \N__6205\,
            in3 => \N__6201\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9140\,
            ce => 'H',
            sr => \N__8958\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNISB5T1_2_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__7699\,
            in1 => \N__7388\,
            in2 => \N__8115\,
            in3 => \N__6494\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_0_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_2_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__7977\,
            in1 => \N__7389\,
            in2 => \N__8116\,
            in3 => \N__6495\,
            lcout => \U712_CHIP_RAM.N_427\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI3F0BF_0_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001000"
        )
    port map (
            in0 => \N__6115\,
            in1 => \N__8122\,
            in2 => \N__6514\,
            in3 => \N__6109\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_sbtinv_3_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6103\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__7359\,
            in1 => \N__8016\,
            in2 => \N__7239\,
            in3 => \N__7694\,
            lcout => \U712_CHIP_RAM.N_296\,
            ltout => \U712_CHIP_RAM.N_296_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000010011"
        )
    port map (
            in0 => \N__7695\,
            in1 => \N__6298\,
            in2 => \N__6316\,
            in3 => \N__6313\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9145\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000001110"
        )
    port map (
            in0 => \N__6307\,
            in1 => \N__7441\,
            in2 => \N__6286\,
            in3 => \N__7073\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9145\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__7384\,
            in1 => \N__7726\,
            in2 => \N__8114\,
            in3 => \N__6296\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9145\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6297\,
            in1 => \N__7899\,
            in2 => \_gnd_net_\,
            in3 => \N__7990\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9145\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111100010"
        )
    port map (
            in0 => \N__7599\,
            in1 => \N__6284\,
            in2 => \N__8425\,
            in3 => \N__7423\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9145\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__6268\,
            in1 => \N__7579\,
            in2 => \_gnd_net_\,
            in3 => \N__6792\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9150\,
            ce => 'H',
            sr => \N__8947\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__7808\,
            in1 => \N__7238\,
            in2 => \_gnd_net_\,
            in3 => \N__6562\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9150\,
            ce => 'H',
            sr => \N__8947\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83_2_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110111"
        )
    port map (
            in0 => \N__7358\,
            in1 => \N__8087\,
            in2 => \N__7730\,
            in3 => \N__7221\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNISSMN4_3_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001010"
        )
    port map (
            in0 => \N__8225\,
            in1 => \N__7975\,
            in2 => \N__6256\,
            in3 => \N__6478\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__6545\,
            in1 => \N__6528\,
            in2 => \_gnd_net_\,
            in3 => \N__7807\,
            lcout => \U712_CHIP_RAM.N_282\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI7MV4_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6546\,
            in2 => \_gnd_net_\,
            in3 => \N__6529\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER46\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER46_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVE5T1_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__8017\,
            in1 => \N__7360\,
            in2 => \N__6517\,
            in3 => \N__7809\,
            lcout => \U712_CHIP_RAM.N_420\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110110111"
        )
    port map (
            in0 => \N__7361\,
            in1 => \N__8113\,
            in2 => \N__7741\,
            in3 => \N__6491\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_a5_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7992\,
            in2 => \N__6445\,
            in3 => \N__7236\,
            lcout => \U712_CHIP_RAM.N_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_i_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111010"
        )
    port map (
            in0 => \N__7581\,
            in1 => \N__6874\,
            in2 => \N__7513\,
            in3 => \N__6426\,
            lcout => \N_218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RASn_LC_15_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7107\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9121\,
            ce => 'H',
            sr => \N__8984\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__8737\,
            in1 => \N__6823\,
            in2 => \N__8595\,
            in3 => \N__8767\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_15_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__6824\,
            in1 => \N__6361\,
            in2 => \N__6340\,
            in3 => \N__6337\,
            lcout => \U712_CHIP_RAM.N_318\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__7183\,
            in1 => \N__7165\,
            in2 => \N__7453\,
            in3 => \N__6812\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9128\,
            ce => \N__6994\,
            sr => \N__8981\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__7135\,
            in1 => \_gnd_net_\,
            in2 => \N__8443\,
            in3 => \N__7102\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9128\,
            ce => \N__6994\,
            sr => \N__8981\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__8437\,
            in1 => \N__7101\,
            in2 => \_gnd_net_\,
            in3 => \N__7021\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9128\,
            ce => \N__6994\,
            sr => \N__8981\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000100"
        )
    port map (
            in0 => \N__6927\,
            in1 => \N__7545\,
            in2 => \N__6889\,
            in3 => \N__6811\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9133\,
            ce => \N__6643\,
            sr => \N__8977\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6634\,
            in2 => \_gnd_net_\,
            in3 => \N__7739\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9141\,
            ce => \N__6592\,
            sr => \N__8969\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_3_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__7600\,
            in1 => \N__7411\,
            in2 => \N__8152\,
            in3 => \N__7288\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9146\,
            ce => \N__6577\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__7410\,
            in1 => \N__8099\,
            in2 => \N__7993\,
            in3 => \N__6553\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_0_i_a2_1_0_a2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7409\,
            in1 => \N__7716\,
            in2 => \_gnd_net_\,
            in3 => \N__8098\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIO6AQ_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7700\,
            in2 => \_gnd_net_\,
            in3 => \N__7819\,
            lcout => \U712_CHIP_RAM.N_284\,
            ltout => \U712_CHIP_RAM.N_284_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101111"
        )
    port map (
            in0 => \N__8141\,
            in1 => \N__7413\,
            in2 => \N__7444\,
            in3 => \N__8036\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110000"
        )
    port map (
            in0 => \N__7412\,
            in1 => \N__7701\,
            in2 => \N__7839\,
            in3 => \N__7435\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__8226\,
            in1 => \N__8035\,
            in2 => \N__7426\,
            in3 => \N__7237\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__7898\,
            in1 => \N__7920\,
            in2 => \N__9031\,
            in3 => \N__7989\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9151\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7988\,
            in1 => \N__7869\,
            in2 => \N__7921\,
            in3 => \N__7897\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c6\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_12_c6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__9027\,
            in1 => \_gnd_net_\,
            in2 => \N__7417\,
            in3 => \N__7273\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9151\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_3_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100101010"
        )
    port map (
            in0 => \N__7702\,
            in1 => \N__7414\,
            in2 => \N__7838\,
            in3 => \N__8034\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__9022\,
            in1 => \N__7272\,
            in2 => \N__7282\,
            in3 => \N__7257\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9153\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__7271\,
            in1 => \N__7862\,
            in2 => \N__7258\,
            in3 => \N__7915\,
            lcout => \U712_CHIP_RAM.N_274\,
            ltout => \U712_CHIP_RAM.N_274_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__8224\,
            in1 => \_gnd_net_\,
            in2 => \N__8155\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_337\,
            ltout => \U712_CHIP_RAM.N_337_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITDHQ2_0_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8125\,
            in3 => \N__7697\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7973\,
            in2 => \_gnd_net_\,
            in3 => \N__8086\,
            lcout => \U712_CHIP_RAM.N_271\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_5_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__7974\,
            in1 => \N__7916\,
            in2 => \N__7873\,
            in3 => \N__7900\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__9021\,
            in1 => \_gnd_net_\,
            in2 => \N__7876\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9153\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVS9V_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100010"
        )
    port map (
            in0 => \N__7823\,
            in1 => \N__7761\,
            in2 => \_gnd_net_\,
            in3 => \N__7698\,
            lcout => \U712_CHIP_RAM.N_303\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_DRDENn_0_a2_0_a2_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7580\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7512\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8761\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9134\,
            ce => \N__8640\,
            sr => \N__8983\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_16_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8796\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9134\,
            ce => \N__8640\,
            sr => \N__8983\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8757\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9142\,
            ce => \N__8728\,
            sr => \N__8982\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8688\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9147\,
            ce => \N__8622\,
            sr => \N__8978\
        );

    \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__9028\,
            in1 => \N__9169\,
            in2 => \_gnd_net_\,
            in3 => \N__9180\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CASn_LC_17_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8596\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9125\,
            ce => 'H',
            sr => \N__8987\
        );

    \U712_CHIP_RAM.WEn_LC_17_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8441\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9129\,
            ce => 'H',
            sr => \N__8986\
        );

    \U712_CHIP_RAM.CRCSn_LC_17_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8329\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9143\,
            ce => 'H',
            sr => \N__8985\
        );

    \U712_CHIP_RAM.RAS_SYNC_0_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8277\,
            in2 => \_gnd_net_\,
            in3 => \N__8248\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9154\,
            ce => 'H',
            sr => \N__8979\
        );

    \U712_CHIP_RAM.RAS_SYNC_1_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9181\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9154\,
            ce => 'H',
            sr => \N__8979\
        );

    \CONSTANT_ONE_LUT4_LC_22_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

----------------------------------------------------------------------------------
--This work is shared under the Attribution-NonCommercial-ShareAlike 4.0 International (CC BY-NC-SA 4.0) License
--https://creativecommons.org/licenses/by-nc-sa/4.0/legalcode
	
--You are free to:
--Share - copy and redistribute the material in any medium or format
--Adapt - remix, transform, and build upon the material

--Under the following terms:

--Attribution - You must give appropriate credit, provide a link to the license, and indicate if changes were made. 
--You may do so in any reasonable manner, but not in any way that suggests the licensor endorses you or your use.

--NonCommercial - You may not use the material for commercial purposes.

--ShareAlike - If you remix, transform, or build upon the material, you must distribute your contributions under the 
--same license as the original.

--No additional restrictions - You may not apply legal terms or technological measures that legally restrict others 
--from doing anything the license permits.
--------------------------------------------------------------------------------------------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity IDE_CONTROLLER is

	Port ( 
	 
			BCLK : IN STD_LOGIC;
			A : in  STD_LOGIC_VECTOR (15 downto 10);
			nIDEEN : IN STD_LOGIC;
			nRESET : IN STD_LOGIC;
			nTIP : IN STD_LOGIC;
			RnW : IN STD_LOGIC;
			IORDY : IN STD_LOGIC;
			
			nCS0A : INOUT  STD_LOGIC;
			nCS1A : INOUT  STD_LOGIC;
			nCS0B : INOUT  STD_LOGIC;
			nCS1B : INOUT  STD_LOGIC;
			
			nDIOWA : OUT STD_LOGIC;
			nDIORA : OUT STD_LOGIC;
			nDIOWB : OUT STD_LOGIC;
			nDIORB : OUT STD_LOGIC;
			--AIDE : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
			nIDERESET : OUT STD_LOGIC;
			nTA : OUT STD_LOGIC;
			nTBI : OUT STD_LOGIC;
			nIDEROMEN : OUT STD_LOGIC
		
		);

end IDE_CONTROLLER;

architecture Behavioral of IDE_CONTROLLER is

	TYPE IDE_STATE IS ( IDLE, DIO, CYCLEACK, CYCLEEND );	
	SIGNAL CURRENT_STATE : IDE_STATE;

	SIGNAL IDECYCLE : STD_LOGIC;
	SIGNAL ENDCYCLE : STD_LOGIC;
	SIGNAL CYCLE16 : STD_LOGIC;
	SIGNAL READWRITECYCLE : STD_LOGIC;

	CONSTANT CLOCKPERIOD : INTEGER := 25; --THIS IS THE CLOCK PERIOD OF BCLK.
	CONSTANT PIO2T1 : INTEGER := (30 + (CLOCKPERIOD - 1)) / CLOCKPERIOD; --THIS FORMULA CAUSES THE QUOTIENT TO ROUND UP TO THE NEXT GREATER WHOLE INTEGER.
	CONSTANT PIO2T2_16 : INTEGER := (100 + (CLOCKPERIOD - 1)) / CLOCKPERIOD; --16 BIT T2 TIME
	CONSTANT PIO2T2_8 : INTEGER := (290 + (CLOCKPERIOD - 1)) / CLOCKPERIOD; --8 BIT T2 TIME
	CONSTANT PIO2T4 : INTEGER := (15 + (CLOCKPERIOD - 1)) / CLOCKPERIOD; 
	CONSTANT PIO2Teoc : INTEGER := (40 + (CLOCKPERIOD - 1)) / CLOCKPERIOD;
	
	CONSTANT T1 : INTEGER := PIO2T1;
	CONSTANT T2 : INTEGER := PIO2T1 + PIO2T2_16;
	CONSTANT T4 : INTEGER := PIO2T1 + PIO2T2_16 + PIO2T4;	
	CONSTANT Teoc : INTEGER := PIO2T1 + PIO2T2_16 + PIO2T4 + PIO2Teoc;
	CONSTANT DIFFERENTIAL : INTEGER := PIO2T2_8 - PIO2T2_16;

	SIGNAL COUNTER : INTEGER RANGE 0 TO Teoc + DIFFERENTIAL;
	

begin

	--IDE TIMINGS TAKEN FROM ATA/ATAPI-4 SPECIFICATIONS.
	--AT-APOLLO.DEVICE CHARACTERISTICS SUPPLIED BY FREDERIC REQUIN.
	
	--IN THIS LOGIC, THE "PRIMARY" PORT IS DEFINED WITH A TRAILING "A".
	--THE "SECONDARY" PORT IS DEFINED WITH A TRAILING "B".

	-----------
	-- RESET --
	-----------
	
	--PASS THE RESET SIGNAL ASYNCHRONOUSLY TO THE IDE PORTS.
	
	nIDERESET <= nRESET;
	
	---------------------
	-- IDE CHIP SELECT --
	---------------------
	
	--nCS0A AND nCS1A ARE CHIP SELECTS FOR THE "PRIMARY" PORT.
	--nCS0B AND nCS1B ARE CHIP SELECTS FOR THE "SECONDARY" PORT.
	--nIDEEN, WHEN ASSERTED, SIGNALS THAT WE ARE IN THE ADDRESS SPACE ASSIGNED TO THE IDE CONTROLLER.
	--nCS0A RESPONDS IN THE $0000 - $1FFC OFFSET WHILE nCS1A RESPONDS IN THE $2000-$3FFC OFFSET.
	--nCS0B RESPONDS IN THE $4000 - $5FFC OFFSET WHILE nCS1B RESPONDS IN THE $6000-$7FFC OFFSET.	
	--nIDEROMEN IS THE AUTO BOOT ROM AND RESPONDS AT OFFSET $8000.
	--THE IDE ADDRESS SIGNALS A2..A0 ARE CONNECTED TO THE MC68040 A12..A10.
	
	--$0000 = b0000000000000000
	--$1FFC = b0001111111111100
	
	--$2000 = b0010000000000000
	--$3FFC = b0011111111111100
	
	--$4000 = b0100000000000000
	--$5FFC = b0101111111111100
	
	--$6000 = b0110000000000000
	--$7FFC = b0111111111111100
	
	--$8000 = b1000000000000000
	
	--HERE, WE ARE PASSING THE DEVICE ADDRESS SIGNALS TO THE SELECTED IDE PORT WHEN WE ARE IN THE 
	--IDE ADDRESS SPACE, THE MC68040 IS IN A DATA TRANSFER CYCLE, AND WE ARE NOT IN RESET.
	
	nCS0A <= '0' WHEN A(15 DOWNTO 13) = "000" AND nIDEEN = '0' AND nTIP = '0' AND nRESET = '1' ELSE '1';
	nCS1A <= '0' WHEN A(15 DOWNTO 13) = "001" AND nIDEEN = '0' AND nTIP = '0' AND nRESET = '1' ELSE '1';
	nCS0B <= '0' WHEN A(15 DOWNTO 13) = "010" AND nIDEEN = '0' AND nTIP = '0' AND nRESET = '1' ELSE '1';
	nCS1B <= '0' WHEN A(15 DOWNTO 13) = "011" AND nIDEEN = '0' AND nTIP = '0' AND nRESET = '1' ELSE '1';
	nIDEROMEN <= '0' WHEN A(15 DOWNTO 13) = "100" AND nIDEEN = '0' AND nTIP = '0' AND nRESET = '1' ELSE '1';
	
	--AIDE <= A(12 DOWNTO 10);
	
	------------------
	-- IDE DATA I/O --
	------------------
	
	--ASSERT READ AND WRITE SIGNALS TO THE ACTIVE IDE PORT.
	
	nDIORA <= NOT (READWRITECYCLE AND RnW AND (NOT nCS0A OR NOT nCS1A)); 
	nDIOWA <= NOT (READWRITECYCLE AND NOT RnW AND (NOT nCS0A OR NOT nCS1A));
	
	nDIORB <= NOT (READWRITECYCLE AND RnW AND (NOT nCS0B OR NOT nCS1B));
	nDIOWB <= NOT (READWRITECYCLE AND NOT RnW AND (NOT nCS0B OR NOT nCS1B));	
	
	-----------------------------------
	-- IDE DATA TRANSFER ACKNOWLEDGE --
	-----------------------------------
	
	nTA <= 
			'Z' WHEN nIDEEN = '1' AND IDECYCLE = '0'
		ELSE
			'0' WHEN nIDEEN = '0' AND ENDCYCLE = '1'
		ELSE
			'1';
			
			
	nTBI <= 
			'Z' WHEN nIDEEN = '1' AND IDECYCLE = '0'
		ELSE
			'0' WHEN nIDEEN = '0' AND ENDCYCLE = '1'
		ELSE
			'1';
	
	------------------------------
	-- IDE DATA TRANSFER TIMING --
	------------------------------	
	
	--ACTIVITIES OF THE IDE DEVICE ARE ASYNCHRONOUS TO THE MC68040 BUS CLOCK.
	--TO IMPLEMENT THE CORRECT SETUP, HOLD, AND END OF CYCLE TIMING, WE 
	--COUNT THE NUMBER OF 40MHz BCLK TICKS TO DETERMINE WHEN WE CAN PROCEED
	--TO THE NEXT STEP.
	
	--WE WILL IMPLEMENT PIO2 TIMINGS. HERE ARE THE 16-BIT COMMAND TIMINGS:
	--T0 = 240ns = TOTAL CYCLE TIME
	--T1 = 30ns = SETUP TIME FOR DIOR/DIOW AFTER ASSERTION OF DEVICE ADDRESS SIGNALS.
	--T2 = 100ns = TIME FROM ASSERTION OF DIOR/DIOW THAT DATA BECOMES VALID (READ) OR LATCHED (WRITE)
	--T4 = 15ns = HOLD TIME NECESSARY AFTER NEGATION OF CHIP SELECT SIGNALS IN A WRITE CYCLE.
	--Teoc = 110ns = 240 - 30 - 100. THIS IS THE TIME BEFORE A NEW CYCLE MAY BE INITIATED.
	--THESE VALUES ARE DEFINED AS CONSTANTS AT THE START OF THIS FILE.
	
	--DATA TRANSFERS ARE 16 BITS. ALL OTHER COMMANDS ARE 8 BIT. THERE ARE DIFFERENT
	--TIMINGS BETWEEN THE 8 AND 16 BIT TRANSFERS. 16 BIT DATA TRANSFERS CAN BE 
	--IDENTIFIED BY CS0=0, CS1=1, DA2=0, DA1=0, DA0=0.			

	PROCESS (BCLK, nRESET) BEGIN
	
		IF nRESET = '0' THEN
		
			COUNTER <= 0;
			IDECYCLE <= '0';
			ENDCYCLE <= '0';
			CYCLE16 <= '0';
			READWRITECYCLE <= '0';
			CURRENT_STATE <= IDLE;
			
		ELSIF FALLING_EDGE (BCLK) THEN
			
			IF COUNTER /= 0 THEN COUNTER <= COUNTER + 1; END IF;
			
			CASE CURRENT_STATE IS
			
				WHEN IDLE =>
				
					IF nIDEEN = '0' AND nTIP = '0' AND COUNTER = 0 THEN --MC68040 TRANSFER HAS STARTED.
					
						COUNTER <= 1; 
						IDECYCLE <= '1';
						
					END IF;
					
					IF COUNTER = T1 THEN 
					
						CURRENT_STATE <= DIO;
						READWRITECYCLE <= '1'; --ASSERT DIOR/DIOW		
						CYCLE16 <= (NOT nCS0A OR NOT nCS0B) AND (nCS1A AND nCS1B) AND NOT A(12) AND NOT A(11) AND NOT A(10);
						
					END IF;
					
				WHEN DIO =>
				
					IF (CYCLE16 = '1' AND COUNTER = T2) OR (CYCLE16 = '0' AND COUNTER = T2 + DIFFERENTIAL) THEN					
						
						--THE DIOR/DIOW SETUP TIME HAS BEEN MET. END THE CYCLE.						
						ENDCYCLE <= '1'; --ASSERT TRANSFER ACK		
						READWRITECYCLE <= RnW; --NEGATE DIOW ON WRITE CYCLES
						CURRENT_STATE <= CYCLEACK;
						
					END IF;			
					
				WHEN CYCLEACK =>		

					--AT T4 WE REACH THE HOLD TIME REQUIRED FOR WRITE CYCLES.
					--WE ALSO APPLY IT TO READ CYCLES FOR SIMPLICITY. WE DO
					--NOT REALLY LOSE ANY TIME HERE BECAUSE OF THE CLOCK CYCLES
					--REQUIRED TO MEET ALL THE TIMINGS.
								
					ENDCYCLE <= '0'; --NEGATE TRANSFER ACK	
					READWRITECYCLE <= '0'; --NEGATE DIOR ON READ CYCLES
				
					IF CYCLE16 = '1' AND COUNTER = T4 THEN					
						
						IDECYCLE <= '0'; --TRISTATE TRANSFER ACK SIGNAL ONE CLOCK AFTER WE NEGATE TRANSFER ACK.
						CURRENT_STATE <= CYCLEEND;
						
					ELSIF CYCLE16 = '0' AND COUNTER >= T4 + DIFFERENTIAL THEN
					
						--DURING 8 BIT CYCLES, WE REACH THE MINIMUM CYCLE TIME HERE AND CAN SKIP THE TIME PADDING
						--REQUIRED BY THE 16 BIT CYCLE.
					
						IDECYCLE <= '0'; --TRISTATE TRANSFER ACK SIGNAL ONE CLOCK AFTER WE NEGATE TRANSFER ACK.
						COUNTER <= 0; --RESET THE IDE CLOCK COUNTER
						CURRENT_STATE <= IDLE;
					
					END IF;			
					
				WHEN CYCLEEND =>
				
					IF CYCLE16 = '1' AND COUNTER = Teoc THEN	
					
						COUNTER <= 0; --RESET THE IDE CLOCK COUNTER
						CURRENT_STATE <= IDLE;
					
					END IF;
					
				WHEN OTHERS =>
				
			END CASE;	
		
		END IF;
	
	END PROCESS;


end Behavioral;


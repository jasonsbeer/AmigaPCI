module U110_ARBITOR (

    output BGn

);

//GIVE THE CPU CONTINUOUS USE OF THE BUS FOR NOW.
assign BGn = 0;

endmodule

module U110_CYCLE_TERMINATION (

    output TEAn //,TACKn

);

//assign TACKn = 1'bz;
assign TEAn = 1;

endmodule

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Sep 14 2025 20:46:27

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    SIZ,
    DRA,
    CMA,
    DA,
    A,
    TBIn,
    RAMSPACEn,
    DBRn,
    RAMENn,
    TSn,
    LMBEn,
    DMA_LATCH_EN,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    UUBEn,
    LDSn,
    LATCH_CLK,
    CASUn,
    RAS1n,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    UMBEn,
    RAS0n,
    PRnW,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    BLSn,
    TCIn,
    WEn,
    REGENn,
    LLBEn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    input [1:0] SIZ;
    input [9:0] DRA;
    output [10:0] CMA;
    output [2:0] DA;
    input [20:0] A;
    output TBIn;
    input RAMSPACEn;
    input DBRn;
    output RAMENn;
    input TSn;
    output LMBEn;
    output DMA_LATCH_EN;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output UUBEn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    input RAS1n;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    output UMBEn;
    input RAS0n;
    output PRnW;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    output BLSn;
    output TCIn;
    output WEn;
    output REGENn;
    output LLBEn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__12997;
    wire N__12996;
    wire N__12995;
    wire N__12988;
    wire N__12987;
    wire N__12986;
    wire N__12979;
    wire N__12978;
    wire N__12977;
    wire N__12970;
    wire N__12969;
    wire N__12968;
    wire N__12961;
    wire N__12960;
    wire N__12959;
    wire N__12952;
    wire N__12951;
    wire N__12950;
    wire N__12943;
    wire N__12942;
    wire N__12941;
    wire N__12934;
    wire N__12933;
    wire N__12932;
    wire N__12925;
    wire N__12924;
    wire N__12923;
    wire N__12916;
    wire N__12915;
    wire N__12914;
    wire N__12907;
    wire N__12906;
    wire N__12905;
    wire N__12898;
    wire N__12897;
    wire N__12896;
    wire N__12889;
    wire N__12888;
    wire N__12887;
    wire N__12880;
    wire N__12879;
    wire N__12878;
    wire N__12871;
    wire N__12870;
    wire N__12869;
    wire N__12862;
    wire N__12861;
    wire N__12860;
    wire N__12853;
    wire N__12852;
    wire N__12851;
    wire N__12844;
    wire N__12843;
    wire N__12842;
    wire N__12835;
    wire N__12834;
    wire N__12833;
    wire N__12826;
    wire N__12825;
    wire N__12824;
    wire N__12817;
    wire N__12816;
    wire N__12815;
    wire N__12808;
    wire N__12807;
    wire N__12806;
    wire N__12799;
    wire N__12798;
    wire N__12797;
    wire N__12790;
    wire N__12789;
    wire N__12788;
    wire N__12781;
    wire N__12780;
    wire N__12779;
    wire N__12772;
    wire N__12771;
    wire N__12770;
    wire N__12763;
    wire N__12762;
    wire N__12761;
    wire N__12754;
    wire N__12753;
    wire N__12752;
    wire N__12745;
    wire N__12744;
    wire N__12743;
    wire N__12736;
    wire N__12735;
    wire N__12734;
    wire N__12727;
    wire N__12726;
    wire N__12725;
    wire N__12718;
    wire N__12717;
    wire N__12716;
    wire N__12709;
    wire N__12708;
    wire N__12707;
    wire N__12700;
    wire N__12699;
    wire N__12698;
    wire N__12691;
    wire N__12690;
    wire N__12689;
    wire N__12682;
    wire N__12681;
    wire N__12680;
    wire N__12673;
    wire N__12672;
    wire N__12671;
    wire N__12664;
    wire N__12663;
    wire N__12662;
    wire N__12655;
    wire N__12654;
    wire N__12653;
    wire N__12646;
    wire N__12645;
    wire N__12644;
    wire N__12637;
    wire N__12636;
    wire N__12635;
    wire N__12628;
    wire N__12627;
    wire N__12626;
    wire N__12619;
    wire N__12618;
    wire N__12617;
    wire N__12610;
    wire N__12609;
    wire N__12608;
    wire N__12601;
    wire N__12600;
    wire N__12599;
    wire N__12592;
    wire N__12591;
    wire N__12590;
    wire N__12583;
    wire N__12582;
    wire N__12581;
    wire N__12574;
    wire N__12573;
    wire N__12572;
    wire N__12565;
    wire N__12564;
    wire N__12563;
    wire N__12556;
    wire N__12555;
    wire N__12554;
    wire N__12547;
    wire N__12546;
    wire N__12545;
    wire N__12538;
    wire N__12537;
    wire N__12536;
    wire N__12529;
    wire N__12528;
    wire N__12527;
    wire N__12520;
    wire N__12519;
    wire N__12518;
    wire N__12511;
    wire N__12510;
    wire N__12509;
    wire N__12502;
    wire N__12501;
    wire N__12500;
    wire N__12493;
    wire N__12492;
    wire N__12491;
    wire N__12484;
    wire N__12483;
    wire N__12482;
    wire N__12475;
    wire N__12474;
    wire N__12473;
    wire N__12466;
    wire N__12465;
    wire N__12464;
    wire N__12457;
    wire N__12456;
    wire N__12455;
    wire N__12448;
    wire N__12447;
    wire N__12446;
    wire N__12439;
    wire N__12438;
    wire N__12437;
    wire N__12430;
    wire N__12429;
    wire N__12428;
    wire N__12421;
    wire N__12420;
    wire N__12419;
    wire N__12412;
    wire N__12411;
    wire N__12410;
    wire N__12403;
    wire N__12402;
    wire N__12401;
    wire N__12394;
    wire N__12393;
    wire N__12392;
    wire N__12385;
    wire N__12384;
    wire N__12383;
    wire N__12376;
    wire N__12375;
    wire N__12374;
    wire N__12367;
    wire N__12366;
    wire N__12365;
    wire N__12358;
    wire N__12357;
    wire N__12356;
    wire N__12349;
    wire N__12348;
    wire N__12347;
    wire N__12340;
    wire N__12339;
    wire N__12338;
    wire N__12331;
    wire N__12330;
    wire N__12329;
    wire N__12322;
    wire N__12321;
    wire N__12320;
    wire N__12313;
    wire N__12312;
    wire N__12311;
    wire N__12304;
    wire N__12303;
    wire N__12302;
    wire N__12295;
    wire N__12294;
    wire N__12293;
    wire N__12286;
    wire N__12285;
    wire N__12284;
    wire N__12277;
    wire N__12276;
    wire N__12275;
    wire N__12268;
    wire N__12267;
    wire N__12266;
    wire N__12259;
    wire N__12258;
    wire N__12257;
    wire N__12250;
    wire N__12249;
    wire N__12248;
    wire N__12241;
    wire N__12240;
    wire N__12239;
    wire N__12232;
    wire N__12231;
    wire N__12230;
    wire N__12223;
    wire N__12222;
    wire N__12221;
    wire N__12214;
    wire N__12213;
    wire N__12212;
    wire N__12205;
    wire N__12204;
    wire N__12203;
    wire N__12196;
    wire N__12195;
    wire N__12194;
    wire N__12187;
    wire N__12186;
    wire N__12185;
    wire N__12178;
    wire N__12177;
    wire N__12176;
    wire N__12169;
    wire N__12168;
    wire N__12167;
    wire N__12160;
    wire N__12159;
    wire N__12158;
    wire N__12151;
    wire N__12150;
    wire N__12149;
    wire N__12142;
    wire N__12141;
    wire N__12140;
    wire N__12133;
    wire N__12132;
    wire N__12131;
    wire N__12124;
    wire N__12123;
    wire N__12122;
    wire N__12105;
    wire N__12104;
    wire N__12103;
    wire N__12102;
    wire N__12099;
    wire N__12096;
    wire N__12091;
    wire N__12088;
    wire N__12083;
    wire N__12078;
    wire N__12075;
    wire N__12072;
    wire N__12069;
    wire N__12066;
    wire N__12063;
    wire N__12060;
    wire N__12057;
    wire N__12054;
    wire N__12051;
    wire N__12048;
    wire N__12045;
    wire N__12042;
    wire N__12039;
    wire N__12036;
    wire N__12035;
    wire N__12032;
    wire N__12029;
    wire N__12026;
    wire N__12023;
    wire N__12018;
    wire N__12015;
    wire N__12012;
    wire N__12009;
    wire N__12006;
    wire N__12005;
    wire N__12004;
    wire N__12003;
    wire N__12002;
    wire N__12001;
    wire N__12000;
    wire N__11999;
    wire N__11996;
    wire N__11995;
    wire N__11994;
    wire N__11993;
    wire N__11992;
    wire N__11991;
    wire N__11990;
    wire N__11989;
    wire N__11988;
    wire N__11987;
    wire N__11986;
    wire N__11977;
    wire N__11976;
    wire N__11975;
    wire N__11974;
    wire N__11973;
    wire N__11970;
    wire N__11965;
    wire N__11960;
    wire N__11953;
    wire N__11950;
    wire N__11943;
    wire N__11938;
    wire N__11935;
    wire N__11932;
    wire N__11931;
    wire N__11930;
    wire N__11927;
    wire N__11926;
    wire N__11925;
    wire N__11924;
    wire N__11923;
    wire N__11922;
    wire N__11921;
    wire N__11920;
    wire N__11919;
    wire N__11916;
    wire N__11913;
    wire N__11912;
    wire N__11911;
    wire N__11906;
    wire N__11903;
    wire N__11894;
    wire N__11889;
    wire N__11886;
    wire N__11883;
    wire N__11880;
    wire N__11873;
    wire N__11870;
    wire N__11865;
    wire N__11862;
    wire N__11853;
    wire N__11850;
    wire N__11847;
    wire N__11846;
    wire N__11835;
    wire N__11834;
    wire N__11833;
    wire N__11832;
    wire N__11829;
    wire N__11820;
    wire N__11815;
    wire N__11812;
    wire N__11809;
    wire N__11806;
    wire N__11803;
    wire N__11798;
    wire N__11795;
    wire N__11792;
    wire N__11789;
    wire N__11784;
    wire N__11781;
    wire N__11776;
    wire N__11771;
    wire N__11768;
    wire N__11761;
    wire N__11754;
    wire N__11751;
    wire N__11748;
    wire N__11745;
    wire N__11742;
    wire N__11739;
    wire N__11738;
    wire N__11737;
    wire N__11736;
    wire N__11735;
    wire N__11734;
    wire N__11733;
    wire N__11732;
    wire N__11731;
    wire N__11730;
    wire N__11729;
    wire N__11728;
    wire N__11727;
    wire N__11726;
    wire N__11725;
    wire N__11724;
    wire N__11723;
    wire N__11722;
    wire N__11721;
    wire N__11720;
    wire N__11719;
    wire N__11718;
    wire N__11717;
    wire N__11716;
    wire N__11715;
    wire N__11714;
    wire N__11713;
    wire N__11712;
    wire N__11711;
    wire N__11710;
    wire N__11709;
    wire N__11708;
    wire N__11707;
    wire N__11706;
    wire N__11705;
    wire N__11704;
    wire N__11703;
    wire N__11702;
    wire N__11701;
    wire N__11700;
    wire N__11699;
    wire N__11698;
    wire N__11697;
    wire N__11696;
    wire N__11695;
    wire N__11694;
    wire N__11693;
    wire N__11690;
    wire N__11689;
    wire N__11592;
    wire N__11589;
    wire N__11586;
    wire N__11585;
    wire N__11584;
    wire N__11583;
    wire N__11580;
    wire N__11577;
    wire N__11572;
    wire N__11569;
    wire N__11564;
    wire N__11561;
    wire N__11558;
    wire N__11555;
    wire N__11550;
    wire N__11547;
    wire N__11544;
    wire N__11543;
    wire N__11542;
    wire N__11541;
    wire N__11538;
    wire N__11535;
    wire N__11530;
    wire N__11527;
    wire N__11522;
    wire N__11519;
    wire N__11516;
    wire N__11513;
    wire N__11508;
    wire N__11505;
    wire N__11502;
    wire N__11499;
    wire N__11496;
    wire N__11495;
    wire N__11494;
    wire N__11493;
    wire N__11490;
    wire N__11487;
    wire N__11484;
    wire N__11481;
    wire N__11474;
    wire N__11471;
    wire N__11468;
    wire N__11465;
    wire N__11462;
    wire N__11459;
    wire N__11456;
    wire N__11453;
    wire N__11448;
    wire N__11447;
    wire N__11444;
    wire N__11441;
    wire N__11440;
    wire N__11439;
    wire N__11434;
    wire N__11431;
    wire N__11428;
    wire N__11423;
    wire N__11420;
    wire N__11417;
    wire N__11414;
    wire N__11411;
    wire N__11408;
    wire N__11405;
    wire N__11400;
    wire N__11397;
    wire N__11396;
    wire N__11395;
    wire N__11394;
    wire N__11393;
    wire N__11390;
    wire N__11387;
    wire N__11386;
    wire N__11385;
    wire N__11384;
    wire N__11383;
    wire N__11380;
    wire N__11379;
    wire N__11378;
    wire N__11377;
    wire N__11376;
    wire N__11375;
    wire N__11370;
    wire N__11367;
    wire N__11360;
    wire N__11357;
    wire N__11356;
    wire N__11353;
    wire N__11352;
    wire N__11351;
    wire N__11350;
    wire N__11347;
    wire N__11344;
    wire N__11339;
    wire N__11334;
    wire N__11331;
    wire N__11326;
    wire N__11317;
    wire N__11314;
    wire N__11311;
    wire N__11308;
    wire N__11305;
    wire N__11304;
    wire N__11299;
    wire N__11298;
    wire N__11297;
    wire N__11286;
    wire N__11281;
    wire N__11278;
    wire N__11275;
    wire N__11272;
    wire N__11269;
    wire N__11266;
    wire N__11263;
    wire N__11254;
    wire N__11251;
    wire N__11248;
    wire N__11243;
    wire N__11240;
    wire N__11237;
    wire N__11232;
    wire N__11231;
    wire N__11228;
    wire N__11225;
    wire N__11222;
    wire N__11219;
    wire N__11216;
    wire N__11213;
    wire N__11208;
    wire N__11207;
    wire N__11206;
    wire N__11205;
    wire N__11204;
    wire N__11203;
    wire N__11190;
    wire N__11187;
    wire N__11184;
    wire N__11183;
    wire N__11182;
    wire N__11181;
    wire N__11180;
    wire N__11179;
    wire N__11178;
    wire N__11177;
    wire N__11176;
    wire N__11175;
    wire N__11174;
    wire N__11151;
    wire N__11148;
    wire N__11145;
    wire N__11144;
    wire N__11143;
    wire N__11142;
    wire N__11141;
    wire N__11140;
    wire N__11139;
    wire N__11136;
    wire N__11131;
    wire N__11128;
    wire N__11125;
    wire N__11122;
    wire N__11119;
    wire N__11118;
    wire N__11117;
    wire N__11116;
    wire N__11115;
    wire N__11114;
    wire N__11113;
    wire N__11112;
    wire N__11111;
    wire N__11110;
    wire N__11109;
    wire N__11108;
    wire N__11107;
    wire N__11106;
    wire N__11105;
    wire N__11104;
    wire N__11103;
    wire N__11102;
    wire N__11099;
    wire N__11098;
    wire N__11097;
    wire N__11096;
    wire N__11093;
    wire N__11092;
    wire N__11089;
    wire N__11086;
    wire N__11085;
    wire N__11084;
    wire N__11083;
    wire N__11082;
    wire N__11081;
    wire N__11080;
    wire N__11079;
    wire N__11078;
    wire N__11077;
    wire N__11076;
    wire N__11075;
    wire N__11074;
    wire N__11073;
    wire N__11070;
    wire N__11069;
    wire N__11068;
    wire N__11067;
    wire N__11064;
    wire N__11063;
    wire N__11062;
    wire N__10971;
    wire N__10968;
    wire N__10965;
    wire N__10964;
    wire N__10963;
    wire N__10960;
    wire N__10959;
    wire N__10956;
    wire N__10955;
    wire N__10952;
    wire N__10949;
    wire N__10946;
    wire N__10943;
    wire N__10940;
    wire N__10935;
    wire N__10932;
    wire N__10929;
    wire N__10926;
    wire N__10923;
    wire N__10920;
    wire N__10917;
    wire N__10914;
    wire N__10909;
    wire N__10904;
    wire N__10901;
    wire N__10896;
    wire N__10893;
    wire N__10890;
    wire N__10889;
    wire N__10886;
    wire N__10883;
    wire N__10882;
    wire N__10881;
    wire N__10878;
    wire N__10875;
    wire N__10870;
    wire N__10869;
    wire N__10864;
    wire N__10861;
    wire N__10858;
    wire N__10857;
    wire N__10852;
    wire N__10849;
    wire N__10846;
    wire N__10843;
    wire N__10840;
    wire N__10837;
    wire N__10834;
    wire N__10831;
    wire N__10828;
    wire N__10821;
    wire N__10818;
    wire N__10815;
    wire N__10814;
    wire N__10811;
    wire N__10808;
    wire N__10807;
    wire N__10804;
    wire N__10801;
    wire N__10798;
    wire N__10795;
    wire N__10792;
    wire N__10789;
    wire N__10782;
    wire N__10779;
    wire N__10778;
    wire N__10777;
    wire N__10772;
    wire N__10771;
    wire N__10770;
    wire N__10767;
    wire N__10764;
    wire N__10759;
    wire N__10756;
    wire N__10753;
    wire N__10750;
    wire N__10747;
    wire N__10746;
    wire N__10743;
    wire N__10740;
    wire N__10737;
    wire N__10734;
    wire N__10731;
    wire N__10728;
    wire N__10725;
    wire N__10722;
    wire N__10717;
    wire N__10712;
    wire N__10707;
    wire N__10704;
    wire N__10701;
    wire N__10698;
    wire N__10695;
    wire N__10692;
    wire N__10689;
    wire N__10686;
    wire N__10683;
    wire N__10680;
    wire N__10677;
    wire N__10674;
    wire N__10671;
    wire N__10668;
    wire N__10665;
    wire N__10662;
    wire N__10659;
    wire N__10658;
    wire N__10655;
    wire N__10654;
    wire N__10653;
    wire N__10650;
    wire N__10647;
    wire N__10644;
    wire N__10641;
    wire N__10638;
    wire N__10631;
    wire N__10628;
    wire N__10625;
    wire N__10622;
    wire N__10619;
    wire N__10614;
    wire N__10611;
    wire N__10608;
    wire N__10605;
    wire N__10602;
    wire N__10601;
    wire N__10600;
    wire N__10599;
    wire N__10596;
    wire N__10591;
    wire N__10590;
    wire N__10587;
    wire N__10582;
    wire N__10579;
    wire N__10572;
    wire N__10569;
    wire N__10566;
    wire N__10563;
    wire N__10560;
    wire N__10557;
    wire N__10554;
    wire N__10551;
    wire N__10548;
    wire N__10545;
    wire N__10542;
    wire N__10539;
    wire N__10536;
    wire N__10533;
    wire N__10530;
    wire N__10529;
    wire N__10528;
    wire N__10525;
    wire N__10522;
    wire N__10519;
    wire N__10518;
    wire N__10517;
    wire N__10516;
    wire N__10515;
    wire N__10514;
    wire N__10511;
    wire N__10510;
    wire N__10507;
    wire N__10504;
    wire N__10501;
    wire N__10500;
    wire N__10499;
    wire N__10498;
    wire N__10495;
    wire N__10494;
    wire N__10489;
    wire N__10486;
    wire N__10485;
    wire N__10484;
    wire N__10483;
    wire N__10480;
    wire N__10477;
    wire N__10476;
    wire N__10475;
    wire N__10474;
    wire N__10469;
    wire N__10468;
    wire N__10467;
    wire N__10466;
    wire N__10463;
    wire N__10460;
    wire N__10457;
    wire N__10454;
    wire N__10449;
    wire N__10448;
    wire N__10445;
    wire N__10442;
    wire N__10439;
    wire N__10436;
    wire N__10435;
    wire N__10432;
    wire N__10429;
    wire N__10426;
    wire N__10423;
    wire N__10418;
    wire N__10415;
    wire N__10412;
    wire N__10407;
    wire N__10402;
    wire N__10399;
    wire N__10396;
    wire N__10393;
    wire N__10390;
    wire N__10389;
    wire N__10384;
    wire N__10381;
    wire N__10378;
    wire N__10375;
    wire N__10368;
    wire N__10359;
    wire N__10354;
    wire N__10345;
    wire N__10342;
    wire N__10323;
    wire N__10320;
    wire N__10317;
    wire N__10314;
    wire N__10311;
    wire N__10308;
    wire N__10305;
    wire N__10302;
    wire N__10301;
    wire N__10298;
    wire N__10295;
    wire N__10294;
    wire N__10293;
    wire N__10292;
    wire N__10291;
    wire N__10290;
    wire N__10289;
    wire N__10286;
    wire N__10283;
    wire N__10276;
    wire N__10273;
    wire N__10270;
    wire N__10267;
    wire N__10266;
    wire N__10265;
    wire N__10260;
    wire N__10257;
    wire N__10254;
    wire N__10249;
    wire N__10246;
    wire N__10243;
    wire N__10230;
    wire N__10229;
    wire N__10228;
    wire N__10227;
    wire N__10224;
    wire N__10221;
    wire N__10218;
    wire N__10215;
    wire N__10212;
    wire N__10209;
    wire N__10208;
    wire N__10207;
    wire N__10204;
    wire N__10201;
    wire N__10198;
    wire N__10195;
    wire N__10194;
    wire N__10191;
    wire N__10188;
    wire N__10185;
    wire N__10182;
    wire N__10179;
    wire N__10176;
    wire N__10173;
    wire N__10168;
    wire N__10165;
    wire N__10162;
    wire N__10157;
    wire N__10146;
    wire N__10143;
    wire N__10140;
    wire N__10137;
    wire N__10134;
    wire N__10131;
    wire N__10128;
    wire N__10125;
    wire N__10122;
    wire N__10119;
    wire N__10116;
    wire N__10113;
    wire N__10112;
    wire N__10109;
    wire N__10108;
    wire N__10105;
    wire N__10102;
    wire N__10099;
    wire N__10098;
    wire N__10097;
    wire N__10096;
    wire N__10093;
    wire N__10088;
    wire N__10085;
    wire N__10084;
    wire N__10081;
    wire N__10080;
    wire N__10077;
    wire N__10070;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10053;
    wire N__10050;
    wire N__10047;
    wire N__10042;
    wire N__10035;
    wire N__10034;
    wire N__10031;
    wire N__10030;
    wire N__10027;
    wire N__10026;
    wire N__10023;
    wire N__10020;
    wire N__10017;
    wire N__10014;
    wire N__10011;
    wire N__10004;
    wire N__10001;
    wire N__9998;
    wire N__9993;
    wire N__9990;
    wire N__9987;
    wire N__9984;
    wire N__9981;
    wire N__9978;
    wire N__9975;
    wire N__9972;
    wire N__9971;
    wire N__9970;
    wire N__9969;
    wire N__9966;
    wire N__9963;
    wire N__9960;
    wire N__9959;
    wire N__9956;
    wire N__9951;
    wire N__9948;
    wire N__9945;
    wire N__9942;
    wire N__9939;
    wire N__9936;
    wire N__9933;
    wire N__9924;
    wire N__9921;
    wire N__9918;
    wire N__9915;
    wire N__9912;
    wire N__9909;
    wire N__9906;
    wire N__9905;
    wire N__9902;
    wire N__9899;
    wire N__9898;
    wire N__9897;
    wire N__9894;
    wire N__9893;
    wire N__9890;
    wire N__9887;
    wire N__9884;
    wire N__9881;
    wire N__9880;
    wire N__9877;
    wire N__9870;
    wire N__9867;
    wire N__9864;
    wire N__9855;
    wire N__9852;
    wire N__9851;
    wire N__9850;
    wire N__9849;
    wire N__9848;
    wire N__9847;
    wire N__9846;
    wire N__9845;
    wire N__9844;
    wire N__9841;
    wire N__9838;
    wire N__9837;
    wire N__9836;
    wire N__9835;
    wire N__9832;
    wire N__9829;
    wire N__9826;
    wire N__9825;
    wire N__9824;
    wire N__9823;
    wire N__9822;
    wire N__9821;
    wire N__9820;
    wire N__9817;
    wire N__9814;
    wire N__9809;
    wire N__9808;
    wire N__9805;
    wire N__9802;
    wire N__9799;
    wire N__9794;
    wire N__9789;
    wire N__9784;
    wire N__9777;
    wire N__9774;
    wire N__9771;
    wire N__9770;
    wire N__9769;
    wire N__9768;
    wire N__9761;
    wire N__9758;
    wire N__9755;
    wire N__9752;
    wire N__9749;
    wire N__9746;
    wire N__9739;
    wire N__9738;
    wire N__9737;
    wire N__9736;
    wire N__9731;
    wire N__9730;
    wire N__9723;
    wire N__9720;
    wire N__9707;
    wire N__9700;
    wire N__9697;
    wire N__9694;
    wire N__9681;
    wire N__9678;
    wire N__9675;
    wire N__9672;
    wire N__9669;
    wire N__9666;
    wire N__9663;
    wire N__9660;
    wire N__9657;
    wire N__9654;
    wire N__9651;
    wire N__9648;
    wire N__9645;
    wire N__9642;
    wire N__9639;
    wire N__9636;
    wire N__9633;
    wire N__9630;
    wire N__9627;
    wire N__9624;
    wire N__9621;
    wire N__9618;
    wire N__9615;
    wire N__9612;
    wire N__9609;
    wire N__9606;
    wire N__9603;
    wire N__9600;
    wire N__9597;
    wire N__9594;
    wire N__9591;
    wire N__9588;
    wire N__9585;
    wire N__9582;
    wire N__9579;
    wire N__9576;
    wire N__9573;
    wire N__9570;
    wire N__9567;
    wire N__9564;
    wire N__9561;
    wire N__9558;
    wire N__9557;
    wire N__9552;
    wire N__9549;
    wire N__9548;
    wire N__9547;
    wire N__9544;
    wire N__9539;
    wire N__9534;
    wire N__9531;
    wire N__9528;
    wire N__9527;
    wire N__9526;
    wire N__9523;
    wire N__9520;
    wire N__9517;
    wire N__9516;
    wire N__9509;
    wire N__9506;
    wire N__9503;
    wire N__9500;
    wire N__9497;
    wire N__9494;
    wire N__9489;
    wire N__9486;
    wire N__9483;
    wire N__9480;
    wire N__9477;
    wire N__9474;
    wire N__9473;
    wire N__9470;
    wire N__9467;
    wire N__9464;
    wire N__9461;
    wire N__9456;
    wire N__9453;
    wire N__9450;
    wire N__9447;
    wire N__9444;
    wire N__9441;
    wire N__9438;
    wire N__9435;
    wire N__9432;
    wire N__9429;
    wire N__9426;
    wire N__9423;
    wire N__9420;
    wire N__9417;
    wire N__9414;
    wire N__9411;
    wire N__9408;
    wire N__9405;
    wire N__9402;
    wire N__9399;
    wire N__9396;
    wire N__9393;
    wire N__9390;
    wire N__9387;
    wire N__9384;
    wire N__9381;
    wire N__9380;
    wire N__9379;
    wire N__9376;
    wire N__9373;
    wire N__9370;
    wire N__9367;
    wire N__9364;
    wire N__9361;
    wire N__9360;
    wire N__9357;
    wire N__9354;
    wire N__9351;
    wire N__9348;
    wire N__9343;
    wire N__9336;
    wire N__9333;
    wire N__9330;
    wire N__9327;
    wire N__9324;
    wire N__9321;
    wire N__9318;
    wire N__9315;
    wire N__9312;
    wire N__9309;
    wire N__9306;
    wire N__9303;
    wire N__9300;
    wire N__9297;
    wire N__9294;
    wire N__9291;
    wire N__9288;
    wire N__9285;
    wire N__9282;
    wire N__9279;
    wire N__9276;
    wire N__9273;
    wire N__9270;
    wire N__9267;
    wire N__9264;
    wire N__9261;
    wire N__9258;
    wire N__9255;
    wire N__9252;
    wire N__9249;
    wire N__9246;
    wire N__9243;
    wire N__9240;
    wire N__9237;
    wire N__9234;
    wire N__9231;
    wire N__9228;
    wire N__9225;
    wire N__9222;
    wire N__9219;
    wire N__9216;
    wire N__9213;
    wire N__9210;
    wire N__9207;
    wire N__9204;
    wire N__9201;
    wire N__9198;
    wire N__9195;
    wire N__9192;
    wire N__9189;
    wire N__9188;
    wire N__9185;
    wire N__9182;
    wire N__9181;
    wire N__9178;
    wire N__9175;
    wire N__9172;
    wire N__9169;
    wire N__9166;
    wire N__9163;
    wire N__9156;
    wire N__9153;
    wire N__9150;
    wire N__9149;
    wire N__9146;
    wire N__9143;
    wire N__9140;
    wire N__9135;
    wire N__9132;
    wire N__9129;
    wire N__9126;
    wire N__9123;
    wire N__9120;
    wire N__9117;
    wire N__9114;
    wire N__9111;
    wire N__9108;
    wire N__9105;
    wire N__9102;
    wire N__9101;
    wire N__9100;
    wire N__9097;
    wire N__9096;
    wire N__9093;
    wire N__9092;
    wire N__9089;
    wire N__9088;
    wire N__9087;
    wire N__9086;
    wire N__9085;
    wire N__9082;
    wire N__9079;
    wire N__9076;
    wire N__9071;
    wire N__9068;
    wire N__9063;
    wire N__9060;
    wire N__9045;
    wire N__9044;
    wire N__9043;
    wire N__9042;
    wire N__9037;
    wire N__9032;
    wire N__9027;
    wire N__9026;
    wire N__9025;
    wire N__9022;
    wire N__9019;
    wire N__9018;
    wire N__9017;
    wire N__9016;
    wire N__9015;
    wire N__9012;
    wire N__9011;
    wire N__9010;
    wire N__9007;
    wire N__9004;
    wire N__9001;
    wire N__8998;
    wire N__8991;
    wire N__8986;
    wire N__8979;
    wire N__8970;
    wire N__8969;
    wire N__8966;
    wire N__8965;
    wire N__8962;
    wire N__8961;
    wire N__8960;
    wire N__8959;
    wire N__8958;
    wire N__8957;
    wire N__8956;
    wire N__8953;
    wire N__8950;
    wire N__8947;
    wire N__8944;
    wire N__8939;
    wire N__8932;
    wire N__8919;
    wire N__8916;
    wire N__8913;
    wire N__8910;
    wire N__8907;
    wire N__8904;
    wire N__8901;
    wire N__8898;
    wire N__8895;
    wire N__8892;
    wire N__8889;
    wire N__8886;
    wire N__8883;
    wire N__8880;
    wire N__8877;
    wire N__8874;
    wire N__8871;
    wire N__8868;
    wire N__8865;
    wire N__8862;
    wire N__8859;
    wire N__8856;
    wire N__8853;
    wire N__8850;
    wire N__8847;
    wire N__8844;
    wire N__8841;
    wire N__8838;
    wire N__8835;
    wire N__8832;
    wire N__8829;
    wire N__8826;
    wire N__8825;
    wire N__8824;
    wire N__8821;
    wire N__8818;
    wire N__8815;
    wire N__8812;
    wire N__8809;
    wire N__8806;
    wire N__8799;
    wire N__8796;
    wire N__8793;
    wire N__8792;
    wire N__8789;
    wire N__8786;
    wire N__8783;
    wire N__8778;
    wire N__8775;
    wire N__8774;
    wire N__8771;
    wire N__8768;
    wire N__8765;
    wire N__8760;
    wire N__8757;
    wire N__8756;
    wire N__8755;
    wire N__8754;
    wire N__8751;
    wire N__8746;
    wire N__8745;
    wire N__8744;
    wire N__8743;
    wire N__8742;
    wire N__8739;
    wire N__8736;
    wire N__8733;
    wire N__8724;
    wire N__8721;
    wire N__8718;
    wire N__8709;
    wire N__8706;
    wire N__8705;
    wire N__8702;
    wire N__8699;
    wire N__8694;
    wire N__8693;
    wire N__8692;
    wire N__8691;
    wire N__8690;
    wire N__8689;
    wire N__8688;
    wire N__8685;
    wire N__8678;
    wire N__8671;
    wire N__8668;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8652;
    wire N__8651;
    wire N__8648;
    wire N__8647;
    wire N__8646;
    wire N__8643;
    wire N__8640;
    wire N__8637;
    wire N__8634;
    wire N__8633;
    wire N__8628;
    wire N__8627;
    wire N__8626;
    wire N__8625;
    wire N__8624;
    wire N__8623;
    wire N__8622;
    wire N__8617;
    wire N__8616;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8596;
    wire N__8593;
    wire N__8590;
    wire N__8585;
    wire N__8568;
    wire N__8565;
    wire N__8562;
    wire N__8559;
    wire N__8556;
    wire N__8553;
    wire N__8550;
    wire N__8549;
    wire N__8548;
    wire N__8547;
    wire N__8542;
    wire N__8541;
    wire N__8538;
    wire N__8535;
    wire N__8532;
    wire N__8529;
    wire N__8526;
    wire N__8523;
    wire N__8522;
    wire N__8521;
    wire N__8516;
    wire N__8511;
    wire N__8508;
    wire N__8505;
    wire N__8502;
    wire N__8499;
    wire N__8494;
    wire N__8487;
    wire N__8486;
    wire N__8485;
    wire N__8484;
    wire N__8477;
    wire N__8474;
    wire N__8469;
    wire N__8468;
    wire N__8467;
    wire N__8464;
    wire N__8461;
    wire N__8458;
    wire N__8453;
    wire N__8450;
    wire N__8447;
    wire N__8442;
    wire N__8441;
    wire N__8440;
    wire N__8439;
    wire N__8438;
    wire N__8437;
    wire N__8436;
    wire N__8435;
    wire N__8434;
    wire N__8431;
    wire N__8430;
    wire N__8427;
    wire N__8426;
    wire N__8425;
    wire N__8424;
    wire N__8423;
    wire N__8418;
    wire N__8417;
    wire N__8410;
    wire N__8409;
    wire N__8406;
    wire N__8405;
    wire N__8404;
    wire N__8403;
    wire N__8402;
    wire N__8401;
    wire N__8400;
    wire N__8397;
    wire N__8394;
    wire N__8391;
    wire N__8388;
    wire N__8385;
    wire N__8384;
    wire N__8379;
    wire N__8376;
    wire N__8373;
    wire N__8372;
    wire N__8371;
    wire N__8368;
    wire N__8365;
    wire N__8358;
    wire N__8351;
    wire N__8348;
    wire N__8347;
    wire N__8346;
    wire N__8343;
    wire N__8340;
    wire N__8333;
    wire N__8328;
    wire N__8321;
    wire N__8314;
    wire N__8307;
    wire N__8300;
    wire N__8297;
    wire N__8280;
    wire N__8277;
    wire N__8274;
    wire N__8271;
    wire N__8268;
    wire N__8265;
    wire N__8264;
    wire N__8261;
    wire N__8258;
    wire N__8253;
    wire N__8250;
    wire N__8247;
    wire N__8244;
    wire N__8243;
    wire N__8240;
    wire N__8239;
    wire N__8236;
    wire N__8235;
    wire N__8232;
    wire N__8229;
    wire N__8226;
    wire N__8223;
    wire N__8218;
    wire N__8215;
    wire N__8212;
    wire N__8205;
    wire N__8202;
    wire N__8201;
    wire N__8200;
    wire N__8199;
    wire N__8196;
    wire N__8191;
    wire N__8188;
    wire N__8181;
    wire N__8178;
    wire N__8175;
    wire N__8172;
    wire N__8171;
    wire N__8168;
    wire N__8167;
    wire N__8166;
    wire N__8165;
    wire N__8164;
    wire N__8163;
    wire N__8162;
    wire N__8161;
    wire N__8158;
    wire N__8153;
    wire N__8150;
    wire N__8147;
    wire N__8142;
    wire N__8137;
    wire N__8130;
    wire N__8121;
    wire N__8118;
    wire N__8115;
    wire N__8114;
    wire N__8113;
    wire N__8112;
    wire N__8111;
    wire N__8110;
    wire N__8107;
    wire N__8106;
    wire N__8105;
    wire N__8100;
    wire N__8099;
    wire N__8098;
    wire N__8095;
    wire N__8094;
    wire N__8085;
    wire N__8084;
    wire N__8083;
    wire N__8082;
    wire N__8081;
    wire N__8080;
    wire N__8079;
    wire N__8076;
    wire N__8073;
    wire N__8064;
    wire N__8061;
    wire N__8056;
    wire N__8051;
    wire N__8048;
    wire N__8045;
    wire N__8028;
    wire N__8027;
    wire N__8024;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8010;
    wire N__8007;
    wire N__8004;
    wire N__8001;
    wire N__7998;
    wire N__7995;
    wire N__7992;
    wire N__7989;
    wire N__7988;
    wire N__7985;
    wire N__7984;
    wire N__7981;
    wire N__7978;
    wire N__7975;
    wire N__7974;
    wire N__7971;
    wire N__7970;
    wire N__7969;
    wire N__7966;
    wire N__7963;
    wire N__7962;
    wire N__7961;
    wire N__7958;
    wire N__7957;
    wire N__7954;
    wire N__7951;
    wire N__7950;
    wire N__7947;
    wire N__7942;
    wire N__7937;
    wire N__7932;
    wire N__7927;
    wire N__7924;
    wire N__7911;
    wire N__7908;
    wire N__7907;
    wire N__7904;
    wire N__7901;
    wire N__7896;
    wire N__7893;
    wire N__7890;
    wire N__7887;
    wire N__7884;
    wire N__7883;
    wire N__7880;
    wire N__7877;
    wire N__7872;
    wire N__7869;
    wire N__7866;
    wire N__7863;
    wire N__7860;
    wire N__7857;
    wire N__7854;
    wire N__7853;
    wire N__7850;
    wire N__7847;
    wire N__7844;
    wire N__7839;
    wire N__7836;
    wire N__7833;
    wire N__7830;
    wire N__7827;
    wire N__7826;
    wire N__7825;
    wire N__7824;
    wire N__7821;
    wire N__7818;
    wire N__7813;
    wire N__7810;
    wire N__7807;
    wire N__7804;
    wire N__7803;
    wire N__7802;
    wire N__7801;
    wire N__7800;
    wire N__7797;
    wire N__7792;
    wire N__7787;
    wire N__7782;
    wire N__7779;
    wire N__7776;
    wire N__7771;
    wire N__7768;
    wire N__7763;
    wire N__7758;
    wire N__7755;
    wire N__7752;
    wire N__7751;
    wire N__7750;
    wire N__7749;
    wire N__7748;
    wire N__7745;
    wire N__7740;
    wire N__7737;
    wire N__7736;
    wire N__7733;
    wire N__7732;
    wire N__7731;
    wire N__7730;
    wire N__7727;
    wire N__7724;
    wire N__7719;
    wire N__7716;
    wire N__7713;
    wire N__7710;
    wire N__7707;
    wire N__7704;
    wire N__7699;
    wire N__7692;
    wire N__7689;
    wire N__7686;
    wire N__7683;
    wire N__7678;
    wire N__7675;
    wire N__7670;
    wire N__7665;
    wire N__7662;
    wire N__7659;
    wire N__7658;
    wire N__7655;
    wire N__7652;
    wire N__7651;
    wire N__7650;
    wire N__7647;
    wire N__7642;
    wire N__7641;
    wire N__7638;
    wire N__7635;
    wire N__7634;
    wire N__7633;
    wire N__7630;
    wire N__7625;
    wire N__7622;
    wire N__7619;
    wire N__7616;
    wire N__7615;
    wire N__7610;
    wire N__7607;
    wire N__7604;
    wire N__7601;
    wire N__7598;
    wire N__7595;
    wire N__7586;
    wire N__7583;
    wire N__7580;
    wire N__7577;
    wire N__7574;
    wire N__7571;
    wire N__7566;
    wire N__7565;
    wire N__7562;
    wire N__7561;
    wire N__7560;
    wire N__7559;
    wire N__7554;
    wire N__7553;
    wire N__7550;
    wire N__7547;
    wire N__7544;
    wire N__7543;
    wire N__7540;
    wire N__7537;
    wire N__7536;
    wire N__7535;
    wire N__7532;
    wire N__7529;
    wire N__7526;
    wire N__7523;
    wire N__7520;
    wire N__7517;
    wire N__7512;
    wire N__7509;
    wire N__7502;
    wire N__7499;
    wire N__7494;
    wire N__7491;
    wire N__7488;
    wire N__7483;
    wire N__7480;
    wire N__7477;
    wire N__7474;
    wire N__7467;
    wire N__7464;
    wire N__7461;
    wire N__7458;
    wire N__7455;
    wire N__7452;
    wire N__7449;
    wire N__7446;
    wire N__7443;
    wire N__7440;
    wire N__7437;
    wire N__7434;
    wire N__7431;
    wire N__7428;
    wire N__7425;
    wire N__7422;
    wire N__7419;
    wire N__7416;
    wire N__7415;
    wire N__7412;
    wire N__7409;
    wire N__7406;
    wire N__7403;
    wire N__7400;
    wire N__7397;
    wire N__7392;
    wire N__7389;
    wire N__7386;
    wire N__7383;
    wire N__7380;
    wire N__7377;
    wire N__7374;
    wire N__7371;
    wire N__7368;
    wire N__7365;
    wire N__7362;
    wire N__7359;
    wire N__7356;
    wire N__7353;
    wire N__7350;
    wire N__7349;
    wire N__7346;
    wire N__7343;
    wire N__7340;
    wire N__7337;
    wire N__7334;
    wire N__7331;
    wire N__7328;
    wire N__7325;
    wire N__7322;
    wire N__7319;
    wire N__7314;
    wire N__7313;
    wire N__7310;
    wire N__7307;
    wire N__7302;
    wire N__7299;
    wire N__7296;
    wire N__7295;
    wire N__7292;
    wire N__7289;
    wire N__7286;
    wire N__7283;
    wire N__7280;
    wire N__7277;
    wire N__7274;
    wire N__7271;
    wire N__7268;
    wire N__7265;
    wire N__7260;
    wire N__7257;
    wire N__7254;
    wire N__7251;
    wire N__7250;
    wire N__7249;
    wire N__7248;
    wire N__7245;
    wire N__7242;
    wire N__7239;
    wire N__7238;
    wire N__7235;
    wire N__7234;
    wire N__7233;
    wire N__7230;
    wire N__7227;
    wire N__7222;
    wire N__7217;
    wire N__7214;
    wire N__7203;
    wire N__7200;
    wire N__7197;
    wire N__7194;
    wire N__7191;
    wire N__7188;
    wire N__7187;
    wire N__7184;
    wire N__7181;
    wire N__7176;
    wire N__7173;
    wire N__7170;
    wire N__7169;
    wire N__7168;
    wire N__7167;
    wire N__7164;
    wire N__7159;
    wire N__7158;
    wire N__7155;
    wire N__7152;
    wire N__7149;
    wire N__7146;
    wire N__7145;
    wire N__7142;
    wire N__7141;
    wire N__7140;
    wire N__7139;
    wire N__7134;
    wire N__7131;
    wire N__7128;
    wire N__7125;
    wire N__7118;
    wire N__7107;
    wire N__7104;
    wire N__7103;
    wire N__7102;
    wire N__7101;
    wire N__7100;
    wire N__7095;
    wire N__7090;
    wire N__7089;
    wire N__7088;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7074;
    wire N__7065;
    wire N__7062;
    wire N__7059;
    wire N__7056;
    wire N__7053;
    wire N__7050;
    wire N__7047;
    wire N__7046;
    wire N__7043;
    wire N__7040;
    wire N__7035;
    wire N__7032;
    wire N__7029;
    wire N__7026;
    wire N__7023;
    wire N__7020;
    wire N__7017;
    wire N__7014;
    wire N__7013;
    wire N__7010;
    wire N__7007;
    wire N__7004;
    wire N__7001;
    wire N__6998;
    wire N__6995;
    wire N__6992;
    wire N__6989;
    wire N__6986;
    wire N__6981;
    wire N__6978;
    wire N__6975;
    wire N__6972;
    wire N__6969;
    wire N__6968;
    wire N__6965;
    wire N__6962;
    wire N__6959;
    wire N__6956;
    wire N__6953;
    wire N__6950;
    wire N__6945;
    wire N__6942;
    wire N__6941;
    wire N__6940;
    wire N__6939;
    wire N__6936;
    wire N__6933;
    wire N__6926;
    wire N__6921;
    wire N__6918;
    wire N__6915;
    wire N__6912;
    wire N__6909;
    wire N__6906;
    wire N__6903;
    wire N__6900;
    wire N__6897;
    wire N__6894;
    wire N__6891;
    wire N__6888;
    wire N__6885;
    wire N__6882;
    wire N__6879;
    wire N__6876;
    wire N__6875;
    wire N__6870;
    wire N__6867;
    wire N__6864;
    wire N__6861;
    wire N__6858;
    wire N__6855;
    wire N__6854;
    wire N__6853;
    wire N__6852;
    wire N__6851;
    wire N__6850;
    wire N__6849;
    wire N__6840;
    wire N__6839;
    wire N__6836;
    wire N__6831;
    wire N__6828;
    wire N__6825;
    wire N__6822;
    wire N__6821;
    wire N__6818;
    wire N__6813;
    wire N__6810;
    wire N__6807;
    wire N__6802;
    wire N__6795;
    wire N__6794;
    wire N__6789;
    wire N__6786;
    wire N__6783;
    wire N__6780;
    wire N__6777;
    wire N__6774;
    wire N__6773;
    wire N__6770;
    wire N__6767;
    wire N__6762;
    wire N__6759;
    wire N__6756;
    wire N__6753;
    wire N__6750;
    wire N__6747;
    wire N__6746;
    wire N__6743;
    wire N__6740;
    wire N__6735;
    wire N__6734;
    wire N__6731;
    wire N__6728;
    wire N__6725;
    wire N__6720;
    wire N__6717;
    wire N__6714;
    wire N__6711;
    wire N__6708;
    wire N__6705;
    wire N__6704;
    wire N__6701;
    wire N__6698;
    wire N__6693;
    wire N__6690;
    wire N__6687;
    wire N__6684;
    wire N__6681;
    wire N__6678;
    wire N__6677;
    wire N__6674;
    wire N__6671;
    wire N__6666;
    wire N__6663;
    wire N__6660;
    wire N__6657;
    wire N__6654;
    wire N__6651;
    wire N__6648;
    wire N__6647;
    wire N__6644;
    wire N__6641;
    wire N__6636;
    wire N__6633;
    wire N__6630;
    wire N__6629;
    wire N__6626;
    wire N__6623;
    wire N__6620;
    wire N__6615;
    wire N__6612;
    wire N__6609;
    wire N__6608;
    wire N__6607;
    wire N__6606;
    wire N__6605;
    wire N__6602;
    wire N__6597;
    wire N__6592;
    wire N__6585;
    wire N__6584;
    wire N__6583;
    wire N__6582;
    wire N__6581;
    wire N__6578;
    wire N__6577;
    wire N__6574;
    wire N__6571;
    wire N__6568;
    wire N__6565;
    wire N__6562;
    wire N__6561;
    wire N__6560;
    wire N__6559;
    wire N__6558;
    wire N__6553;
    wire N__6550;
    wire N__6545;
    wire N__6542;
    wire N__6535;
    wire N__6532;
    wire N__6519;
    wire N__6516;
    wire N__6513;
    wire N__6510;
    wire N__6507;
    wire N__6504;
    wire N__6501;
    wire N__6498;
    wire N__6495;
    wire N__6492;
    wire N__6489;
    wire N__6486;
    wire N__6483;
    wire N__6480;
    wire N__6477;
    wire N__6474;
    wire N__6471;
    wire N__6468;
    wire N__6465;
    wire N__6462;
    wire N__6459;
    wire N__6456;
    wire N__6453;
    wire N__6450;
    wire N__6449;
    wire N__6446;
    wire N__6441;
    wire N__6438;
    wire N__6435;
    wire N__6432;
    wire N__6429;
    wire N__6426;
    wire N__6423;
    wire N__6420;
    wire N__6417;
    wire N__6414;
    wire N__6411;
    wire N__6408;
    wire N__6405;
    wire N__6402;
    wire N__6399;
    wire N__6396;
    wire N__6393;
    wire N__6390;
    wire N__6387;
    wire N__6384;
    wire N__6381;
    wire N__6378;
    wire N__6375;
    wire N__6372;
    wire N__6369;
    wire N__6366;
    wire N__6363;
    wire N__6360;
    wire N__6357;
    wire N__6354;
    wire N__6353;
    wire N__6350;
    wire N__6349;
    wire N__6348;
    wire N__6345;
    wire N__6342;
    wire N__6339;
    wire N__6334;
    wire N__6333;
    wire N__6330;
    wire N__6327;
    wire N__6324;
    wire N__6321;
    wire N__6312;
    wire N__6309;
    wire N__6306;
    wire N__6303;
    wire N__6300;
    wire N__6297;
    wire N__6294;
    wire N__6291;
    wire N__6288;
    wire N__6285;
    wire N__6282;
    wire N__6279;
    wire N__6276;
    wire N__6273;
    wire N__6270;
    wire N__6269;
    wire N__6266;
    wire N__6263;
    wire N__6258;
    wire N__6255;
    wire N__6254;
    wire N__6251;
    wire N__6248;
    wire N__6243;
    wire N__6240;
    wire N__6239;
    wire N__6236;
    wire N__6233;
    wire N__6232;
    wire N__6229;
    wire N__6226;
    wire N__6223;
    wire N__6220;
    wire N__6215;
    wire N__6212;
    wire N__6209;
    wire N__6206;
    wire N__6203;
    wire N__6198;
    wire N__6197;
    wire N__6194;
    wire N__6191;
    wire N__6188;
    wire N__6183;
    wire N__6180;
    wire N__6179;
    wire N__6178;
    wire N__6173;
    wire N__6170;
    wire N__6167;
    wire N__6162;
    wire N__6159;
    wire N__6156;
    wire N__6153;
    wire N__6150;
    wire N__6149;
    wire N__6146;
    wire N__6143;
    wire N__6140;
    wire N__6135;
    wire N__6132;
    wire N__6129;
    wire N__6126;
    wire N__6123;
    wire N__6120;
    wire N__6117;
    wire N__6116;
    wire N__6113;
    wire N__6110;
    wire N__6107;
    wire N__6104;
    wire N__6101;
    wire N__6098;
    wire N__6095;
    wire N__6092;
    wire N__6089;
    wire N__6086;
    wire N__6081;
    wire N__6078;
    wire N__6075;
    wire N__6072;
    wire N__6069;
    wire N__6066;
    wire N__6063;
    wire N__6060;
    wire N__6057;
    wire N__6054;
    wire N__6051;
    wire N__6048;
    wire N__6045;
    wire N__6042;
    wire N__6039;
    wire N__6036;
    wire N__6033;
    wire N__6030;
    wire N__6027;
    wire N__6024;
    wire N__6021;
    wire N__6018;
    wire N__6015;
    wire N__6012;
    wire N__6009;
    wire N__6006;
    wire N__6003;
    wire N__6000;
    wire N__5997;
    wire N__5994;
    wire N__5991;
    wire N__5988;
    wire N__5985;
    wire N__5982;
    wire N__5979;
    wire N__5976;
    wire N__5973;
    wire N__5970;
    wire N__5967;
    wire N__5964;
    wire N__5961;
    wire N__5958;
    wire N__5957;
    wire N__5954;
    wire N__5951;
    wire N__5946;
    wire N__5945;
    wire N__5942;
    wire N__5937;
    wire N__5934;
    wire N__5931;
    wire N__5928;
    wire N__5925;
    wire N__5922;
    wire N__5919;
    wire N__5918;
    wire N__5915;
    wire N__5912;
    wire N__5907;
    wire N__5904;
    wire N__5901;
    wire N__5898;
    wire N__5895;
    wire N__5892;
    wire N__5889;
    wire N__5886;
    wire N__5883;
    wire N__5880;
    wire N__5877;
    wire N__5874;
    wire N__5871;
    wire N__5868;
    wire N__5865;
    wire N__5862;
    wire N__5861;
    wire N__5860;
    wire N__5855;
    wire N__5852;
    wire N__5849;
    wire N__5846;
    wire N__5843;
    wire N__5840;
    wire N__5835;
    wire N__5832;
    wire N__5829;
    wire N__5826;
    wire N__5823;
    wire N__5820;
    wire N__5817;
    wire N__5814;
    wire N__5811;
    wire N__5808;
    wire N__5805;
    wire N__5802;
    wire N__5799;
    wire N__5796;
    wire N__5793;
    wire N__5792;
    wire N__5787;
    wire N__5784;
    wire N__5781;
    wire N__5778;
    wire N__5775;
    wire N__5772;
    wire N__5769;
    wire N__5766;
    wire N__5763;
    wire N__5760;
    wire N__5757;
    wire N__5754;
    wire N__5751;
    wire N__5748;
    wire N__5745;
    wire N__5742;
    wire N__5739;
    wire N__5736;
    wire N__5733;
    wire N__5730;
    wire N__5727;
    wire N__5724;
    wire N__5721;
    wire N__5718;
    wire N__5715;
    wire N__5712;
    wire N__5709;
    wire N__5706;
    wire N__5705;
    wire N__5702;
    wire N__5699;
    wire N__5696;
    wire N__5691;
    wire N__5688;
    wire N__5685;
    wire N__5682;
    wire N__5679;
    wire N__5676;
    wire N__5673;
    wire N__5670;
    wire N__5667;
    wire N__5664;
    wire N__5663;
    wire N__5662;
    wire N__5659;
    wire N__5656;
    wire N__5653;
    wire N__5652;
    wire N__5651;
    wire N__5650;
    wire N__5649;
    wire N__5648;
    wire N__5645;
    wire N__5640;
    wire N__5635;
    wire N__5628;
    wire N__5619;
    wire N__5616;
    wire N__5613;
    wire N__5610;
    wire N__5609;
    wire N__5606;
    wire N__5603;
    wire N__5600;
    wire N__5595;
    wire N__5592;
    wire N__5589;
    wire N__5586;
    wire N__5583;
    wire N__5580;
    wire N__5577;
    wire N__5574;
    wire N__5571;
    wire N__5568;
    wire N__5565;
    wire N__5562;
    wire N__5559;
    wire N__5556;
    wire N__5553;
    wire N__5550;
    wire N__5549;
    wire N__5544;
    wire N__5541;
    wire N__5538;
    wire N__5537;
    wire N__5534;
    wire N__5531;
    wire N__5530;
    wire N__5527;
    wire N__5524;
    wire N__5521;
    wire N__5514;
    wire N__5511;
    wire N__5508;
    wire N__5505;
    wire N__5504;
    wire N__5501;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5489;
    wire N__5486;
    wire N__5483;
    wire N__5480;
    wire N__5479;
    wire N__5476;
    wire N__5473;
    wire N__5470;
    wire N__5465;
    wire N__5462;
    wire N__5457;
    wire N__5454;
    wire N__5453;
    wire N__5452;
    wire N__5449;
    wire N__5446;
    wire N__5443;
    wire N__5442;
    wire N__5437;
    wire N__5432;
    wire N__5427;
    wire N__5424;
    wire N__5421;
    wire N__5418;
    wire N__5417;
    wire N__5416;
    wire N__5415;
    wire N__5412;
    wire N__5409;
    wire N__5404;
    wire N__5397;
    wire N__5396;
    wire N__5395;
    wire N__5390;
    wire N__5387;
    wire N__5384;
    wire N__5379;
    wire N__5378;
    wire N__5373;
    wire N__5370;
    wire N__5367;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5359;
    wire N__5356;
    wire N__5353;
    wire N__5350;
    wire N__5343;
    wire N__5342;
    wire N__5341;
    wire N__5340;
    wire N__5337;
    wire N__5336;
    wire N__5333;
    wire N__5328;
    wire N__5325;
    wire N__5322;
    wire N__5313;
    wire N__5312;
    wire N__5311;
    wire N__5310;
    wire N__5307;
    wire N__5304;
    wire N__5299;
    wire N__5292;
    wire N__5291;
    wire N__5290;
    wire N__5289;
    wire N__5288;
    wire N__5285;
    wire N__5280;
    wire N__5275;
    wire N__5268;
    wire N__5265;
    wire N__5262;
    wire N__5261;
    wire N__5258;
    wire N__5257;
    wire N__5254;
    wire N__5251;
    wire N__5248;
    wire N__5245;
    wire N__5242;
    wire N__5239;
    wire N__5236;
    wire N__5233;
    wire N__5230;
    wire N__5229;
    wire N__5226;
    wire N__5223;
    wire N__5220;
    wire N__5219;
    wire N__5216;
    wire N__5213;
    wire N__5210;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5194;
    wire N__5191;
    wire N__5188;
    wire N__5181;
    wire N__5178;
    wire N__5175;
    wire N__5172;
    wire N__5169;
    wire N__5166;
    wire N__5163;
    wire N__5160;
    wire N__5157;
    wire N__5154;
    wire N__5151;
    wire N__5148;
    wire N__5145;
    wire N__5142;
    wire N__5139;
    wire N__5136;
    wire N__5133;
    wire N__5132;
    wire N__5131;
    wire N__5128;
    wire N__5125;
    wire N__5122;
    wire N__5115;
    wire N__5112;
    wire N__5109;
    wire N__5106;
    wire N__5103;
    wire N__5100;
    wire N__5097;
    wire N__5094;
    wire N__5091;
    wire N__5088;
    wire N__5085;
    wire N__5084;
    wire N__5081;
    wire N__5078;
    wire N__5075;
    wire N__5070;
    wire N__5067;
    wire N__5064;
    wire N__5061;
    wire N__5058;
    wire N__5055;
    wire N__5052;
    wire N__5049;
    wire N__5046;
    wire N__5043;
    wire N__5040;
    wire N__5039;
    wire N__5036;
    wire N__5033;
    wire N__5030;
    wire N__5027;
    wire N__5024;
    wire N__5021;
    wire N__5018;
    wire N__5015;
    wire N__5010;
    wire N__5007;
    wire N__5004;
    wire N__5001;
    wire N__5000;
    wire N__4997;
    wire N__4994;
    wire N__4989;
    wire N__4986;
    wire N__4983;
    wire N__4980;
    wire N__4977;
    wire N__4974;
    wire N__4971;
    wire N__4970;
    wire N__4969;
    wire N__4966;
    wire N__4961;
    wire N__4956;
    wire N__4955;
    wire N__4952;
    wire N__4951;
    wire N__4948;
    wire N__4943;
    wire N__4942;
    wire N__4937;
    wire N__4934;
    wire N__4931;
    wire N__4926;
    wire N__4925;
    wire N__4924;
    wire N__4923;
    wire N__4922;
    wire N__4919;
    wire N__4910;
    wire N__4905;
    wire N__4902;
    wire N__4901;
    wire N__4898;
    wire N__4895;
    wire N__4894;
    wire N__4891;
    wire N__4888;
    wire N__4885;
    wire N__4882;
    wire N__4879;
    wire N__4876;
    wire N__4873;
    wire N__4870;
    wire N__4867;
    wire N__4864;
    wire N__4861;
    wire N__4858;
    wire N__4857;
    wire N__4850;
    wire N__4847;
    wire N__4842;
    wire N__4839;
    wire N__4836;
    wire N__4833;
    wire N__4830;
    wire N__4827;
    wire N__4824;
    wire N__4821;
    wire N__4818;
    wire N__4815;
    wire N__4812;
    wire N__4811;
    wire N__4806;
    wire N__4803;
    wire N__4800;
    wire N__4797;
    wire N__4794;
    wire N__4791;
    wire N__4788;
    wire N__4785;
    wire N__4782;
    wire N__4779;
    wire N__4778;
    wire N__4775;
    wire N__4772;
    wire N__4767;
    wire N__4764;
    wire N__4761;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4748;
    wire N__4745;
    wire N__4742;
    wire N__4739;
    wire N__4736;
    wire N__4733;
    wire N__4732;
    wire N__4727;
    wire N__4724;
    wire N__4719;
    wire N__4716;
    wire N__4713;
    wire N__4710;
    wire N__4707;
    wire N__4704;
    wire N__4701;
    wire N__4698;
    wire N__4697;
    wire N__4692;
    wire N__4689;
    wire N__4688;
    wire N__4685;
    wire N__4682;
    wire N__4677;
    wire N__4676;
    wire N__4673;
    wire N__4670;
    wire N__4665;
    wire N__4664;
    wire N__4661;
    wire N__4658;
    wire N__4655;
    wire N__4650;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4638;
    wire N__4635;
    wire N__4632;
    wire N__4629;
    wire N__4628;
    wire N__4625;
    wire N__4622;
    wire N__4617;
    wire N__4614;
    wire N__4611;
    wire N__4608;
    wire N__4605;
    wire N__4602;
    wire N__4599;
    wire N__4596;
    wire N__4593;
    wire N__4590;
    wire N__4587;
    wire N__4584;
    wire N__4583;
    wire N__4582;
    wire N__4581;
    wire N__4580;
    wire N__4579;
    wire N__4578;
    wire N__4563;
    wire N__4560;
    wire N__4557;
    wire N__4556;
    wire N__4553;
    wire N__4550;
    wire N__4545;
    wire N__4544;
    wire N__4541;
    wire N__4538;
    wire N__4533;
    wire N__4530;
    wire N__4527;
    wire N__4524;
    wire N__4521;
    wire N__4520;
    wire N__4517;
    wire N__4514;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4502;
    wire N__4497;
    wire N__4494;
    wire N__4491;
    wire N__4488;
    wire N__4485;
    wire N__4484;
    wire N__4481;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4463;
    wire N__4460;
    wire N__4457;
    wire N__4452;
    wire N__4449;
    wire N__4446;
    wire N__4443;
    wire N__4440;
    wire N__4437;
    wire N__4434;
    wire N__4431;
    wire N__4428;
    wire N__4425;
    wire N__4422;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4407;
    wire N__4404;
    wire N__4401;
    wire N__4398;
    wire N__4395;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire CLK80_PLL_i_i;
    wire DBRn_c_i_cascade_;
    wire DBRn_c_i_0;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire bfn_10_6_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire C1_c_g;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire C3_c;
    wire DBRn_c;
    wire N_58_i;
    wire \U712_BYTE_ENABLE.N_352 ;
    wire \INVU712_CYCLE_TERM.TACK_ENC_net ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ;
    wire DBDIR_c;
    wire DBR_SYNCZ0Z_0;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_4 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_5 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_6 ;
    wire PRnW_c;
    wire \U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1 ;
    wire BLSn_c;
    wire REG_TACK;
    wire VBENn_c;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_CYCLE_TERM.TACK_STARTZ0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_CYCLE_TERM.N_36_0_cascade_ ;
    wire TACK_OUT;
    wire \INVU712_CYCLE_TERM.TACK_STATE_0C_net ;
    wire A_c_16;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_ ;
    wire CMA_c_1;
    wire \U712_REG_SM.START_RSTZ0 ;
    wire REGSPACEn_c;
    wire \U712_REG_SM.N_455_cascade_ ;
    wire A_c_10;
    wire \U712_CHIP_RAM.N_387 ;
    wire \U712_REG_SM.N_185_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_7 ;
    wire \U712_REG_SM.N_368_cascade_ ;
    wire \U712_CHIP_RAM.N_378 ;
    wire \U712_REG_SM.N_441 ;
    wire \U712_REG_SM.N_358_cascade_ ;
    wire \U712_REG_SM.N_368 ;
    wire \U712_REG_SM.N_366 ;
    wire \U712_REG_SM.N_366_cascade_ ;
    wire \U712_REG_SM.un1_STATE_COUNT_1_sqmuxa_0 ;
    wire CLK40_PLL;
    wire CLK40_PLL_iso_i;
    wire \U712_REG_SM.WRITE_CYCLEZ0 ;
    wire \U712_REG_SM.N_375 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_0 ;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.N_483 ;
    wire \U712_REG_SM.N_483_cascade_ ;
    wire \U712_REG_SM.N_367 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_1 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire \U712_REG_SM.N_358 ;
    wire \U712_REG_SM.N_592 ;
    wire TACK_EN;
    wire \U712_CYCLE_TERM.TACK_RST_0_i ;
    wire RESETn_c_i;
    wire A_c_15;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.N_407 ;
    wire \U712_REG_SM.N_369_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_2 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0 ;
    wire A_c_17;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8 ;
    wire \U712_CHIP_RAM.un1_CMA25_0_i_cascade_ ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_3 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_4 ;
    wire A_c_8;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ;
    wire A_c_18;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ;
    wire A_c_20;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ;
    wire \U712_REG_SM.N_481 ;
    wire LDSn_c;
    wire \U712_REG_SM.N_185 ;
    wire UDSn_c;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_0Z0Z_0 ;
    wire \U712_BYTE_ENABLE.N_468 ;
    wire N_65_i;
    wire \U712_BYTE_ENABLE.N_343_i ;
    wire \U712_BYTE_ENABLE.N_466_cascade_ ;
    wire N_67_i;
    wire ASn_c;
    wire \U712_REG_SM.N_185_0 ;
    wire \U712_REG_SM.N_482 ;
    wire C1_c;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ;
    wire CMA_c_7;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8 ;
    wire CMA_c_8;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire \U712_CHIP_RAM.N_362_cascade_ ;
    wire \U712_CHIP_RAM.N_493_cascade_ ;
    wire \U712_CHIP_RAM.N_503_cascade_ ;
    wire \U712_CHIP_RAM.N_596_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.N_596 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0 ;
    wire AWEn_c;
    wire \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_i_i_a2_0_cascade_ ;
    wire \U712_CHIP_RAM.WRITE_CYCLEZ0 ;
    wire \U712_CHIP_RAM.N_365 ;
    wire \U712_CHIP_RAM.N_365_cascade_ ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_ ;
    wire A_c_2;
    wire A_c_3;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ;
    wire A_c_4;
    wire A_c_7;
    wire DBENn_c;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_1Z0Z_0 ;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_1Z0Z_0_cascade_ ;
    wire N_62_i;
    wire \U712_CHIP_RAM.N_452_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_0_2 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_1_cascade_ ;
    wire \U712_REG_SM.N_406 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_8 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire \U712_REG_SM.N_445_cascade_ ;
    wire \U712_REG_SM.REG_CYCLE_5_iv_0_0 ;
    wire \U712_BYTE_ENABLE.LMBE_0_i_o3_0_oZ0Z2 ;
    wire N_282_i;
    wire N_219;
    wire N_60_i;
    wire \U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ;
    wire DBR_SYNC_i_1;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0 ;
    wire bfn_15_4_0_;
    wire \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2 ;
    wire \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3_cascade_ ;
    wire \U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3 ;
    wire \U712_CHIP_RAM.N_451_cascade_ ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1 ;
    wire DBR_SYNCZ0Z_1;
    wire \U712_CHIP_RAM.CAS_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.N_362 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_165_i_i_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_o2_0_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_a2_1_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER19 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0 ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0 ;
    wire \U712_CHIP_RAM.N_344_cascade_ ;
    wire \U712_CHIP_RAM.N_435 ;
    wire \U712_CHIP_RAM.N_430 ;
    wire \U712_CHIP_RAM.N_347_cascade_ ;
    wire \U712_CHIP_RAM.N_590 ;
    wire \U712_CHIP_RAM.N_590_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0 ;
    wire \U712_CHIP_RAM.N_509_cascade_ ;
    wire \U712_CHIP_RAM.DBENn_8_0_0 ;
    wire TSn_c;
    wire \U712_CHIP_RAM.N_458_cascade_ ;
    wire RAMENn_c;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3 ;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ;
    wire A_c_11;
    wire \U712_CHIP_RAM.N_350 ;
    wire \U712_CHIP_RAM.N_452 ;
    wire A_c_9;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a2_1_cascade_ ;
    wire \U712_CHIP_RAM.N_344 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_0 ;
    wire \U712_CHIP_RAM.N_72_cascade_ ;
    wire CPU_TACKm;
    wire \U712_CHIP_RAM.N_462 ;
    wire \U712_CHIP_RAM.N_503 ;
    wire \U712_CHIP_RAM.N_462_cascade_ ;
    wire \U712_CHIP_RAM.N_510 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0_cascade_ ;
    wire LATCH_CLK_c;
    wire DBRn_c_i;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ;
    wire N_119_i;
    wire A_c_1;
    wire A_c_0;
    wire SIZ_c_0;
    wire SIZ_c_1;
    wire N_61_i;
    wire CMA_c_2;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ;
    wire CONSTANT_ONE_NET;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_0 ;
    wire \U712_CHIP_RAM.N_431 ;
    wire \U712_CHIP_RAM.N_359 ;
    wire \U712_CHIP_RAM.N_595 ;
    wire \U712_CHIP_RAM.N_348 ;
    wire \U712_CHIP_RAM.N_595_cascade_ ;
    wire \U712_CHIP_RAM.N_577 ;
    wire \U712_CHIP_RAM.N_279 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_i_a2_0_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_a2_0 ;
    wire bfn_16_6_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.N_132_i ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.N_436 ;
    wire \U712_CHIP_RAM.N_499 ;
    wire DMA_CYCLEm;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.N_506_cascade_ ;
    wire \U712_CHIP_RAM.N_147_i_i_a2_0 ;
    wire \U712_CHIP_RAM.N_147_i_i_a2_0_cascade_ ;
    wire \U712_CHIP_RAM.N_500_i ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH5lto7_0 ;
    wire \U712_CHIP_RAM.REFRESH5lt7 ;
    wire \U712_CHIP_RAM.N_509 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_508 ;
    wire \U712_CHIP_RAM.N_494 ;
    wire A_c_12;
    wire A_c_13;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ;
    wire A_c_5;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ;
    wire A_c_6;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ;
    wire REG_CYCLEm;
    wire N_207_i;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire A_c_14;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ;
    wire CMA_c_0;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire DRA_c_7;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \INVU712_CHIP_RAM.DMA_A1_nesrC_net ;
    wire RASn_c;
    wire CRCSn_c;
    wire CASn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CMA_c_10;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire \U712_CHIP_RAM.N_354_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ;
    wire CMA_c_5;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire CMA_c_3;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire DRA_c_1;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire WEn_c;
    wire \U712_CHIP_RAM.CMA_5_i_0_9 ;
    wire A_c_19;
    wire CPU_CYCLEm;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.N_354 ;
    wire \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ;
    wire CMA_c_4;
    wire \U712_CHIP_RAM.un1_CMA25_0_i_0 ;
    wire DRA_c_9;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_2 ;
    wire RAS0n_c;
    wire RAS1n_c;
    wire RESETn_c;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_1 ;
    wire CLK80_PLL;
    wire DRA_c_3;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire DRA_c_5;
    wire DRA_c_6;
    wire AGNUS_REV_c;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire C3_c_g;
    wire DBRn_c_i_0_g;
    wire RESETn_c_i_g;
    wire RnW_c;
    wire CASUn_c;
    wire DMA_WRITE_CYCLE;
    wire CASLn_c;
    wire N_409;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL),
            .REFERENCECLK(N__4413),
            .RESETB(N__7416),
            .BYPASS(GNDG0),
            .PLLOUTCOREA(),
            .SDI(GNDG0),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(GNDG0),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK(GNDG0));
    IO_PAD DBENn_obuf_iopad (
            .OE(N__12997),
            .DIN(N__12996),
            .DOUT(N__12995),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__12997),
            .PADOUT(N__12996),
            .PADIN(N__12995),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6363),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__12988),
            .DIN(N__12987),
            .DOUT(N__12986),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__12988),
            .PADOUT(N__12987),
            .PADIN(N__12986),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__12979),
            .DIN(N__12978),
            .DOUT(N__12977),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__12979),
            .PADOUT(N__12978),
            .PADIN(N__12977),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9399),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__12970),
            .DIN(N__12969),
            .DOUT(N__12968),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__12970),
            .PADOUT(N__12969),
            .PADIN(N__12968),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10707),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__12961),
            .DIN(N__12960),
            .DOUT(N__12959),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__12961),
            .PADOUT(N__12960),
            .PADIN(N__12959),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__12952),
            .DIN(N__12951),
            .DOUT(N__12950),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__12952),
            .PADOUT(N__12951),
            .PADIN(N__12950),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__12943),
            .DIN(N__12942),
            .DOUT(N__12941),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__12943),
            .PADOUT(N__12942),
            .PADIN(N__12941),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__12934),
            .DIN(N__12933),
            .DOUT(N__12932),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__12934),
            .PADOUT(N__12933),
            .PADIN(N__12932),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__12925),
            .DIN(N__12924),
            .DOUT(N__12923),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__12925),
            .PADOUT(N__12924),
            .PADIN(N__12923),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS1n_ibuf_iopad (
            .OE(N__12916),
            .DIN(N__12915),
            .DOUT(N__12914),
            .PACKAGEPIN(RAS1n));
    defparam RAS1n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS1n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS1n_ibuf_preio (
            .PADOEN(N__12916),
            .PADOUT(N__12915),
            .PADIN(N__12914),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS1n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__12907),
            .DIN(N__12906),
            .DOUT(N__12905),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__12907),
            .PADOUT(N__12906),
            .PADIN(N__12905),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__12898),
            .DIN(N__12897),
            .DOUT(N__12896),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__12898),
            .PADOUT(N__12897),
            .PADIN(N__12896),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6033),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__12889),
            .DIN(N__12888),
            .DOUT(N__12887),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__12889),
            .PADOUT(N__12888),
            .PADIN(N__12887),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6465),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__12880),
            .DIN(N__12879),
            .DOUT(N__12878),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__12880),
            .PADOUT(N__12879),
            .PADIN(N__12878),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMENn_obuf_iopad (
            .OE(N__12871),
            .DIN(N__12870),
            .DOUT(N__12869),
            .PACKAGEPIN(RAMENn));
    defparam RAMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMENn_obuf_preio (
            .PADOEN(N__12871),
            .PADOUT(N__12870),
            .PADIN(N__12869),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6968),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__12862),
            .DIN(N__12861),
            .DOUT(N__12860),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__12862),
            .PADOUT(N__12861),
            .PADIN(N__12860),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__12853),
            .DIN(N__12852),
            .DOUT(N__12851),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__12853),
            .PADOUT(N__12852),
            .PADIN(N__12851),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__12844),
            .DIN(N__12843),
            .DOUT(N__12842),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__12844),
            .PADOUT(N__12843),
            .PADIN(N__12842),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4989),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__12835),
            .DIN(N__12834),
            .DOUT(N__12833),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__12835),
            .PADOUT(N__12834),
            .PADIN(N__12833),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__12826),
            .DIN(N__12825),
            .DOUT(N__12824),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__12826),
            .PADOUT(N__12825),
            .PADIN(N__12824),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__12817),
            .DIN(N__12816),
            .DOUT(N__12815),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__12817),
            .PADOUT(N__12816),
            .PADIN(N__12815),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9222),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__12808),
            .DIN(N__12807),
            .DOUT(N__12806),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__12808),
            .PADOUT(N__12807),
            .PADIN(N__12806),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__12799),
            .DIN(N__12798),
            .DOUT(N__12797),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__12799),
            .PADOUT(N__12798),
            .PADIN(N__12797),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9417),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__12790),
            .DIN(N__12789),
            .DOUT(N__12788),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__12790),
            .PADOUT(N__12789),
            .PADIN(N__12788),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__12781),
            .DIN(N__12780),
            .DOUT(N__12779),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__12781),
            .PADOUT(N__12780),
            .PADIN(N__12779),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6480),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_obuft_iopad (
            .OE(N__12772),
            .DIN(N__12771),
            .DOUT(N__12770),
            .PACKAGEPIN(TBIn));
    defparam TBIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TBIn_obuft_preio (
            .PADOEN(N__12772),
            .PADOUT(N__12771),
            .PADIN(N__12770),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5257),
            .DIN0(),
            .DOUT0(N__4894),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__12763),
            .DIN(N__12762),
            .DOUT(N__12761),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__12763),
            .PADOUT(N__12762),
            .PADIN(N__12761),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__12754),
            .DIN(N__12753),
            .DOUT(N__12752),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__12754),
            .PADOUT(N__12753),
            .PADIN(N__12752),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__12745),
            .DIN(N__12744),
            .DOUT(N__12743),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__12745),
            .PADOUT(N__12744),
            .PADIN(N__12743),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__12736),
            .DIN(N__12735),
            .DOUT(N__12734),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__12736),
            .PADOUT(N__12735),
            .PADIN(N__12734),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__12727),
            .DIN(N__12726),
            .DOUT(N__12725),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__12727),
            .PADOUT(N__12726),
            .PADIN(N__12725),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_EN_obuf_iopad (
            .OE(N__12718),
            .DIN(N__12717),
            .DOUT(N__12716),
            .PACKAGEPIN(DMA_LATCH_EN));
    defparam DMA_LATCH_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_EN_obuf_preio (
            .PADOEN(N__12718),
            .PADOUT(N__12717),
            .PADIN(N__12716),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6501),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__12709),
            .DIN(N__12708),
            .DOUT(N__12707),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__12709),
            .PADOUT(N__12708),
            .PADIN(N__12707),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__12700),
            .DIN(N__12699),
            .DOUT(N__12698),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__12700),
            .PADOUT(N__12699),
            .PADIN(N__12698),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__12691),
            .DIN(N__12690),
            .DOUT(N__12689),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__12691),
            .PADOUT(N__12690),
            .PADIN(N__12689),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__12682),
            .DIN(N__12681),
            .DOUT(N__12680),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__12682),
            .PADOUT(N__12681),
            .PADIN(N__12680),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__12673),
            .DIN(N__12672),
            .DOUT(N__12671),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__12673),
            .PADOUT(N__12672),
            .PADIN(N__12671),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__12664),
            .DIN(N__12663),
            .DOUT(N__12662),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__12664),
            .PADOUT(N__12663),
            .PADIN(N__12662),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9432),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__12655),
            .DIN(N__12654),
            .DOUT(N__12653),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__12655),
            .PADOUT(N__12654),
            .PADIN(N__12653),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__12646),
            .DIN(N__12645),
            .DOUT(N__12644),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__12646),
            .PADOUT(N__12645),
            .PADIN(N__12644),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__12637),
            .DIN(N__12636),
            .DOUT(N__12635),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__12637),
            .PADOUT(N__12636),
            .PADIN(N__12635),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5817),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_0_iopad (
            .OE(N__12628),
            .DIN(N__12627),
            .DOUT(N__12626),
            .PACKAGEPIN(DA[0]));
    defparam DA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_0_preio (
            .PADOEN(N__12628),
            .PADOUT(N__12627),
            .PADIN(N__12626),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7296),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__12619),
            .DIN(N__12618),
            .DOUT(N__12617),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__12619),
            .PADOUT(N__12618),
            .PADIN(N__12617),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__12610),
            .DIN(N__12609),
            .DOUT(N__12608),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__12610),
            .PADOUT(N__12609),
            .PADIN(N__12608),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9924),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__12601),
            .DIN(N__12600),
            .DOUT(N__12599),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__12601),
            .PADOUT(N__12600),
            .PADIN(N__12599),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10134),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__12592),
            .DIN(N__12591),
            .DOUT(N__12590),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__12592),
            .PADOUT(N__12591),
            .PADIN(N__12590),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4761),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__12583),
            .DIN(N__12582),
            .DOUT(N__12581),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__12583),
            .PADOUT(N__12582),
            .PADIN(N__12581),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__12574),
            .DIN(N__12573),
            .DOUT(N__12572),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__12574),
            .PADOUT(N__12573),
            .PADIN(N__12572),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__12565),
            .DIN(N__12564),
            .DOUT(N__12563),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__12565),
            .PADOUT(N__12564),
            .PADIN(N__12563),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6303),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_obuft_iopad (
            .OE(N__12556),
            .DIN(N__12555),
            .DOUT(N__12554),
            .PACKAGEPIN(TCIn));
    defparam TCIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TCIn_obuft_preio (
            .PADOEN(N__12556),
            .PADOUT(N__12555),
            .PADIN(N__12554),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5262),
            .DIN0(),
            .DOUT0(N__4901),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__12547),
            .DIN(N__12546),
            .DOUT(N__12545),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__12547),
            .PADOUT(N__12546),
            .PADIN(N__12545),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10572),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__12538),
            .DIN(N__12537),
            .DOUT(N__12536),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__12538),
            .PADOUT(N__12537),
            .PADIN(N__12536),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4638),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__12529),
            .DIN(N__12528),
            .DOUT(N__12527),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__12529),
            .PADOUT(N__12528),
            .PADIN(N__12527),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5886),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__12520),
            .DIN(N__12519),
            .DOUT(N__12518),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__12520),
            .PADOUT(N__12519),
            .PADIN(N__12518),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__12511),
            .DIN(N__12510),
            .DOUT(N__12509),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__12511),
            .PADOUT(N__12510),
            .PADIN(N__12509),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_2_iopad (
            .OE(N__12502),
            .DIN(N__12501),
            .DOUT(N__12500),
            .PACKAGEPIN(DA[2]));
    defparam DA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_2_preio (
            .PADOEN(N__12502),
            .PADOUT(N__12501),
            .PADIN(N__12500),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7359),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__12493),
            .DIN(N__12492),
            .DOUT(N__12491),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__12493),
            .PADOUT(N__12492),
            .PADIN(N__12491),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__12484),
            .DIN(N__12483),
            .DOUT(N__12482),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__12484),
            .PADOUT(N__12483),
            .PADIN(N__12482),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__12475),
            .DIN(N__12474),
            .DOUT(N__12473),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__12475),
            .PADOUT(N__12474),
            .PADIN(N__12473),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5097),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__12466),
            .DIN(N__12465),
            .DOUT(N__12464),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__12466),
            .PADOUT(N__12465),
            .PADIN(N__12464),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7467),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__12457),
            .DIN(N__12456),
            .DOUT(N__12455),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__12457),
            .PADOUT(N__12456),
            .PADIN(N__12455),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__12448),
            .DIN(N__12447),
            .DOUT(N__12446),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__12448),
            .PADOUT(N__12447),
            .PADIN(N__12446),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5832),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__12439),
            .DIN(N__12438),
            .DOUT(N__12437),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__12439),
            .PADOUT(N__12438),
            .PADIN(N__12437),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5261),
            .DIN0(),
            .DOUT0(N__4902),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__12430),
            .DIN(N__12429),
            .DOUT(N__12428),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__12430),
            .PADOUT(N__12429),
            .PADIN(N__12428),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7455),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__12421),
            .DIN(N__12420),
            .DOUT(N__12419),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__12421),
            .PADOUT(N__12420),
            .PADIN(N__12419),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__12412),
            .DIN(N__12411),
            .DOUT(N__12410),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__12412),
            .PADOUT(N__12411),
            .PADIN(N__12410),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__12403),
            .DIN(N__12402),
            .DOUT(N__12401),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__12403),
            .PADOUT(N__12402),
            .PADIN(N__12401),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6006),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__12394),
            .DIN(N__12393),
            .DOUT(N__12392),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__12394),
            .PADOUT(N__12393),
            .PADIN(N__12392),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__12385),
            .DIN(N__12384),
            .DOUT(N__12383),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__12385),
            .PADOUT(N__12384),
            .PADIN(N__12383),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_1_iopad (
            .OE(N__12376),
            .DIN(N__12375),
            .DOUT(N__12374),
            .PACKAGEPIN(DA[1]));
    defparam DA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_1_preio (
            .PADOEN(N__12376),
            .PADOUT(N__12375),
            .PADIN(N__12374),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5049),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__12367),
            .DIN(N__12366),
            .DOUT(N__12365),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__12367),
            .PADOUT(N__12366),
            .PADIN(N__12365),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__12358),
            .DIN(N__12357),
            .DOUT(N__12356),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__12358),
            .PADOUT(N__12357),
            .PADIN(N__12356),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__12349),
            .DIN(N__12348),
            .DOUT(N__12347),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__12349),
            .PADOUT(N__12348),
            .PADIN(N__12347),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9660),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__12340),
            .DIN(N__12339),
            .DOUT(N__12338),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__12340),
            .PADOUT(N__12339),
            .PADIN(N__12338),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5934),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__12331),
            .DIN(N__12330),
            .DOUT(N__12329),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__12331),
            .PADOUT(N__12330),
            .PADIN(N__12329),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7839),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__12322),
            .DIN(N__12321),
            .DOUT(N__12320),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__12322),
            .PADOUT(N__12321),
            .PADIN(N__12320),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6912),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__12313),
            .DIN(N__12312),
            .DOUT(N__12311),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__12313),
            .PADOUT(N__12312),
            .PADIN(N__12311),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__12304),
            .DIN(N__12303),
            .DOUT(N__12302),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__12304),
            .PADOUT(N__12303),
            .PADIN(N__12302),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__12295),
            .DIN(N__12294),
            .DOUT(N__12293),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__12295),
            .PADOUT(N__12294),
            .PADIN(N__12293),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6063),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__12286),
            .DIN(N__12285),
            .DOUT(N__12284),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__12286),
            .PADOUT(N__12285),
            .PADIN(N__12284),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__12277),
            .DIN(N__12276),
            .DOUT(N__12275),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__12277),
            .PADOUT(N__12276),
            .PADIN(N__12275),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__12268),
            .DIN(N__12267),
            .DOUT(N__12266),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__12268),
            .PADOUT(N__12267),
            .PADIN(N__12266),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7893),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__12259),
            .DIN(N__12258),
            .DOUT(N__12257),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__12259),
            .PADOUT(N__12258),
            .PADIN(N__12257),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5973),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__12250),
            .DIN(N__12249),
            .DOUT(N__12248),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__12250),
            .PADOUT(N__12249),
            .PADIN(N__12248),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5505),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PRnW_obuf_iopad (
            .OE(N__12241),
            .DIN(N__12240),
            .DOUT(N__12239),
            .PACKAGEPIN(PRnW));
    defparam PRnW_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PRnW_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PRnW_obuf_preio (
            .PADOEN(N__12241),
            .PADOUT(N__12240),
            .PADIN(N__12239),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4797),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__12232),
            .DIN(N__12231),
            .DOUT(N__12230),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__12232),
            .PADOUT(N__12231),
            .PADIN(N__12230),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__12223),
            .DIN(N__12222),
            .DOUT(N__12221),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__12223),
            .PADOUT(N__12222),
            .PADIN(N__12221),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5504),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__12214),
            .DIN(N__12213),
            .DOUT(N__12212),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__12214),
            .PADOUT(N__12213),
            .PADIN(N__12212),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4452),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__12205),
            .DIN(N__12204),
            .DOUT(N__12203),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__12205),
            .PADOUT(N__12204),
            .PADIN(N__12203),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9633),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__12196),
            .DIN(N__12195),
            .DOUT(N__12194),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__12196),
            .PADOUT(N__12195),
            .PADIN(N__12194),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__12187),
            .DIN(N__12186),
            .DOUT(N__12185),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__12187),
            .PADOUT(N__12186),
            .PADIN(N__12185),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__12178),
            .DIN(N__12177),
            .DOUT(N__12176),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__12178),
            .PADOUT(N__12177),
            .PADIN(N__12176),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BLSn_obuf_iopad (
            .OE(N__12169),
            .DIN(N__12168),
            .DOUT(N__12167),
            .PACKAGEPIN(BLSn));
    defparam BLSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BLSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BLSn_obuf_preio (
            .PADOEN(N__12169),
            .PADOUT(N__12168),
            .PADIN(N__12167),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4760),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__12160),
            .DIN(N__12159),
            .DOUT(N__12158),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__12160),
            .PADOUT(N__12159),
            .PADIN(N__12158),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__12151),
            .DIN(N__12150),
            .DOUT(N__12149),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__12151),
            .PADOUT(N__12150),
            .PADIN(N__12149),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5479),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__12142),
            .DIN(N__12141),
            .DOUT(N__12140),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__12142),
            .PADOUT(N__12141),
            .PADIN(N__12140),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9336),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__12133),
            .DIN(N__12132),
            .DOUT(N__12131),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__12133),
            .PADOUT(N__12132),
            .PADIN(N__12131),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4719),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__12124),
            .DIN(N__12123),
            .DOUT(N__12122),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__12124),
            .PADOUT(N__12123),
            .PADIN(N__12122),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10323),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2950 (
            .O(N__12105),
            .I(N__12099));
    InMux I__2949 (
            .O(N__12104),
            .I(N__12096));
    InMux I__2948 (
            .O(N__12103),
            .I(N__12091));
    InMux I__2947 (
            .O(N__12102),
            .I(N__12091));
    LocalMux I__2946 (
            .O(N__12099),
            .I(N__12088));
    LocalMux I__2945 (
            .O(N__12096),
            .I(N__12083));
    LocalMux I__2944 (
            .O(N__12091),
            .I(N__12083));
    Span4Mux_v I__2943 (
            .O(N__12088),
            .I(N__12078));
    Span4Mux_v I__2942 (
            .O(N__12083),
            .I(N__12078));
    Span4Mux_v I__2941 (
            .O(N__12078),
            .I(N__12075));
    Sp12to4 I__2940 (
            .O(N__12075),
            .I(N__12072));
    Odrv12 I__2939 (
            .O(N__12072),
            .I(DRA_c_4));
    InMux I__2938 (
            .O(N__12069),
            .I(N__12066));
    LocalMux I__2937 (
            .O(N__12066),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__2936 (
            .O(N__12063),
            .I(N__12060));
    LocalMux I__2935 (
            .O(N__12060),
            .I(N__12057));
    Span4Mux_h I__2934 (
            .O(N__12057),
            .I(N__12054));
    Odrv4 I__2933 (
            .O(N__12054),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__2932 (
            .O(N__12051),
            .I(N__12048));
    LocalMux I__2931 (
            .O(N__12048),
            .I(N__12045));
    Odrv12 I__2930 (
            .O(N__12045),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_2 ));
    InMux I__2929 (
            .O(N__12042),
            .I(N__12039));
    LocalMux I__2928 (
            .O(N__12039),
            .I(N__12036));
    Span4Mux_v I__2927 (
            .O(N__12036),
            .I(N__12032));
    InMux I__2926 (
            .O(N__12035),
            .I(N__12029));
    Span4Mux_h I__2925 (
            .O(N__12032),
            .I(N__12026));
    LocalMux I__2924 (
            .O(N__12029),
            .I(N__12023));
    Odrv4 I__2923 (
            .O(N__12026),
            .I(RAS0n_c));
    Odrv12 I__2922 (
            .O(N__12023),
            .I(RAS0n_c));
    InMux I__2921 (
            .O(N__12018),
            .I(N__12015));
    LocalMux I__2920 (
            .O(N__12015),
            .I(N__12012));
    Span12Mux_v I__2919 (
            .O(N__12012),
            .I(N__12009));
    Odrv12 I__2918 (
            .O(N__12009),
            .I(RAS1n_c));
    CascadeMux I__2917 (
            .O(N__12006),
            .I(N__11996));
    InMux I__2916 (
            .O(N__12005),
            .I(N__11977));
    InMux I__2915 (
            .O(N__12004),
            .I(N__11977));
    InMux I__2914 (
            .O(N__12003),
            .I(N__11977));
    InMux I__2913 (
            .O(N__12002),
            .I(N__11977));
    InMux I__2912 (
            .O(N__12001),
            .I(N__11970));
    InMux I__2911 (
            .O(N__12000),
            .I(N__11965));
    InMux I__2910 (
            .O(N__11999),
            .I(N__11965));
    InMux I__2909 (
            .O(N__11996),
            .I(N__11960));
    InMux I__2908 (
            .O(N__11995),
            .I(N__11960));
    InMux I__2907 (
            .O(N__11994),
            .I(N__11953));
    InMux I__2906 (
            .O(N__11993),
            .I(N__11953));
    InMux I__2905 (
            .O(N__11992),
            .I(N__11953));
    InMux I__2904 (
            .O(N__11991),
            .I(N__11950));
    InMux I__2903 (
            .O(N__11990),
            .I(N__11943));
    InMux I__2902 (
            .O(N__11989),
            .I(N__11943));
    InMux I__2901 (
            .O(N__11988),
            .I(N__11943));
    InMux I__2900 (
            .O(N__11987),
            .I(N__11938));
    InMux I__2899 (
            .O(N__11986),
            .I(N__11938));
    LocalMux I__2898 (
            .O(N__11977),
            .I(N__11935));
    InMux I__2897 (
            .O(N__11976),
            .I(N__11932));
    InMux I__2896 (
            .O(N__11975),
            .I(N__11927));
    CascadeMux I__2895 (
            .O(N__11974),
            .I(N__11916));
    CascadeMux I__2894 (
            .O(N__11973),
            .I(N__11913));
    LocalMux I__2893 (
            .O(N__11970),
            .I(N__11906));
    LocalMux I__2892 (
            .O(N__11965),
            .I(N__11906));
    LocalMux I__2891 (
            .O(N__11960),
            .I(N__11903));
    LocalMux I__2890 (
            .O(N__11953),
            .I(N__11894));
    LocalMux I__2889 (
            .O(N__11950),
            .I(N__11894));
    LocalMux I__2888 (
            .O(N__11943),
            .I(N__11894));
    LocalMux I__2887 (
            .O(N__11938),
            .I(N__11894));
    Span4Mux_v I__2886 (
            .O(N__11935),
            .I(N__11889));
    LocalMux I__2885 (
            .O(N__11932),
            .I(N__11889));
    InMux I__2884 (
            .O(N__11931),
            .I(N__11886));
    InMux I__2883 (
            .O(N__11930),
            .I(N__11883));
    LocalMux I__2882 (
            .O(N__11927),
            .I(N__11880));
    InMux I__2881 (
            .O(N__11926),
            .I(N__11873));
    InMux I__2880 (
            .O(N__11925),
            .I(N__11873));
    InMux I__2879 (
            .O(N__11924),
            .I(N__11873));
    InMux I__2878 (
            .O(N__11923),
            .I(N__11870));
    InMux I__2877 (
            .O(N__11922),
            .I(N__11865));
    InMux I__2876 (
            .O(N__11921),
            .I(N__11865));
    InMux I__2875 (
            .O(N__11920),
            .I(N__11862));
    InMux I__2874 (
            .O(N__11919),
            .I(N__11853));
    InMux I__2873 (
            .O(N__11916),
            .I(N__11853));
    InMux I__2872 (
            .O(N__11913),
            .I(N__11853));
    InMux I__2871 (
            .O(N__11912),
            .I(N__11853));
    InMux I__2870 (
            .O(N__11911),
            .I(N__11850));
    Span4Mux_v I__2869 (
            .O(N__11906),
            .I(N__11847));
    Span4Mux_v I__2868 (
            .O(N__11903),
            .I(N__11835));
    Span4Mux_v I__2867 (
            .O(N__11894),
            .I(N__11835));
    Span4Mux_h I__2866 (
            .O(N__11889),
            .I(N__11835));
    LocalMux I__2865 (
            .O(N__11886),
            .I(N__11835));
    LocalMux I__2864 (
            .O(N__11883),
            .I(N__11835));
    Span12Mux_v I__2863 (
            .O(N__11880),
            .I(N__11829));
    LocalMux I__2862 (
            .O(N__11873),
            .I(N__11820));
    LocalMux I__2861 (
            .O(N__11870),
            .I(N__11820));
    LocalMux I__2860 (
            .O(N__11865),
            .I(N__11820));
    LocalMux I__2859 (
            .O(N__11862),
            .I(N__11820));
    LocalMux I__2858 (
            .O(N__11853),
            .I(N__11815));
    LocalMux I__2857 (
            .O(N__11850),
            .I(N__11815));
    Span4Mux_v I__2856 (
            .O(N__11847),
            .I(N__11812));
    InMux I__2855 (
            .O(N__11846),
            .I(N__11809));
    Span4Mux_v I__2854 (
            .O(N__11835),
            .I(N__11806));
    InMux I__2853 (
            .O(N__11834),
            .I(N__11803));
    InMux I__2852 (
            .O(N__11833),
            .I(N__11798));
    InMux I__2851 (
            .O(N__11832),
            .I(N__11798));
    Span12Mux_h I__2850 (
            .O(N__11829),
            .I(N__11795));
    Span12Mux_v I__2849 (
            .O(N__11820),
            .I(N__11792));
    Span12Mux_v I__2848 (
            .O(N__11815),
            .I(N__11789));
    Sp12to4 I__2847 (
            .O(N__11812),
            .I(N__11784));
    LocalMux I__2846 (
            .O(N__11809),
            .I(N__11784));
    Span4Mux_h I__2845 (
            .O(N__11806),
            .I(N__11781));
    LocalMux I__2844 (
            .O(N__11803),
            .I(N__11776));
    LocalMux I__2843 (
            .O(N__11798),
            .I(N__11776));
    Span12Mux_v I__2842 (
            .O(N__11795),
            .I(N__11771));
    Span12Mux_h I__2841 (
            .O(N__11792),
            .I(N__11771));
    Span12Mux_h I__2840 (
            .O(N__11789),
            .I(N__11768));
    Span12Mux_h I__2839 (
            .O(N__11784),
            .I(N__11761));
    Sp12to4 I__2838 (
            .O(N__11781),
            .I(N__11761));
    Span12Mux_v I__2837 (
            .O(N__11776),
            .I(N__11761));
    Odrv12 I__2836 (
            .O(N__11771),
            .I(RESETn_c));
    Odrv12 I__2835 (
            .O(N__11768),
            .I(RESETn_c));
    Odrv12 I__2834 (
            .O(N__11761),
            .I(RESETn_c));
    InMux I__2833 (
            .O(N__11754),
            .I(N__11751));
    LocalMux I__2832 (
            .O(N__11751),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ));
    InMux I__2831 (
            .O(N__11748),
            .I(N__11745));
    LocalMux I__2830 (
            .O(N__11745),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ));
    InMux I__2829 (
            .O(N__11742),
            .I(N__11739));
    LocalMux I__2828 (
            .O(N__11739),
            .I(N__11690));
    ClkMux I__2827 (
            .O(N__11738),
            .I(N__11592));
    ClkMux I__2826 (
            .O(N__11737),
            .I(N__11592));
    ClkMux I__2825 (
            .O(N__11736),
            .I(N__11592));
    ClkMux I__2824 (
            .O(N__11735),
            .I(N__11592));
    ClkMux I__2823 (
            .O(N__11734),
            .I(N__11592));
    ClkMux I__2822 (
            .O(N__11733),
            .I(N__11592));
    ClkMux I__2821 (
            .O(N__11732),
            .I(N__11592));
    ClkMux I__2820 (
            .O(N__11731),
            .I(N__11592));
    ClkMux I__2819 (
            .O(N__11730),
            .I(N__11592));
    ClkMux I__2818 (
            .O(N__11729),
            .I(N__11592));
    ClkMux I__2817 (
            .O(N__11728),
            .I(N__11592));
    ClkMux I__2816 (
            .O(N__11727),
            .I(N__11592));
    ClkMux I__2815 (
            .O(N__11726),
            .I(N__11592));
    ClkMux I__2814 (
            .O(N__11725),
            .I(N__11592));
    ClkMux I__2813 (
            .O(N__11724),
            .I(N__11592));
    ClkMux I__2812 (
            .O(N__11723),
            .I(N__11592));
    ClkMux I__2811 (
            .O(N__11722),
            .I(N__11592));
    ClkMux I__2810 (
            .O(N__11721),
            .I(N__11592));
    ClkMux I__2809 (
            .O(N__11720),
            .I(N__11592));
    ClkMux I__2808 (
            .O(N__11719),
            .I(N__11592));
    ClkMux I__2807 (
            .O(N__11718),
            .I(N__11592));
    ClkMux I__2806 (
            .O(N__11717),
            .I(N__11592));
    ClkMux I__2805 (
            .O(N__11716),
            .I(N__11592));
    ClkMux I__2804 (
            .O(N__11715),
            .I(N__11592));
    ClkMux I__2803 (
            .O(N__11714),
            .I(N__11592));
    ClkMux I__2802 (
            .O(N__11713),
            .I(N__11592));
    ClkMux I__2801 (
            .O(N__11712),
            .I(N__11592));
    ClkMux I__2800 (
            .O(N__11711),
            .I(N__11592));
    ClkMux I__2799 (
            .O(N__11710),
            .I(N__11592));
    ClkMux I__2798 (
            .O(N__11709),
            .I(N__11592));
    ClkMux I__2797 (
            .O(N__11708),
            .I(N__11592));
    ClkMux I__2796 (
            .O(N__11707),
            .I(N__11592));
    ClkMux I__2795 (
            .O(N__11706),
            .I(N__11592));
    ClkMux I__2794 (
            .O(N__11705),
            .I(N__11592));
    ClkMux I__2793 (
            .O(N__11704),
            .I(N__11592));
    ClkMux I__2792 (
            .O(N__11703),
            .I(N__11592));
    ClkMux I__2791 (
            .O(N__11702),
            .I(N__11592));
    ClkMux I__2790 (
            .O(N__11701),
            .I(N__11592));
    ClkMux I__2789 (
            .O(N__11700),
            .I(N__11592));
    ClkMux I__2788 (
            .O(N__11699),
            .I(N__11592));
    ClkMux I__2787 (
            .O(N__11698),
            .I(N__11592));
    ClkMux I__2786 (
            .O(N__11697),
            .I(N__11592));
    ClkMux I__2785 (
            .O(N__11696),
            .I(N__11592));
    ClkMux I__2784 (
            .O(N__11695),
            .I(N__11592));
    ClkMux I__2783 (
            .O(N__11694),
            .I(N__11592));
    ClkMux I__2782 (
            .O(N__11693),
            .I(N__11592));
    Glb2LocalMux I__2781 (
            .O(N__11690),
            .I(N__11592));
    ClkMux I__2780 (
            .O(N__11689),
            .I(N__11592));
    GlobalMux I__2779 (
            .O(N__11592),
            .I(CLK80_PLL));
    InMux I__2778 (
            .O(N__11589),
            .I(N__11586));
    LocalMux I__2777 (
            .O(N__11586),
            .I(N__11580));
    InMux I__2776 (
            .O(N__11585),
            .I(N__11577));
    InMux I__2775 (
            .O(N__11584),
            .I(N__11572));
    InMux I__2774 (
            .O(N__11583),
            .I(N__11572));
    Span4Mux_v I__2773 (
            .O(N__11580),
            .I(N__11569));
    LocalMux I__2772 (
            .O(N__11577),
            .I(N__11564));
    LocalMux I__2771 (
            .O(N__11572),
            .I(N__11564));
    Span4Mux_v I__2770 (
            .O(N__11569),
            .I(N__11561));
    Span12Mux_v I__2769 (
            .O(N__11564),
            .I(N__11558));
    Span4Mux_h I__2768 (
            .O(N__11561),
            .I(N__11555));
    Odrv12 I__2767 (
            .O(N__11558),
            .I(DRA_c_3));
    Odrv4 I__2766 (
            .O(N__11555),
            .I(DRA_c_3));
    InMux I__2765 (
            .O(N__11550),
            .I(N__11547));
    LocalMux I__2764 (
            .O(N__11547),
            .I(N__11544));
    Span4Mux_v I__2763 (
            .O(N__11544),
            .I(N__11538));
    InMux I__2762 (
            .O(N__11543),
            .I(N__11535));
    InMux I__2761 (
            .O(N__11542),
            .I(N__11530));
    InMux I__2760 (
            .O(N__11541),
            .I(N__11530));
    Span4Mux_v I__2759 (
            .O(N__11538),
            .I(N__11527));
    LocalMux I__2758 (
            .O(N__11535),
            .I(N__11522));
    LocalMux I__2757 (
            .O(N__11530),
            .I(N__11522));
    Span4Mux_h I__2756 (
            .O(N__11527),
            .I(N__11519));
    Span12Mux_v I__2755 (
            .O(N__11522),
            .I(N__11516));
    IoSpan4Mux I__2754 (
            .O(N__11519),
            .I(N__11513));
    Odrv12 I__2753 (
            .O(N__11516),
            .I(DRA_c_2));
    Odrv4 I__2752 (
            .O(N__11513),
            .I(DRA_c_2));
    InMux I__2751 (
            .O(N__11508),
            .I(N__11505));
    LocalMux I__2750 (
            .O(N__11505),
            .I(N__11502));
    Span12Mux_h I__2749 (
            .O(N__11502),
            .I(N__11499));
    Odrv12 I__2748 (
            .O(N__11499),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__2747 (
            .O(N__11496),
            .I(N__11490));
    InMux I__2746 (
            .O(N__11495),
            .I(N__11487));
    InMux I__2745 (
            .O(N__11494),
            .I(N__11484));
    InMux I__2744 (
            .O(N__11493),
            .I(N__11481));
    LocalMux I__2743 (
            .O(N__11490),
            .I(N__11474));
    LocalMux I__2742 (
            .O(N__11487),
            .I(N__11474));
    LocalMux I__2741 (
            .O(N__11484),
            .I(N__11474));
    LocalMux I__2740 (
            .O(N__11481),
            .I(N__11471));
    Span4Mux_v I__2739 (
            .O(N__11474),
            .I(N__11468));
    Span4Mux_v I__2738 (
            .O(N__11471),
            .I(N__11465));
    Span4Mux_v I__2737 (
            .O(N__11468),
            .I(N__11462));
    Span4Mux_h I__2736 (
            .O(N__11465),
            .I(N__11459));
    Sp12to4 I__2735 (
            .O(N__11462),
            .I(N__11456));
    IoSpan4Mux I__2734 (
            .O(N__11459),
            .I(N__11453));
    Odrv12 I__2733 (
            .O(N__11456),
            .I(DRA_c_5));
    Odrv4 I__2732 (
            .O(N__11453),
            .I(DRA_c_5));
    InMux I__2731 (
            .O(N__11448),
            .I(N__11444));
    InMux I__2730 (
            .O(N__11447),
            .I(N__11441));
    LocalMux I__2729 (
            .O(N__11444),
            .I(N__11434));
    LocalMux I__2728 (
            .O(N__11441),
            .I(N__11434));
    InMux I__2727 (
            .O(N__11440),
            .I(N__11431));
    InMux I__2726 (
            .O(N__11439),
            .I(N__11428));
    Span4Mux_h I__2725 (
            .O(N__11434),
            .I(N__11423));
    LocalMux I__2724 (
            .O(N__11431),
            .I(N__11423));
    LocalMux I__2723 (
            .O(N__11428),
            .I(N__11420));
    Span4Mux_h I__2722 (
            .O(N__11423),
            .I(N__11417));
    Span4Mux_v I__2721 (
            .O(N__11420),
            .I(N__11414));
    Span4Mux_v I__2720 (
            .O(N__11417),
            .I(N__11411));
    Sp12to4 I__2719 (
            .O(N__11414),
            .I(N__11408));
    Span4Mux_h I__2718 (
            .O(N__11411),
            .I(N__11405));
    Odrv12 I__2717 (
            .O(N__11408),
            .I(DRA_c_6));
    Odrv4 I__2716 (
            .O(N__11405),
            .I(DRA_c_6));
    InMux I__2715 (
            .O(N__11400),
            .I(N__11397));
    LocalMux I__2714 (
            .O(N__11397),
            .I(N__11390));
    CascadeMux I__2713 (
            .O(N__11396),
            .I(N__11387));
    InMux I__2712 (
            .O(N__11395),
            .I(N__11380));
    InMux I__2711 (
            .O(N__11394),
            .I(N__11370));
    InMux I__2710 (
            .O(N__11393),
            .I(N__11370));
    Span4Mux_v I__2709 (
            .O(N__11390),
            .I(N__11367));
    InMux I__2708 (
            .O(N__11387),
            .I(N__11360));
    InMux I__2707 (
            .O(N__11386),
            .I(N__11360));
    InMux I__2706 (
            .O(N__11385),
            .I(N__11360));
    CascadeMux I__2705 (
            .O(N__11384),
            .I(N__11357));
    CascadeMux I__2704 (
            .O(N__11383),
            .I(N__11353));
    LocalMux I__2703 (
            .O(N__11380),
            .I(N__11347));
    InMux I__2702 (
            .O(N__11379),
            .I(N__11344));
    InMux I__2701 (
            .O(N__11378),
            .I(N__11339));
    InMux I__2700 (
            .O(N__11377),
            .I(N__11339));
    InMux I__2699 (
            .O(N__11376),
            .I(N__11334));
    InMux I__2698 (
            .O(N__11375),
            .I(N__11334));
    LocalMux I__2697 (
            .O(N__11370),
            .I(N__11331));
    Span4Mux_h I__2696 (
            .O(N__11367),
            .I(N__11326));
    LocalMux I__2695 (
            .O(N__11360),
            .I(N__11326));
    InMux I__2694 (
            .O(N__11357),
            .I(N__11317));
    InMux I__2693 (
            .O(N__11356),
            .I(N__11317));
    InMux I__2692 (
            .O(N__11353),
            .I(N__11317));
    InMux I__2691 (
            .O(N__11352),
            .I(N__11317));
    InMux I__2690 (
            .O(N__11351),
            .I(N__11314));
    InMux I__2689 (
            .O(N__11350),
            .I(N__11311));
    Span4Mux_v I__2688 (
            .O(N__11347),
            .I(N__11308));
    LocalMux I__2687 (
            .O(N__11344),
            .I(N__11305));
    LocalMux I__2686 (
            .O(N__11339),
            .I(N__11299));
    LocalMux I__2685 (
            .O(N__11334),
            .I(N__11299));
    Span4Mux_h I__2684 (
            .O(N__11331),
            .I(N__11286));
    Span4Mux_v I__2683 (
            .O(N__11326),
            .I(N__11286));
    LocalMux I__2682 (
            .O(N__11317),
            .I(N__11286));
    LocalMux I__2681 (
            .O(N__11314),
            .I(N__11286));
    LocalMux I__2680 (
            .O(N__11311),
            .I(N__11286));
    Span4Mux_h I__2679 (
            .O(N__11308),
            .I(N__11281));
    Span4Mux_v I__2678 (
            .O(N__11305),
            .I(N__11281));
    InMux I__2677 (
            .O(N__11304),
            .I(N__11278));
    Span4Mux_v I__2676 (
            .O(N__11299),
            .I(N__11275));
    InMux I__2675 (
            .O(N__11298),
            .I(N__11272));
    InMux I__2674 (
            .O(N__11297),
            .I(N__11269));
    Span4Mux_h I__2673 (
            .O(N__11286),
            .I(N__11266));
    Sp12to4 I__2672 (
            .O(N__11281),
            .I(N__11263));
    LocalMux I__2671 (
            .O(N__11278),
            .I(N__11254));
    Sp12to4 I__2670 (
            .O(N__11275),
            .I(N__11254));
    LocalMux I__2669 (
            .O(N__11272),
            .I(N__11254));
    LocalMux I__2668 (
            .O(N__11269),
            .I(N__11254));
    Span4Mux_h I__2667 (
            .O(N__11266),
            .I(N__11251));
    Span12Mux_h I__2666 (
            .O(N__11263),
            .I(N__11248));
    Span12Mux_h I__2665 (
            .O(N__11254),
            .I(N__11243));
    Sp12to4 I__2664 (
            .O(N__11251),
            .I(N__11243));
    Span12Mux_v I__2663 (
            .O(N__11248),
            .I(N__11240));
    Span12Mux_v I__2662 (
            .O(N__11243),
            .I(N__11237));
    Odrv12 I__2661 (
            .O(N__11240),
            .I(AGNUS_REV_c));
    Odrv12 I__2660 (
            .O(N__11237),
            .I(AGNUS_REV_c));
    InMux I__2659 (
            .O(N__11232),
            .I(N__11228));
    InMux I__2658 (
            .O(N__11231),
            .I(N__11225));
    LocalMux I__2657 (
            .O(N__11228),
            .I(N__11222));
    LocalMux I__2656 (
            .O(N__11225),
            .I(N__11219));
    Span4Mux_h I__2655 (
            .O(N__11222),
            .I(N__11216));
    Span4Mux_h I__2654 (
            .O(N__11219),
            .I(N__11213));
    Odrv4 I__2653 (
            .O(N__11216),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    Odrv4 I__2652 (
            .O(N__11213),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    ClkMux I__2651 (
            .O(N__11208),
            .I(N__11190));
    ClkMux I__2650 (
            .O(N__11207),
            .I(N__11190));
    ClkMux I__2649 (
            .O(N__11206),
            .I(N__11190));
    ClkMux I__2648 (
            .O(N__11205),
            .I(N__11190));
    ClkMux I__2647 (
            .O(N__11204),
            .I(N__11190));
    ClkMux I__2646 (
            .O(N__11203),
            .I(N__11190));
    GlobalMux I__2645 (
            .O(N__11190),
            .I(N__11187));
    gio2CtrlBuf I__2644 (
            .O(N__11187),
            .I(C3_c_g));
    CEMux I__2643 (
            .O(N__11184),
            .I(N__11151));
    CEMux I__2642 (
            .O(N__11183),
            .I(N__11151));
    CEMux I__2641 (
            .O(N__11182),
            .I(N__11151));
    CEMux I__2640 (
            .O(N__11181),
            .I(N__11151));
    CEMux I__2639 (
            .O(N__11180),
            .I(N__11151));
    CEMux I__2638 (
            .O(N__11179),
            .I(N__11151));
    CEMux I__2637 (
            .O(N__11178),
            .I(N__11151));
    CEMux I__2636 (
            .O(N__11177),
            .I(N__11151));
    CEMux I__2635 (
            .O(N__11176),
            .I(N__11151));
    CEMux I__2634 (
            .O(N__11175),
            .I(N__11151));
    CEMux I__2633 (
            .O(N__11174),
            .I(N__11151));
    GlobalMux I__2632 (
            .O(N__11151),
            .I(N__11148));
    gio2CtrlBuf I__2631 (
            .O(N__11148),
            .I(DBRn_c_i_0_g));
    InMux I__2630 (
            .O(N__11145),
            .I(N__11136));
    InMux I__2629 (
            .O(N__11144),
            .I(N__11131));
    InMux I__2628 (
            .O(N__11143),
            .I(N__11131));
    InMux I__2627 (
            .O(N__11142),
            .I(N__11128));
    InMux I__2626 (
            .O(N__11141),
            .I(N__11125));
    InMux I__2625 (
            .O(N__11140),
            .I(N__11122));
    InMux I__2624 (
            .O(N__11139),
            .I(N__11119));
    LocalMux I__2623 (
            .O(N__11136),
            .I(N__11099));
    LocalMux I__2622 (
            .O(N__11131),
            .I(N__11093));
    LocalMux I__2621 (
            .O(N__11128),
            .I(N__11089));
    LocalMux I__2620 (
            .O(N__11125),
            .I(N__11086));
    LocalMux I__2619 (
            .O(N__11122),
            .I(N__11070));
    LocalMux I__2618 (
            .O(N__11119),
            .I(N__11064));
    SRMux I__2617 (
            .O(N__11118),
            .I(N__10971));
    SRMux I__2616 (
            .O(N__11117),
            .I(N__10971));
    SRMux I__2615 (
            .O(N__11116),
            .I(N__10971));
    SRMux I__2614 (
            .O(N__11115),
            .I(N__10971));
    SRMux I__2613 (
            .O(N__11114),
            .I(N__10971));
    SRMux I__2612 (
            .O(N__11113),
            .I(N__10971));
    SRMux I__2611 (
            .O(N__11112),
            .I(N__10971));
    SRMux I__2610 (
            .O(N__11111),
            .I(N__10971));
    SRMux I__2609 (
            .O(N__11110),
            .I(N__10971));
    SRMux I__2608 (
            .O(N__11109),
            .I(N__10971));
    SRMux I__2607 (
            .O(N__11108),
            .I(N__10971));
    SRMux I__2606 (
            .O(N__11107),
            .I(N__10971));
    SRMux I__2605 (
            .O(N__11106),
            .I(N__10971));
    SRMux I__2604 (
            .O(N__11105),
            .I(N__10971));
    SRMux I__2603 (
            .O(N__11104),
            .I(N__10971));
    SRMux I__2602 (
            .O(N__11103),
            .I(N__10971));
    SRMux I__2601 (
            .O(N__11102),
            .I(N__10971));
    Glb2LocalMux I__2600 (
            .O(N__11099),
            .I(N__10971));
    SRMux I__2599 (
            .O(N__11098),
            .I(N__10971));
    SRMux I__2598 (
            .O(N__11097),
            .I(N__10971));
    SRMux I__2597 (
            .O(N__11096),
            .I(N__10971));
    Glb2LocalMux I__2596 (
            .O(N__11093),
            .I(N__10971));
    SRMux I__2595 (
            .O(N__11092),
            .I(N__10971));
    Glb2LocalMux I__2594 (
            .O(N__11089),
            .I(N__10971));
    Glb2LocalMux I__2593 (
            .O(N__11086),
            .I(N__10971));
    SRMux I__2592 (
            .O(N__11085),
            .I(N__10971));
    SRMux I__2591 (
            .O(N__11084),
            .I(N__10971));
    SRMux I__2590 (
            .O(N__11083),
            .I(N__10971));
    SRMux I__2589 (
            .O(N__11082),
            .I(N__10971));
    SRMux I__2588 (
            .O(N__11081),
            .I(N__10971));
    SRMux I__2587 (
            .O(N__11080),
            .I(N__10971));
    SRMux I__2586 (
            .O(N__11079),
            .I(N__10971));
    SRMux I__2585 (
            .O(N__11078),
            .I(N__10971));
    SRMux I__2584 (
            .O(N__11077),
            .I(N__10971));
    SRMux I__2583 (
            .O(N__11076),
            .I(N__10971));
    SRMux I__2582 (
            .O(N__11075),
            .I(N__10971));
    SRMux I__2581 (
            .O(N__11074),
            .I(N__10971));
    SRMux I__2580 (
            .O(N__11073),
            .I(N__10971));
    Glb2LocalMux I__2579 (
            .O(N__11070),
            .I(N__10971));
    SRMux I__2578 (
            .O(N__11069),
            .I(N__10971));
    SRMux I__2577 (
            .O(N__11068),
            .I(N__10971));
    SRMux I__2576 (
            .O(N__11067),
            .I(N__10971));
    Glb2LocalMux I__2575 (
            .O(N__11064),
            .I(N__10971));
    SRMux I__2574 (
            .O(N__11063),
            .I(N__10971));
    SRMux I__2573 (
            .O(N__11062),
            .I(N__10971));
    GlobalMux I__2572 (
            .O(N__10971),
            .I(N__10968));
    gio2CtrlBuf I__2571 (
            .O(N__10968),
            .I(RESETn_c_i_g));
    InMux I__2570 (
            .O(N__10965),
            .I(N__10960));
    InMux I__2569 (
            .O(N__10964),
            .I(N__10956));
    InMux I__2568 (
            .O(N__10963),
            .I(N__10952));
    LocalMux I__2567 (
            .O(N__10960),
            .I(N__10949));
    InMux I__2566 (
            .O(N__10959),
            .I(N__10946));
    LocalMux I__2565 (
            .O(N__10956),
            .I(N__10943));
    InMux I__2564 (
            .O(N__10955),
            .I(N__10940));
    LocalMux I__2563 (
            .O(N__10952),
            .I(N__10935));
    Span4Mux_v I__2562 (
            .O(N__10949),
            .I(N__10935));
    LocalMux I__2561 (
            .O(N__10946),
            .I(N__10932));
    Span4Mux_v I__2560 (
            .O(N__10943),
            .I(N__10929));
    LocalMux I__2559 (
            .O(N__10940),
            .I(N__10926));
    Span4Mux_h I__2558 (
            .O(N__10935),
            .I(N__10923));
    Span4Mux_v I__2557 (
            .O(N__10932),
            .I(N__10920));
    Sp12to4 I__2556 (
            .O(N__10929),
            .I(N__10917));
    Sp12to4 I__2555 (
            .O(N__10926),
            .I(N__10914));
    Sp12to4 I__2554 (
            .O(N__10923),
            .I(N__10909));
    Sp12to4 I__2553 (
            .O(N__10920),
            .I(N__10909));
    Span12Mux_h I__2552 (
            .O(N__10917),
            .I(N__10904));
    Span12Mux_v I__2551 (
            .O(N__10914),
            .I(N__10904));
    Span12Mux_h I__2550 (
            .O(N__10909),
            .I(N__10901));
    Span12Mux_h I__2549 (
            .O(N__10904),
            .I(N__10896));
    Span12Mux_v I__2548 (
            .O(N__10901),
            .I(N__10896));
    Odrv12 I__2547 (
            .O(N__10896),
            .I(RnW_c));
    InMux I__2546 (
            .O(N__10893),
            .I(N__10890));
    LocalMux I__2545 (
            .O(N__10890),
            .I(N__10886));
    InMux I__2544 (
            .O(N__10889),
            .I(N__10883));
    Span4Mux_v I__2543 (
            .O(N__10886),
            .I(N__10878));
    LocalMux I__2542 (
            .O(N__10883),
            .I(N__10875));
    InMux I__2541 (
            .O(N__10882),
            .I(N__10870));
    InMux I__2540 (
            .O(N__10881),
            .I(N__10870));
    Span4Mux_v I__2539 (
            .O(N__10878),
            .I(N__10864));
    Span4Mux_v I__2538 (
            .O(N__10875),
            .I(N__10864));
    LocalMux I__2537 (
            .O(N__10870),
            .I(N__10861));
    InMux I__2536 (
            .O(N__10869),
            .I(N__10858));
    Span4Mux_h I__2535 (
            .O(N__10864),
            .I(N__10852));
    Span4Mux_h I__2534 (
            .O(N__10861),
            .I(N__10852));
    LocalMux I__2533 (
            .O(N__10858),
            .I(N__10849));
    InMux I__2532 (
            .O(N__10857),
            .I(N__10846));
    Sp12to4 I__2531 (
            .O(N__10852),
            .I(N__10843));
    Span12Mux_v I__2530 (
            .O(N__10849),
            .I(N__10840));
    LocalMux I__2529 (
            .O(N__10846),
            .I(N__10837));
    Span12Mux_v I__2528 (
            .O(N__10843),
            .I(N__10834));
    Span12Mux_h I__2527 (
            .O(N__10840),
            .I(N__10831));
    Span4Mux_v I__2526 (
            .O(N__10837),
            .I(N__10828));
    Odrv12 I__2525 (
            .O(N__10834),
            .I(CASUn_c));
    Odrv12 I__2524 (
            .O(N__10831),
            .I(CASUn_c));
    Odrv4 I__2523 (
            .O(N__10828),
            .I(CASUn_c));
    CascadeMux I__2522 (
            .O(N__10821),
            .I(N__10818));
    InMux I__2521 (
            .O(N__10818),
            .I(N__10815));
    LocalMux I__2520 (
            .O(N__10815),
            .I(N__10811));
    InMux I__2519 (
            .O(N__10814),
            .I(N__10808));
    Span12Mux_s7_v I__2518 (
            .O(N__10811),
            .I(N__10804));
    LocalMux I__2517 (
            .O(N__10808),
            .I(N__10801));
    CascadeMux I__2516 (
            .O(N__10807),
            .I(N__10798));
    Span12Mux_v I__2515 (
            .O(N__10804),
            .I(N__10795));
    Span12Mux_v I__2514 (
            .O(N__10801),
            .I(N__10792));
    InMux I__2513 (
            .O(N__10798),
            .I(N__10789));
    Odrv12 I__2512 (
            .O(N__10795),
            .I(DMA_WRITE_CYCLE));
    Odrv12 I__2511 (
            .O(N__10792),
            .I(DMA_WRITE_CYCLE));
    LocalMux I__2510 (
            .O(N__10789),
            .I(DMA_WRITE_CYCLE));
    CascadeMux I__2509 (
            .O(N__10782),
            .I(N__10779));
    InMux I__2508 (
            .O(N__10779),
            .I(N__10772));
    InMux I__2507 (
            .O(N__10778),
            .I(N__10772));
    InMux I__2506 (
            .O(N__10777),
            .I(N__10767));
    LocalMux I__2505 (
            .O(N__10772),
            .I(N__10764));
    InMux I__2504 (
            .O(N__10771),
            .I(N__10759));
    InMux I__2503 (
            .O(N__10770),
            .I(N__10759));
    LocalMux I__2502 (
            .O(N__10767),
            .I(N__10756));
    Span4Mux_h I__2501 (
            .O(N__10764),
            .I(N__10753));
    LocalMux I__2500 (
            .O(N__10759),
            .I(N__10750));
    Span4Mux_h I__2499 (
            .O(N__10756),
            .I(N__10747));
    Sp12to4 I__2498 (
            .O(N__10753),
            .I(N__10743));
    Span12Mux_v I__2497 (
            .O(N__10750),
            .I(N__10740));
    Span4Mux_v I__2496 (
            .O(N__10747),
            .I(N__10737));
    InMux I__2495 (
            .O(N__10746),
            .I(N__10734));
    Span12Mux_v I__2494 (
            .O(N__10743),
            .I(N__10731));
    Span12Mux_h I__2493 (
            .O(N__10740),
            .I(N__10728));
    Sp12to4 I__2492 (
            .O(N__10737),
            .I(N__10725));
    LocalMux I__2491 (
            .O(N__10734),
            .I(N__10722));
    Span12Mux_h I__2490 (
            .O(N__10731),
            .I(N__10717));
    Span12Mux_v I__2489 (
            .O(N__10728),
            .I(N__10717));
    Span12Mux_h I__2488 (
            .O(N__10725),
            .I(N__10712));
    Span12Mux_v I__2487 (
            .O(N__10722),
            .I(N__10712));
    Odrv12 I__2486 (
            .O(N__10717),
            .I(CASLn_c));
    Odrv12 I__2485 (
            .O(N__10712),
            .I(CASLn_c));
    IoInMux I__2484 (
            .O(N__10707),
            .I(N__10704));
    LocalMux I__2483 (
            .O(N__10704),
            .I(N__10701));
    IoSpan4Mux I__2482 (
            .O(N__10701),
            .I(N__10698));
    IoSpan4Mux I__2481 (
            .O(N__10698),
            .I(N__10695));
    Span4Mux_s3_v I__2480 (
            .O(N__10695),
            .I(N__10692));
    Odrv4 I__2479 (
            .O(N__10692),
            .I(N_409));
    InMux I__2478 (
            .O(N__10689),
            .I(N__10686));
    LocalMux I__2477 (
            .O(N__10686),
            .I(N__10683));
    Odrv12 I__2476 (
            .O(N__10683),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__2475 (
            .O(N__10680),
            .I(N__10677));
    LocalMux I__2474 (
            .O(N__10677),
            .I(N__10674));
    Span4Mux_h I__2473 (
            .O(N__10674),
            .I(N__10671));
    Span4Mux_v I__2472 (
            .O(N__10671),
            .I(N__10668));
    Odrv4 I__2471 (
            .O(N__10668),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__2470 (
            .O(N__10665),
            .I(N__10662));
    LocalMux I__2469 (
            .O(N__10662),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__2468 (
            .O(N__10659),
            .I(N__10655));
    InMux I__2467 (
            .O(N__10658),
            .I(N__10650));
    LocalMux I__2466 (
            .O(N__10655),
            .I(N__10647));
    InMux I__2465 (
            .O(N__10654),
            .I(N__10644));
    InMux I__2464 (
            .O(N__10653),
            .I(N__10641));
    LocalMux I__2463 (
            .O(N__10650),
            .I(N__10638));
    Span4Mux_v I__2462 (
            .O(N__10647),
            .I(N__10631));
    LocalMux I__2461 (
            .O(N__10644),
            .I(N__10631));
    LocalMux I__2460 (
            .O(N__10641),
            .I(N__10631));
    Span12Mux_h I__2459 (
            .O(N__10638),
            .I(N__10628));
    Sp12to4 I__2458 (
            .O(N__10631),
            .I(N__10625));
    Span12Mux_v I__2457 (
            .O(N__10628),
            .I(N__10622));
    Span12Mux_v I__2456 (
            .O(N__10625),
            .I(N__10619));
    Odrv12 I__2455 (
            .O(N__10622),
            .I(DRA_c_1));
    Odrv12 I__2454 (
            .O(N__10619),
            .I(DRA_c_1));
    InMux I__2453 (
            .O(N__10614),
            .I(N__10611));
    LocalMux I__2452 (
            .O(N__10611),
            .I(N__10608));
    Odrv4 I__2451 (
            .O(N__10608),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__2450 (
            .O(N__10605),
            .I(N__10602));
    LocalMux I__2449 (
            .O(N__10602),
            .I(N__10596));
    InMux I__2448 (
            .O(N__10601),
            .I(N__10591));
    InMux I__2447 (
            .O(N__10600),
            .I(N__10591));
    InMux I__2446 (
            .O(N__10599),
            .I(N__10587));
    Span4Mux_v I__2445 (
            .O(N__10596),
            .I(N__10582));
    LocalMux I__2444 (
            .O(N__10591),
            .I(N__10582));
    InMux I__2443 (
            .O(N__10590),
            .I(N__10579));
    LocalMux I__2442 (
            .O(N__10587),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__2441 (
            .O(N__10582),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__2440 (
            .O(N__10579),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    IoInMux I__2439 (
            .O(N__10572),
            .I(N__10569));
    LocalMux I__2438 (
            .O(N__10569),
            .I(N__10566));
    IoSpan4Mux I__2437 (
            .O(N__10566),
            .I(N__10563));
    Sp12to4 I__2436 (
            .O(N__10563),
            .I(N__10560));
    Span12Mux_s9_v I__2435 (
            .O(N__10560),
            .I(N__10557));
    Odrv12 I__2434 (
            .O(N__10557),
            .I(WEn_c));
    InMux I__2433 (
            .O(N__10554),
            .I(N__10551));
    LocalMux I__2432 (
            .O(N__10551),
            .I(\U712_CHIP_RAM.CMA_5_i_0_9 ));
    InMux I__2431 (
            .O(N__10548),
            .I(N__10545));
    LocalMux I__2430 (
            .O(N__10545),
            .I(N__10542));
    Sp12to4 I__2429 (
            .O(N__10542),
            .I(N__10539));
    Span12Mux_v I__2428 (
            .O(N__10539),
            .I(N__10536));
    Span12Mux_h I__2427 (
            .O(N__10536),
            .I(N__10533));
    Odrv12 I__2426 (
            .O(N__10533),
            .I(A_c_19));
    CascadeMux I__2425 (
            .O(N__10530),
            .I(N__10525));
    InMux I__2424 (
            .O(N__10529),
            .I(N__10522));
    CascadeMux I__2423 (
            .O(N__10528),
            .I(N__10519));
    InMux I__2422 (
            .O(N__10525),
            .I(N__10511));
    LocalMux I__2421 (
            .O(N__10522),
            .I(N__10507));
    InMux I__2420 (
            .O(N__10519),
            .I(N__10504));
    CascadeMux I__2419 (
            .O(N__10518),
            .I(N__10501));
    CascadeMux I__2418 (
            .O(N__10517),
            .I(N__10495));
    InMux I__2417 (
            .O(N__10516),
            .I(N__10489));
    InMux I__2416 (
            .O(N__10515),
            .I(N__10489));
    InMux I__2415 (
            .O(N__10514),
            .I(N__10486));
    LocalMux I__2414 (
            .O(N__10511),
            .I(N__10480));
    InMux I__2413 (
            .O(N__10510),
            .I(N__10477));
    Span4Mux_h I__2412 (
            .O(N__10507),
            .I(N__10469));
    LocalMux I__2411 (
            .O(N__10504),
            .I(N__10469));
    InMux I__2410 (
            .O(N__10501),
            .I(N__10463));
    InMux I__2409 (
            .O(N__10500),
            .I(N__10460));
    InMux I__2408 (
            .O(N__10499),
            .I(N__10457));
    InMux I__2407 (
            .O(N__10498),
            .I(N__10454));
    InMux I__2406 (
            .O(N__10495),
            .I(N__10449));
    InMux I__2405 (
            .O(N__10494),
            .I(N__10449));
    LocalMux I__2404 (
            .O(N__10489),
            .I(N__10445));
    LocalMux I__2403 (
            .O(N__10486),
            .I(N__10442));
    CascadeMux I__2402 (
            .O(N__10485),
            .I(N__10439));
    InMux I__2401 (
            .O(N__10484),
            .I(N__10436));
    InMux I__2400 (
            .O(N__10483),
            .I(N__10432));
    Span4Mux_v I__2399 (
            .O(N__10480),
            .I(N__10429));
    LocalMux I__2398 (
            .O(N__10477),
            .I(N__10426));
    InMux I__2397 (
            .O(N__10476),
            .I(N__10423));
    InMux I__2396 (
            .O(N__10475),
            .I(N__10418));
    InMux I__2395 (
            .O(N__10474),
            .I(N__10418));
    Span4Mux_v I__2394 (
            .O(N__10469),
            .I(N__10415));
    InMux I__2393 (
            .O(N__10468),
            .I(N__10412));
    InMux I__2392 (
            .O(N__10467),
            .I(N__10407));
    InMux I__2391 (
            .O(N__10466),
            .I(N__10407));
    LocalMux I__2390 (
            .O(N__10463),
            .I(N__10402));
    LocalMux I__2389 (
            .O(N__10460),
            .I(N__10402));
    LocalMux I__2388 (
            .O(N__10457),
            .I(N__10399));
    LocalMux I__2387 (
            .O(N__10454),
            .I(N__10396));
    LocalMux I__2386 (
            .O(N__10449),
            .I(N__10393));
    InMux I__2385 (
            .O(N__10448),
            .I(N__10390));
    Span4Mux_v I__2384 (
            .O(N__10445),
            .I(N__10384));
    Span4Mux_v I__2383 (
            .O(N__10442),
            .I(N__10384));
    InMux I__2382 (
            .O(N__10439),
            .I(N__10381));
    LocalMux I__2381 (
            .O(N__10436),
            .I(N__10378));
    InMux I__2380 (
            .O(N__10435),
            .I(N__10375));
    LocalMux I__2379 (
            .O(N__10432),
            .I(N__10368));
    Span4Mux_h I__2378 (
            .O(N__10429),
            .I(N__10368));
    Span4Mux_v I__2377 (
            .O(N__10426),
            .I(N__10368));
    LocalMux I__2376 (
            .O(N__10423),
            .I(N__10359));
    LocalMux I__2375 (
            .O(N__10418),
            .I(N__10359));
    Sp12to4 I__2374 (
            .O(N__10415),
            .I(N__10359));
    LocalMux I__2373 (
            .O(N__10412),
            .I(N__10359));
    LocalMux I__2372 (
            .O(N__10407),
            .I(N__10354));
    Span12Mux_h I__2371 (
            .O(N__10402),
            .I(N__10354));
    Span4Mux_v I__2370 (
            .O(N__10399),
            .I(N__10345));
    Span4Mux_h I__2369 (
            .O(N__10396),
            .I(N__10345));
    Span4Mux_h I__2368 (
            .O(N__10393),
            .I(N__10345));
    LocalMux I__2367 (
            .O(N__10390),
            .I(N__10345));
    InMux I__2366 (
            .O(N__10389),
            .I(N__10342));
    Odrv4 I__2365 (
            .O(N__10384),
            .I(CPU_CYCLEm));
    LocalMux I__2364 (
            .O(N__10381),
            .I(CPU_CYCLEm));
    Odrv4 I__2363 (
            .O(N__10378),
            .I(CPU_CYCLEm));
    LocalMux I__2362 (
            .O(N__10375),
            .I(CPU_CYCLEm));
    Odrv4 I__2361 (
            .O(N__10368),
            .I(CPU_CYCLEm));
    Odrv12 I__2360 (
            .O(N__10359),
            .I(CPU_CYCLEm));
    Odrv12 I__2359 (
            .O(N__10354),
            .I(CPU_CYCLEm));
    Odrv4 I__2358 (
            .O(N__10345),
            .I(CPU_CYCLEm));
    LocalMux I__2357 (
            .O(N__10342),
            .I(CPU_CYCLEm));
    IoInMux I__2356 (
            .O(N__10323),
            .I(N__10320));
    LocalMux I__2355 (
            .O(N__10320),
            .I(N__10317));
    IoSpan4Mux I__2354 (
            .O(N__10317),
            .I(N__10314));
    Sp12to4 I__2353 (
            .O(N__10314),
            .I(N__10311));
    Span12Mux_s9_h I__2352 (
            .O(N__10311),
            .I(N__10308));
    Odrv12 I__2351 (
            .O(N__10308),
            .I(CMA_c_9));
    InMux I__2350 (
            .O(N__10305),
            .I(N__10302));
    LocalMux I__2349 (
            .O(N__10302),
            .I(N__10298));
    InMux I__2348 (
            .O(N__10301),
            .I(N__10295));
    Span4Mux_h I__2347 (
            .O(N__10298),
            .I(N__10286));
    LocalMux I__2346 (
            .O(N__10295),
            .I(N__10283));
    InMux I__2345 (
            .O(N__10294),
            .I(N__10276));
    InMux I__2344 (
            .O(N__10293),
            .I(N__10276));
    InMux I__2343 (
            .O(N__10292),
            .I(N__10276));
    InMux I__2342 (
            .O(N__10291),
            .I(N__10273));
    InMux I__2341 (
            .O(N__10290),
            .I(N__10270));
    InMux I__2340 (
            .O(N__10289),
            .I(N__10267));
    Span4Mux_h I__2339 (
            .O(N__10286),
            .I(N__10260));
    Span4Mux_h I__2338 (
            .O(N__10283),
            .I(N__10260));
    LocalMux I__2337 (
            .O(N__10276),
            .I(N__10257));
    LocalMux I__2336 (
            .O(N__10273),
            .I(N__10254));
    LocalMux I__2335 (
            .O(N__10270),
            .I(N__10249));
    LocalMux I__2334 (
            .O(N__10267),
            .I(N__10249));
    InMux I__2333 (
            .O(N__10266),
            .I(N__10246));
    InMux I__2332 (
            .O(N__10265),
            .I(N__10243));
    Odrv4 I__2331 (
            .O(N__10260),
            .I(\U712_CHIP_RAM.N_354 ));
    Odrv12 I__2330 (
            .O(N__10257),
            .I(\U712_CHIP_RAM.N_354 ));
    Odrv4 I__2329 (
            .O(N__10254),
            .I(\U712_CHIP_RAM.N_354 ));
    Odrv4 I__2328 (
            .O(N__10249),
            .I(\U712_CHIP_RAM.N_354 ));
    LocalMux I__2327 (
            .O(N__10246),
            .I(\U712_CHIP_RAM.N_354 ));
    LocalMux I__2326 (
            .O(N__10243),
            .I(\U712_CHIP_RAM.N_354 ));
    CascadeMux I__2325 (
            .O(N__10230),
            .I(N__10224));
    CascadeMux I__2324 (
            .O(N__10229),
            .I(N__10221));
    CascadeMux I__2323 (
            .O(N__10228),
            .I(N__10218));
    CascadeMux I__2322 (
            .O(N__10227),
            .I(N__10215));
    InMux I__2321 (
            .O(N__10224),
            .I(N__10212));
    InMux I__2320 (
            .O(N__10221),
            .I(N__10209));
    InMux I__2319 (
            .O(N__10218),
            .I(N__10204));
    InMux I__2318 (
            .O(N__10215),
            .I(N__10201));
    LocalMux I__2317 (
            .O(N__10212),
            .I(N__10198));
    LocalMux I__2316 (
            .O(N__10209),
            .I(N__10195));
    CascadeMux I__2315 (
            .O(N__10208),
            .I(N__10191));
    CascadeMux I__2314 (
            .O(N__10207),
            .I(N__10188));
    LocalMux I__2313 (
            .O(N__10204),
            .I(N__10185));
    LocalMux I__2312 (
            .O(N__10201),
            .I(N__10182));
    Span4Mux_v I__2311 (
            .O(N__10198),
            .I(N__10179));
    Span4Mux_v I__2310 (
            .O(N__10195),
            .I(N__10176));
    InMux I__2309 (
            .O(N__10194),
            .I(N__10173));
    InMux I__2308 (
            .O(N__10191),
            .I(N__10168));
    InMux I__2307 (
            .O(N__10188),
            .I(N__10168));
    Span4Mux_v I__2306 (
            .O(N__10185),
            .I(N__10165));
    Span12Mux_s11_v I__2305 (
            .O(N__10182),
            .I(N__10162));
    Span4Mux_h I__2304 (
            .O(N__10179),
            .I(N__10157));
    Span4Mux_h I__2303 (
            .O(N__10176),
            .I(N__10157));
    LocalMux I__2302 (
            .O(N__10173),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9 ));
    LocalMux I__2301 (
            .O(N__10168),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9 ));
    Odrv4 I__2300 (
            .O(N__10165),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9 ));
    Odrv12 I__2299 (
            .O(N__10162),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9 ));
    Odrv4 I__2298 (
            .O(N__10157),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9 ));
    InMux I__2297 (
            .O(N__10146),
            .I(N__10143));
    LocalMux I__2296 (
            .O(N__10143),
            .I(N__10140));
    Span4Mux_h I__2295 (
            .O(N__10140),
            .I(N__10137));
    Odrv4 I__2294 (
            .O(N__10137),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ));
    IoInMux I__2293 (
            .O(N__10134),
            .I(N__10131));
    LocalMux I__2292 (
            .O(N__10131),
            .I(N__10128));
    IoSpan4Mux I__2291 (
            .O(N__10128),
            .I(N__10125));
    IoSpan4Mux I__2290 (
            .O(N__10125),
            .I(N__10122));
    Sp12to4 I__2289 (
            .O(N__10122),
            .I(N__10119));
    Span12Mux_s9_h I__2288 (
            .O(N__10119),
            .I(N__10116));
    Odrv12 I__2287 (
            .O(N__10116),
            .I(CMA_c_4));
    CEMux I__2286 (
            .O(N__10113),
            .I(N__10109));
    CEMux I__2285 (
            .O(N__10112),
            .I(N__10105));
    LocalMux I__2284 (
            .O(N__10109),
            .I(N__10102));
    CEMux I__2283 (
            .O(N__10108),
            .I(N__10099));
    LocalMux I__2282 (
            .O(N__10105),
            .I(N__10093));
    Span4Mux_v I__2281 (
            .O(N__10102),
            .I(N__10088));
    LocalMux I__2280 (
            .O(N__10099),
            .I(N__10088));
    CEMux I__2279 (
            .O(N__10098),
            .I(N__10085));
    CEMux I__2278 (
            .O(N__10097),
            .I(N__10081));
    CEMux I__2277 (
            .O(N__10096),
            .I(N__10077));
    Span4Mux_h I__2276 (
            .O(N__10093),
            .I(N__10070));
    Span4Mux_h I__2275 (
            .O(N__10088),
            .I(N__10070));
    LocalMux I__2274 (
            .O(N__10085),
            .I(N__10070));
    CEMux I__2273 (
            .O(N__10084),
            .I(N__10067));
    LocalMux I__2272 (
            .O(N__10081),
            .I(N__10064));
    CEMux I__2271 (
            .O(N__10080),
            .I(N__10061));
    LocalMux I__2270 (
            .O(N__10077),
            .I(N__10058));
    Span4Mux_h I__2269 (
            .O(N__10070),
            .I(N__10053));
    LocalMux I__2268 (
            .O(N__10067),
            .I(N__10053));
    Span4Mux_h I__2267 (
            .O(N__10064),
            .I(N__10050));
    LocalMux I__2266 (
            .O(N__10061),
            .I(N__10047));
    Span4Mux_h I__2265 (
            .O(N__10058),
            .I(N__10042));
    Span4Mux_h I__2264 (
            .O(N__10053),
            .I(N__10042));
    Odrv4 I__2263 (
            .O(N__10050),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    Odrv4 I__2262 (
            .O(N__10047),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    Odrv4 I__2261 (
            .O(N__10042),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    CascadeMux I__2260 (
            .O(N__10035),
            .I(N__10031));
    InMux I__2259 (
            .O(N__10034),
            .I(N__10027));
    InMux I__2258 (
            .O(N__10031),
            .I(N__10023));
    InMux I__2257 (
            .O(N__10030),
            .I(N__10020));
    LocalMux I__2256 (
            .O(N__10027),
            .I(N__10017));
    InMux I__2255 (
            .O(N__10026),
            .I(N__10014));
    LocalMux I__2254 (
            .O(N__10023),
            .I(N__10011));
    LocalMux I__2253 (
            .O(N__10020),
            .I(N__10004));
    Span4Mux_h I__2252 (
            .O(N__10017),
            .I(N__10004));
    LocalMux I__2251 (
            .O(N__10014),
            .I(N__10004));
    Span4Mux_v I__2250 (
            .O(N__10011),
            .I(N__10001));
    Span4Mux_v I__2249 (
            .O(N__10004),
            .I(N__9998));
    Sp12to4 I__2248 (
            .O(N__10001),
            .I(N__9993));
    Sp12to4 I__2247 (
            .O(N__9998),
            .I(N__9993));
    Span12Mux_h I__2246 (
            .O(N__9993),
            .I(N__9990));
    Span12Mux_v I__2245 (
            .O(N__9990),
            .I(N__9987));
    Odrv12 I__2244 (
            .O(N__9987),
            .I(DRA_c_9));
    InMux I__2243 (
            .O(N__9984),
            .I(N__9981));
    LocalMux I__2242 (
            .O(N__9981),
            .I(N__9978));
    Odrv4 I__2241 (
            .O(N__9978),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    InMux I__2240 (
            .O(N__9975),
            .I(N__9972));
    LocalMux I__2239 (
            .O(N__9972),
            .I(N__9966));
    InMux I__2238 (
            .O(N__9971),
            .I(N__9963));
    InMux I__2237 (
            .O(N__9970),
            .I(N__9960));
    CascadeMux I__2236 (
            .O(N__9969),
            .I(N__9956));
    Span4Mux_v I__2235 (
            .O(N__9966),
            .I(N__9951));
    LocalMux I__2234 (
            .O(N__9963),
            .I(N__9951));
    LocalMux I__2233 (
            .O(N__9960),
            .I(N__9948));
    CascadeMux I__2232 (
            .O(N__9959),
            .I(N__9945));
    InMux I__2231 (
            .O(N__9956),
            .I(N__9942));
    Span4Mux_h I__2230 (
            .O(N__9951),
            .I(N__9939));
    Span4Mux_v I__2229 (
            .O(N__9948),
            .I(N__9936));
    InMux I__2228 (
            .O(N__9945),
            .I(N__9933));
    LocalMux I__2227 (
            .O(N__9942),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__2226 (
            .O(N__9939),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__2225 (
            .O(N__9936),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__2224 (
            .O(N__9933),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__2223 (
            .O(N__9924),
            .I(N__9921));
    LocalMux I__2222 (
            .O(N__9921),
            .I(N__9918));
    Span4Mux_s1_v I__2221 (
            .O(N__9918),
            .I(N__9915));
    Span4Mux_v I__2220 (
            .O(N__9915),
            .I(N__9912));
    Span4Mux_v I__2219 (
            .O(N__9912),
            .I(N__9909));
    Odrv4 I__2218 (
            .O(N__9909),
            .I(CMA_c_10));
    CascadeMux I__2217 (
            .O(N__9906),
            .I(N__9902));
    InMux I__2216 (
            .O(N__9905),
            .I(N__9899));
    InMux I__2215 (
            .O(N__9902),
            .I(N__9894));
    LocalMux I__2214 (
            .O(N__9899),
            .I(N__9890));
    InMux I__2213 (
            .O(N__9898),
            .I(N__9887));
    InMux I__2212 (
            .O(N__9897),
            .I(N__9884));
    LocalMux I__2211 (
            .O(N__9894),
            .I(N__9881));
    InMux I__2210 (
            .O(N__9893),
            .I(N__9877));
    Span4Mux_v I__2209 (
            .O(N__9890),
            .I(N__9870));
    LocalMux I__2208 (
            .O(N__9887),
            .I(N__9870));
    LocalMux I__2207 (
            .O(N__9884),
            .I(N__9870));
    Span4Mux_h I__2206 (
            .O(N__9881),
            .I(N__9867));
    InMux I__2205 (
            .O(N__9880),
            .I(N__9864));
    LocalMux I__2204 (
            .O(N__9877),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__2203 (
            .O(N__9870),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__2202 (
            .O(N__9867),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__2201 (
            .O(N__9864),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    CascadeMux I__2200 (
            .O(N__9855),
            .I(\U712_CHIP_RAM.N_354_cascade_ ));
    CascadeMux I__2199 (
            .O(N__9852),
            .I(N__9841));
    CascadeMux I__2198 (
            .O(N__9851),
            .I(N__9838));
    CascadeMux I__2197 (
            .O(N__9850),
            .I(N__9832));
    CascadeMux I__2196 (
            .O(N__9849),
            .I(N__9829));
    CascadeMux I__2195 (
            .O(N__9848),
            .I(N__9826));
    InMux I__2194 (
            .O(N__9847),
            .I(N__9817));
    InMux I__2193 (
            .O(N__9846),
            .I(N__9814));
    InMux I__2192 (
            .O(N__9845),
            .I(N__9809));
    InMux I__2191 (
            .O(N__9844),
            .I(N__9809));
    InMux I__2190 (
            .O(N__9841),
            .I(N__9805));
    InMux I__2189 (
            .O(N__9838),
            .I(N__9802));
    InMux I__2188 (
            .O(N__9837),
            .I(N__9799));
    InMux I__2187 (
            .O(N__9836),
            .I(N__9794));
    InMux I__2186 (
            .O(N__9835),
            .I(N__9794));
    InMux I__2185 (
            .O(N__9832),
            .I(N__9789));
    InMux I__2184 (
            .O(N__9829),
            .I(N__9789));
    InMux I__2183 (
            .O(N__9826),
            .I(N__9784));
    InMux I__2182 (
            .O(N__9825),
            .I(N__9784));
    InMux I__2181 (
            .O(N__9824),
            .I(N__9777));
    InMux I__2180 (
            .O(N__9823),
            .I(N__9777));
    InMux I__2179 (
            .O(N__9822),
            .I(N__9777));
    InMux I__2178 (
            .O(N__9821),
            .I(N__9774));
    InMux I__2177 (
            .O(N__9820),
            .I(N__9771));
    LocalMux I__2176 (
            .O(N__9817),
            .I(N__9761));
    LocalMux I__2175 (
            .O(N__9814),
            .I(N__9761));
    LocalMux I__2174 (
            .O(N__9809),
            .I(N__9761));
    InMux I__2173 (
            .O(N__9808),
            .I(N__9758));
    LocalMux I__2172 (
            .O(N__9805),
            .I(N__9755));
    LocalMux I__2171 (
            .O(N__9802),
            .I(N__9752));
    LocalMux I__2170 (
            .O(N__9799),
            .I(N__9749));
    LocalMux I__2169 (
            .O(N__9794),
            .I(N__9746));
    LocalMux I__2168 (
            .O(N__9789),
            .I(N__9739));
    LocalMux I__2167 (
            .O(N__9784),
            .I(N__9739));
    LocalMux I__2166 (
            .O(N__9777),
            .I(N__9739));
    LocalMux I__2165 (
            .O(N__9774),
            .I(N__9731));
    LocalMux I__2164 (
            .O(N__9771),
            .I(N__9731));
    InMux I__2163 (
            .O(N__9770),
            .I(N__9723));
    InMux I__2162 (
            .O(N__9769),
            .I(N__9723));
    InMux I__2161 (
            .O(N__9768),
            .I(N__9723));
    Span4Mux_v I__2160 (
            .O(N__9761),
            .I(N__9720));
    LocalMux I__2159 (
            .O(N__9758),
            .I(N__9707));
    Span4Mux_v I__2158 (
            .O(N__9755),
            .I(N__9707));
    Span4Mux_v I__2157 (
            .O(N__9752),
            .I(N__9707));
    Span4Mux_h I__2156 (
            .O(N__9749),
            .I(N__9707));
    Span4Mux_v I__2155 (
            .O(N__9746),
            .I(N__9707));
    Span4Mux_v I__2154 (
            .O(N__9739),
            .I(N__9707));
    InMux I__2153 (
            .O(N__9738),
            .I(N__9700));
    InMux I__2152 (
            .O(N__9737),
            .I(N__9700));
    InMux I__2151 (
            .O(N__9736),
            .I(N__9700));
    Span4Mux_v I__2150 (
            .O(N__9731),
            .I(N__9697));
    InMux I__2149 (
            .O(N__9730),
            .I(N__9694));
    LocalMux I__2148 (
            .O(N__9723),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2147 (
            .O(N__9720),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2146 (
            .O(N__9707),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2145 (
            .O(N__9700),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2144 (
            .O(N__9697),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2143 (
            .O(N__9694),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    InMux I__2142 (
            .O(N__9681),
            .I(N__9678));
    LocalMux I__2141 (
            .O(N__9678),
            .I(N__9675));
    Odrv4 I__2140 (
            .O(N__9675),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ));
    InMux I__2139 (
            .O(N__9672),
            .I(N__9669));
    LocalMux I__2138 (
            .O(N__9669),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ));
    InMux I__2137 (
            .O(N__9666),
            .I(N__9663));
    LocalMux I__2136 (
            .O(N__9663),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ));
    IoInMux I__2135 (
            .O(N__9660),
            .I(N__9657));
    LocalMux I__2134 (
            .O(N__9657),
            .I(N__9654));
    IoSpan4Mux I__2133 (
            .O(N__9654),
            .I(N__9651));
    Span4Mux_s2_h I__2132 (
            .O(N__9651),
            .I(N__9648));
    Sp12to4 I__2131 (
            .O(N__9648),
            .I(N__9645));
    Span12Mux_s10_h I__2130 (
            .O(N__9645),
            .I(N__9642));
    Odrv12 I__2129 (
            .O(N__9642),
            .I(CMA_c_5));
    InMux I__2128 (
            .O(N__9639),
            .I(N__9636));
    LocalMux I__2127 (
            .O(N__9636),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    IoInMux I__2126 (
            .O(N__9633),
            .I(N__9630));
    LocalMux I__2125 (
            .O(N__9630),
            .I(N__9627));
    Span4Mux_s1_h I__2124 (
            .O(N__9627),
            .I(N__9624));
    Sp12to4 I__2123 (
            .O(N__9624),
            .I(N__9621));
    Span12Mux_v I__2122 (
            .O(N__9621),
            .I(N__9618));
    Odrv12 I__2121 (
            .O(N__9618),
            .I(CMA_c_3));
    InMux I__2120 (
            .O(N__9615),
            .I(N__9612));
    LocalMux I__2119 (
            .O(N__9612),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__2118 (
            .O(N__9609),
            .I(N__9606));
    LocalMux I__2117 (
            .O(N__9606),
            .I(N__9603));
    Odrv12 I__2116 (
            .O(N__9603),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__2115 (
            .O(N__9600),
            .I(N__9597));
    LocalMux I__2114 (
            .O(N__9597),
            .I(N__9594));
    Span4Mux_h I__2113 (
            .O(N__9594),
            .I(N__9591));
    Odrv4 I__2112 (
            .O(N__9591),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__2111 (
            .O(N__9588),
            .I(N__9585));
    LocalMux I__2110 (
            .O(N__9585),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__2109 (
            .O(N__9582),
            .I(N__9579));
    LocalMux I__2108 (
            .O(N__9579),
            .I(N__9576));
    Odrv4 I__2107 (
            .O(N__9576),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__2106 (
            .O(N__9573),
            .I(N__9570));
    LocalMux I__2105 (
            .O(N__9570),
            .I(N__9567));
    Span4Mux_h I__2104 (
            .O(N__9567),
            .I(N__9564));
    Span4Mux_v I__2103 (
            .O(N__9564),
            .I(N__9561));
    Odrv4 I__2102 (
            .O(N__9561),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__2101 (
            .O(N__9558),
            .I(N__9552));
    InMux I__2100 (
            .O(N__9557),
            .I(N__9552));
    LocalMux I__2099 (
            .O(N__9552),
            .I(N__9549));
    Span4Mux_v I__2098 (
            .O(N__9549),
            .I(N__9544));
    InMux I__2097 (
            .O(N__9548),
            .I(N__9539));
    InMux I__2096 (
            .O(N__9547),
            .I(N__9539));
    Sp12to4 I__2095 (
            .O(N__9544),
            .I(N__9534));
    LocalMux I__2094 (
            .O(N__9539),
            .I(N__9534));
    Span12Mux_h I__2093 (
            .O(N__9534),
            .I(N__9531));
    Odrv12 I__2092 (
            .O(N__9531),
            .I(DRA_c_7));
    InMux I__2091 (
            .O(N__9528),
            .I(N__9523));
    InMux I__2090 (
            .O(N__9527),
            .I(N__9520));
    InMux I__2089 (
            .O(N__9526),
            .I(N__9517));
    LocalMux I__2088 (
            .O(N__9523),
            .I(N__9509));
    LocalMux I__2087 (
            .O(N__9520),
            .I(N__9509));
    LocalMux I__2086 (
            .O(N__9517),
            .I(N__9509));
    InMux I__2085 (
            .O(N__9516),
            .I(N__9506));
    Span4Mux_v I__2084 (
            .O(N__9509),
            .I(N__9503));
    LocalMux I__2083 (
            .O(N__9506),
            .I(N__9500));
    Sp12to4 I__2082 (
            .O(N__9503),
            .I(N__9497));
    Span12Mux_h I__2081 (
            .O(N__9500),
            .I(N__9494));
    Odrv12 I__2080 (
            .O(N__9497),
            .I(DRA_c_8));
    Odrv12 I__2079 (
            .O(N__9494),
            .I(DRA_c_8));
    CascadeMux I__2078 (
            .O(N__9489),
            .I(N__9486));
    InMux I__2077 (
            .O(N__9486),
            .I(N__9483));
    LocalMux I__2076 (
            .O(N__9483),
            .I(N__9480));
    Span12Mux_v I__2075 (
            .O(N__9480),
            .I(N__9477));
    Odrv12 I__2074 (
            .O(N__9477),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    CascadeMux I__2073 (
            .O(N__9474),
            .I(N__9470));
    InMux I__2072 (
            .O(N__9473),
            .I(N__9467));
    InMux I__2071 (
            .O(N__9470),
            .I(N__9464));
    LocalMux I__2070 (
            .O(N__9467),
            .I(N__9461));
    LocalMux I__2069 (
            .O(N__9464),
            .I(N__9456));
    Span4Mux_v I__2068 (
            .O(N__9461),
            .I(N__9456));
    Sp12to4 I__2067 (
            .O(N__9456),
            .I(N__9453));
    Span12Mux_h I__2066 (
            .O(N__9453),
            .I(N__9450));
    Span12Mux_v I__2065 (
            .O(N__9450),
            .I(N__9447));
    Odrv12 I__2064 (
            .O(N__9447),
            .I(DRA_c_0));
    InMux I__2063 (
            .O(N__9444),
            .I(N__9441));
    LocalMux I__2062 (
            .O(N__9441),
            .I(N__9438));
    Span4Mux_h I__2061 (
            .O(N__9438),
            .I(N__9435));
    Odrv4 I__2060 (
            .O(N__9435),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    IoInMux I__2059 (
            .O(N__9432),
            .I(N__9429));
    LocalMux I__2058 (
            .O(N__9429),
            .I(N__9426));
    Span4Mux_s3_v I__2057 (
            .O(N__9426),
            .I(N__9423));
    Span4Mux_v I__2056 (
            .O(N__9423),
            .I(N__9420));
    Odrv4 I__2055 (
            .O(N__9420),
            .I(RASn_c));
    IoInMux I__2054 (
            .O(N__9417),
            .I(N__9414));
    LocalMux I__2053 (
            .O(N__9414),
            .I(N__9411));
    IoSpan4Mux I__2052 (
            .O(N__9411),
            .I(N__9408));
    Span4Mux_s3_v I__2051 (
            .O(N__9408),
            .I(N__9405));
    Span4Mux_v I__2050 (
            .O(N__9405),
            .I(N__9402));
    Odrv4 I__2049 (
            .O(N__9402),
            .I(CRCSn_c));
    IoInMux I__2048 (
            .O(N__9399),
            .I(N__9396));
    LocalMux I__2047 (
            .O(N__9396),
            .I(N__9393));
    Span4Mux_s1_v I__2046 (
            .O(N__9393),
            .I(N__9390));
    Sp12to4 I__2045 (
            .O(N__9390),
            .I(N__9387));
    Span12Mux_s10_h I__2044 (
            .O(N__9387),
            .I(N__9384));
    Odrv12 I__2043 (
            .O(N__9384),
            .I(CASn_c));
    InMux I__2042 (
            .O(N__9381),
            .I(N__9376));
    CascadeMux I__2041 (
            .O(N__9380),
            .I(N__9373));
    InMux I__2040 (
            .O(N__9379),
            .I(N__9370));
    LocalMux I__2039 (
            .O(N__9376),
            .I(N__9367));
    InMux I__2038 (
            .O(N__9373),
            .I(N__9364));
    LocalMux I__2037 (
            .O(N__9370),
            .I(N__9361));
    Span4Mux_v I__2036 (
            .O(N__9367),
            .I(N__9357));
    LocalMux I__2035 (
            .O(N__9364),
            .I(N__9354));
    Span4Mux_h I__2034 (
            .O(N__9361),
            .I(N__9351));
    InMux I__2033 (
            .O(N__9360),
            .I(N__9348));
    Span4Mux_v I__2032 (
            .O(N__9357),
            .I(N__9343));
    Span4Mux_h I__2031 (
            .O(N__9354),
            .I(N__9343));
    Odrv4 I__2030 (
            .O(N__9351),
            .I(REG_CYCLEm));
    LocalMux I__2029 (
            .O(N__9348),
            .I(REG_CYCLEm));
    Odrv4 I__2028 (
            .O(N__9343),
            .I(REG_CYCLEm));
    IoInMux I__2027 (
            .O(N__9336),
            .I(N__9333));
    LocalMux I__2026 (
            .O(N__9333),
            .I(N__9330));
    Span4Mux_s1_v I__2025 (
            .O(N__9330),
            .I(N__9327));
    Span4Mux_v I__2024 (
            .O(N__9327),
            .I(N__9324));
    Sp12to4 I__2023 (
            .O(N__9324),
            .I(N__9321));
    Span12Mux_h I__2022 (
            .O(N__9321),
            .I(N__9318));
    Span12Mux_v I__2021 (
            .O(N__9318),
            .I(N__9315));
    Odrv12 I__2020 (
            .O(N__9315),
            .I(N_207_i));
    InMux I__2019 (
            .O(N__9312),
            .I(N__9309));
    LocalMux I__2018 (
            .O(N__9309),
            .I(N__9306));
    Odrv4 I__2017 (
            .O(N__9306),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    InMux I__2016 (
            .O(N__9303),
            .I(N__9300));
    LocalMux I__2015 (
            .O(N__9300),
            .I(N__9297));
    Span4Mux_v I__2014 (
            .O(N__9297),
            .I(N__9294));
    Span4Mux_v I__2013 (
            .O(N__9294),
            .I(N__9291));
    Span4Mux_v I__2012 (
            .O(N__9291),
            .I(N__9288));
    Sp12to4 I__2011 (
            .O(N__9288),
            .I(N__9285));
    Span12Mux_h I__2010 (
            .O(N__9285),
            .I(N__9282));
    Odrv12 I__2009 (
            .O(N__9282),
            .I(A_c_14));
    CascadeMux I__2008 (
            .O(N__9279),
            .I(N__9276));
    InMux I__2007 (
            .O(N__9276),
            .I(N__9273));
    LocalMux I__2006 (
            .O(N__9273),
            .I(N__9270));
    Odrv4 I__2005 (
            .O(N__9270),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ));
    InMux I__2004 (
            .O(N__9267),
            .I(N__9264));
    LocalMux I__2003 (
            .O(N__9264),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ));
    InMux I__2002 (
            .O(N__9261),
            .I(N__9258));
    LocalMux I__2001 (
            .O(N__9258),
            .I(N__9255));
    Span4Mux_h I__2000 (
            .O(N__9255),
            .I(N__9252));
    Span4Mux_v I__1999 (
            .O(N__9252),
            .I(N__9249));
    Odrv4 I__1998 (
            .O(N__9249),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__1997 (
            .O(N__9246),
            .I(N__9243));
    LocalMux I__1996 (
            .O(N__9243),
            .I(N__9240));
    Span4Mux_h I__1995 (
            .O(N__9240),
            .I(N__9237));
    Span4Mux_v I__1994 (
            .O(N__9237),
            .I(N__9234));
    Odrv4 I__1993 (
            .O(N__9234),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__1992 (
            .O(N__9231),
            .I(N__9228));
    LocalMux I__1991 (
            .O(N__9228),
            .I(N__9225));
    Odrv4 I__1990 (
            .O(N__9225),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ));
    IoInMux I__1989 (
            .O(N__9222),
            .I(N__9219));
    LocalMux I__1988 (
            .O(N__9219),
            .I(N__9216));
    Span12Mux_s0_v I__1987 (
            .O(N__9216),
            .I(N__9213));
    Span12Mux_v I__1986 (
            .O(N__9213),
            .I(N__9210));
    Odrv12 I__1985 (
            .O(N__9210),
            .I(CMA_c_0));
    InMux I__1984 (
            .O(N__9207),
            .I(N__9204));
    LocalMux I__1983 (
            .O(N__9204),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5 ));
    InMux I__1982 (
            .O(N__9201),
            .I(N__9198));
    LocalMux I__1981 (
            .O(N__9198),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ));
    CascadeMux I__1980 (
            .O(N__9195),
            .I(\U712_CHIP_RAM.N_147_i_i_a2_0_cascade_ ));
    CEMux I__1979 (
            .O(N__9192),
            .I(N__9189));
    LocalMux I__1978 (
            .O(N__9189),
            .I(N__9185));
    CEMux I__1977 (
            .O(N__9188),
            .I(N__9182));
    Span4Mux_v I__1976 (
            .O(N__9185),
            .I(N__9178));
    LocalMux I__1975 (
            .O(N__9182),
            .I(N__9175));
    CEMux I__1974 (
            .O(N__9181),
            .I(N__9172));
    Span4Mux_h I__1973 (
            .O(N__9178),
            .I(N__9169));
    Span4Mux_h I__1972 (
            .O(N__9175),
            .I(N__9166));
    LocalMux I__1971 (
            .O(N__9172),
            .I(N__9163));
    Odrv4 I__1970 (
            .O(N__9169),
            .I(\U712_CHIP_RAM.N_500_i ));
    Odrv4 I__1969 (
            .O(N__9166),
            .I(\U712_CHIP_RAM.N_500_i ));
    Odrv4 I__1968 (
            .O(N__9163),
            .I(\U712_CHIP_RAM.N_500_i ));
    InMux I__1967 (
            .O(N__9156),
            .I(N__9153));
    LocalMux I__1966 (
            .O(N__9153),
            .I(N__9150));
    Span4Mux_h I__1965 (
            .O(N__9150),
            .I(N__9146));
    InMux I__1964 (
            .O(N__9149),
            .I(N__9143));
    Span4Mux_h I__1963 (
            .O(N__9146),
            .I(N__9140));
    LocalMux I__1962 (
            .O(N__9143),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    Odrv4 I__1961 (
            .O(N__9140),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__1960 (
            .O(N__9135),
            .I(N__9132));
    LocalMux I__1959 (
            .O(N__9132),
            .I(N__9129));
    Span4Mux_h I__1958 (
            .O(N__9129),
            .I(N__9126));
    Odrv4 I__1957 (
            .O(N__9126),
            .I(\U712_CHIP_RAM.REFRESH5lto7_0 ));
    InMux I__1956 (
            .O(N__9123),
            .I(N__9120));
    LocalMux I__1955 (
            .O(N__9120),
            .I(N__9117));
    Span4Mux_h I__1954 (
            .O(N__9117),
            .I(N__9114));
    Span4Mux_h I__1953 (
            .O(N__9114),
            .I(N__9111));
    Odrv4 I__1952 (
            .O(N__9111),
            .I(\U712_CHIP_RAM.REFRESH5lt7 ));
    CascadeMux I__1951 (
            .O(N__9108),
            .I(N__9105));
    InMux I__1950 (
            .O(N__9105),
            .I(N__9102));
    LocalMux I__1949 (
            .O(N__9102),
            .I(N__9097));
    InMux I__1948 (
            .O(N__9101),
            .I(N__9093));
    CascadeMux I__1947 (
            .O(N__9100),
            .I(N__9089));
    Span4Mux_h I__1946 (
            .O(N__9097),
            .I(N__9082));
    InMux I__1945 (
            .O(N__9096),
            .I(N__9079));
    LocalMux I__1944 (
            .O(N__9093),
            .I(N__9076));
    InMux I__1943 (
            .O(N__9092),
            .I(N__9071));
    InMux I__1942 (
            .O(N__9089),
            .I(N__9071));
    InMux I__1941 (
            .O(N__9088),
            .I(N__9068));
    InMux I__1940 (
            .O(N__9087),
            .I(N__9063));
    InMux I__1939 (
            .O(N__9086),
            .I(N__9063));
    InMux I__1938 (
            .O(N__9085),
            .I(N__9060));
    Odrv4 I__1937 (
            .O(N__9082),
            .I(\U712_CHIP_RAM.N_509 ));
    LocalMux I__1936 (
            .O(N__9079),
            .I(\U712_CHIP_RAM.N_509 ));
    Odrv12 I__1935 (
            .O(N__9076),
            .I(\U712_CHIP_RAM.N_509 ));
    LocalMux I__1934 (
            .O(N__9071),
            .I(\U712_CHIP_RAM.N_509 ));
    LocalMux I__1933 (
            .O(N__9068),
            .I(\U712_CHIP_RAM.N_509 ));
    LocalMux I__1932 (
            .O(N__9063),
            .I(\U712_CHIP_RAM.N_509 ));
    LocalMux I__1931 (
            .O(N__9060),
            .I(\U712_CHIP_RAM.N_509 ));
    InMux I__1930 (
            .O(N__9045),
            .I(N__9037));
    InMux I__1929 (
            .O(N__9044),
            .I(N__9037));
    InMux I__1928 (
            .O(N__9043),
            .I(N__9032));
    InMux I__1927 (
            .O(N__9042),
            .I(N__9032));
    LocalMux I__1926 (
            .O(N__9037),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__1925 (
            .O(N__9032),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    InMux I__1924 (
            .O(N__9027),
            .I(N__9022));
    InMux I__1923 (
            .O(N__9026),
            .I(N__9019));
    CascadeMux I__1922 (
            .O(N__9025),
            .I(N__9012));
    LocalMux I__1921 (
            .O(N__9022),
            .I(N__9007));
    LocalMux I__1920 (
            .O(N__9019),
            .I(N__9004));
    InMux I__1919 (
            .O(N__9018),
            .I(N__9001));
    InMux I__1918 (
            .O(N__9017),
            .I(N__8998));
    InMux I__1917 (
            .O(N__9016),
            .I(N__8991));
    InMux I__1916 (
            .O(N__9015),
            .I(N__8991));
    InMux I__1915 (
            .O(N__9012),
            .I(N__8991));
    InMux I__1914 (
            .O(N__9011),
            .I(N__8986));
    InMux I__1913 (
            .O(N__9010),
            .I(N__8986));
    Span4Mux_v I__1912 (
            .O(N__9007),
            .I(N__8979));
    Span4Mux_v I__1911 (
            .O(N__9004),
            .I(N__8979));
    LocalMux I__1910 (
            .O(N__9001),
            .I(N__8979));
    LocalMux I__1909 (
            .O(N__8998),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1908 (
            .O(N__8991),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1907 (
            .O(N__8986),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1906 (
            .O(N__8979),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    InMux I__1905 (
            .O(N__8970),
            .I(N__8966));
    CascadeMux I__1904 (
            .O(N__8969),
            .I(N__8962));
    LocalMux I__1903 (
            .O(N__8966),
            .I(N__8953));
    InMux I__1902 (
            .O(N__8965),
            .I(N__8950));
    InMux I__1901 (
            .O(N__8962),
            .I(N__8947));
    InMux I__1900 (
            .O(N__8961),
            .I(N__8944));
    InMux I__1899 (
            .O(N__8960),
            .I(N__8939));
    InMux I__1898 (
            .O(N__8959),
            .I(N__8939));
    InMux I__1897 (
            .O(N__8958),
            .I(N__8932));
    InMux I__1896 (
            .O(N__8957),
            .I(N__8932));
    InMux I__1895 (
            .O(N__8956),
            .I(N__8932));
    Odrv4 I__1894 (
            .O(N__8953),
            .I(\U712_CHIP_RAM.N_508 ));
    LocalMux I__1893 (
            .O(N__8950),
            .I(\U712_CHIP_RAM.N_508 ));
    LocalMux I__1892 (
            .O(N__8947),
            .I(\U712_CHIP_RAM.N_508 ));
    LocalMux I__1891 (
            .O(N__8944),
            .I(\U712_CHIP_RAM.N_508 ));
    LocalMux I__1890 (
            .O(N__8939),
            .I(\U712_CHIP_RAM.N_508 ));
    LocalMux I__1889 (
            .O(N__8932),
            .I(\U712_CHIP_RAM.N_508 ));
    InMux I__1888 (
            .O(N__8919),
            .I(N__8916));
    LocalMux I__1887 (
            .O(N__8916),
            .I(\U712_CHIP_RAM.N_494 ));
    InMux I__1886 (
            .O(N__8913),
            .I(N__8910));
    LocalMux I__1885 (
            .O(N__8910),
            .I(N__8907));
    Span4Mux_v I__1884 (
            .O(N__8907),
            .I(N__8904));
    Sp12to4 I__1883 (
            .O(N__8904),
            .I(N__8901));
    Span12Mux_h I__1882 (
            .O(N__8901),
            .I(N__8898));
    Span12Mux_h I__1881 (
            .O(N__8898),
            .I(N__8895));
    Odrv12 I__1880 (
            .O(N__8895),
            .I(A_c_12));
    InMux I__1879 (
            .O(N__8892),
            .I(N__8889));
    LocalMux I__1878 (
            .O(N__8889),
            .I(N__8886));
    Span12Mux_v I__1877 (
            .O(N__8886),
            .I(N__8883));
    Span12Mux_h I__1876 (
            .O(N__8883),
            .I(N__8880));
    Odrv12 I__1875 (
            .O(N__8880),
            .I(A_c_13));
    CascadeMux I__1874 (
            .O(N__8877),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ));
    InMux I__1873 (
            .O(N__8874),
            .I(N__8871));
    LocalMux I__1872 (
            .O(N__8871),
            .I(N__8868));
    Span12Mux_v I__1871 (
            .O(N__8868),
            .I(N__8865));
    Span12Mux_h I__1870 (
            .O(N__8865),
            .I(N__8862));
    Odrv12 I__1869 (
            .O(N__8862),
            .I(A_c_5));
    InMux I__1868 (
            .O(N__8859),
            .I(N__8856));
    LocalMux I__1867 (
            .O(N__8856),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ));
    InMux I__1866 (
            .O(N__8853),
            .I(N__8850));
    LocalMux I__1865 (
            .O(N__8850),
            .I(N__8847));
    Span4Mux_h I__1864 (
            .O(N__8847),
            .I(N__8844));
    Span4Mux_v I__1863 (
            .O(N__8844),
            .I(N__8841));
    Sp12to4 I__1862 (
            .O(N__8841),
            .I(N__8838));
    Span12Mux_h I__1861 (
            .O(N__8838),
            .I(N__8835));
    Odrv12 I__1860 (
            .O(N__8835),
            .I(A_c_6));
    InMux I__1859 (
            .O(N__8832),
            .I(N__8829));
    LocalMux I__1858 (
            .O(N__8829),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ));
    CEMux I__1857 (
            .O(N__8826),
            .I(N__8821));
    CEMux I__1856 (
            .O(N__8825),
            .I(N__8818));
    CEMux I__1855 (
            .O(N__8824),
            .I(N__8815));
    LocalMux I__1854 (
            .O(N__8821),
            .I(N__8812));
    LocalMux I__1853 (
            .O(N__8818),
            .I(N__8809));
    LocalMux I__1852 (
            .O(N__8815),
            .I(N__8806));
    Odrv4 I__1851 (
            .O(N__8812),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ));
    Odrv12 I__1850 (
            .O(N__8809),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ));
    Odrv4 I__1849 (
            .O(N__8806),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ));
    InMux I__1848 (
            .O(N__8799),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    CascadeMux I__1847 (
            .O(N__8796),
            .I(N__8793));
    InMux I__1846 (
            .O(N__8793),
            .I(N__8789));
    InMux I__1845 (
            .O(N__8792),
            .I(N__8786));
    LocalMux I__1844 (
            .O(N__8789),
            .I(N__8783));
    LocalMux I__1843 (
            .O(N__8786),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    Odrv4 I__1842 (
            .O(N__8783),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    InMux I__1841 (
            .O(N__8778),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__1840 (
            .O(N__8775),
            .I(N__8771));
    InMux I__1839 (
            .O(N__8774),
            .I(N__8768));
    LocalMux I__1838 (
            .O(N__8771),
            .I(N__8765));
    LocalMux I__1837 (
            .O(N__8768),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    Odrv4 I__1836 (
            .O(N__8765),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__1835 (
            .O(N__8760),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    InMux I__1834 (
            .O(N__8757),
            .I(N__8751));
    InMux I__1833 (
            .O(N__8756),
            .I(N__8746));
    InMux I__1832 (
            .O(N__8755),
            .I(N__8746));
    InMux I__1831 (
            .O(N__8754),
            .I(N__8739));
    LocalMux I__1830 (
            .O(N__8751),
            .I(N__8736));
    LocalMux I__1829 (
            .O(N__8746),
            .I(N__8733));
    InMux I__1828 (
            .O(N__8745),
            .I(N__8724));
    InMux I__1827 (
            .O(N__8744),
            .I(N__8724));
    InMux I__1826 (
            .O(N__8743),
            .I(N__8724));
    InMux I__1825 (
            .O(N__8742),
            .I(N__8724));
    LocalMux I__1824 (
            .O(N__8739),
            .I(N__8721));
    Span4Mux_v I__1823 (
            .O(N__8736),
            .I(N__8718));
    Odrv4 I__1822 (
            .O(N__8733),
            .I(\U712_CHIP_RAM.N_132_i ));
    LocalMux I__1821 (
            .O(N__8724),
            .I(\U712_CHIP_RAM.N_132_i ));
    Odrv4 I__1820 (
            .O(N__8721),
            .I(\U712_CHIP_RAM.N_132_i ));
    Odrv4 I__1819 (
            .O(N__8718),
            .I(\U712_CHIP_RAM.N_132_i ));
    InMux I__1818 (
            .O(N__8709),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    InMux I__1817 (
            .O(N__8706),
            .I(N__8702));
    InMux I__1816 (
            .O(N__8705),
            .I(N__8699));
    LocalMux I__1815 (
            .O(N__8702),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__1814 (
            .O(N__8699),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    InMux I__1813 (
            .O(N__8694),
            .I(N__8685));
    InMux I__1812 (
            .O(N__8693),
            .I(N__8678));
    InMux I__1811 (
            .O(N__8692),
            .I(N__8678));
    InMux I__1810 (
            .O(N__8691),
            .I(N__8678));
    InMux I__1809 (
            .O(N__8690),
            .I(N__8671));
    InMux I__1808 (
            .O(N__8689),
            .I(N__8671));
    InMux I__1807 (
            .O(N__8688),
            .I(N__8671));
    LocalMux I__1806 (
            .O(N__8685),
            .I(N__8668));
    LocalMux I__1805 (
            .O(N__8678),
            .I(N__8663));
    LocalMux I__1804 (
            .O(N__8671),
            .I(N__8663));
    Span4Mux_v I__1803 (
            .O(N__8668),
            .I(N__8660));
    Span4Mux_h I__1802 (
            .O(N__8663),
            .I(N__8657));
    Odrv4 I__1801 (
            .O(N__8660),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    Odrv4 I__1800 (
            .O(N__8657),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    CascadeMux I__1799 (
            .O(N__8652),
            .I(N__8648));
    InMux I__1798 (
            .O(N__8651),
            .I(N__8643));
    InMux I__1797 (
            .O(N__8648),
            .I(N__8640));
    InMux I__1796 (
            .O(N__8647),
            .I(N__8637));
    InMux I__1795 (
            .O(N__8646),
            .I(N__8634));
    LocalMux I__1794 (
            .O(N__8643),
            .I(N__8628));
    LocalMux I__1793 (
            .O(N__8640),
            .I(N__8628));
    LocalMux I__1792 (
            .O(N__8637),
            .I(N__8617));
    LocalMux I__1791 (
            .O(N__8634),
            .I(N__8617));
    InMux I__1790 (
            .O(N__8633),
            .I(N__8612));
    Span4Mux_v I__1789 (
            .O(N__8628),
            .I(N__8609));
    InMux I__1788 (
            .O(N__8627),
            .I(N__8606));
    InMux I__1787 (
            .O(N__8626),
            .I(N__8603));
    InMux I__1786 (
            .O(N__8625),
            .I(N__8596));
    InMux I__1785 (
            .O(N__8624),
            .I(N__8596));
    InMux I__1784 (
            .O(N__8623),
            .I(N__8596));
    InMux I__1783 (
            .O(N__8622),
            .I(N__8593));
    Span4Mux_h I__1782 (
            .O(N__8617),
            .I(N__8590));
    InMux I__1781 (
            .O(N__8616),
            .I(N__8585));
    InMux I__1780 (
            .O(N__8615),
            .I(N__8585));
    LocalMux I__1779 (
            .O(N__8612),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1778 (
            .O(N__8609),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1777 (
            .O(N__8606),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1776 (
            .O(N__8603),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1775 (
            .O(N__8596),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1774 (
            .O(N__8593),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1773 (
            .O(N__8590),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1772 (
            .O(N__8585),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__1771 (
            .O(N__8568),
            .I(N__8565));
    LocalMux I__1770 (
            .O(N__8565),
            .I(\U712_CHIP_RAM.N_436 ));
    InMux I__1769 (
            .O(N__8562),
            .I(N__8559));
    LocalMux I__1768 (
            .O(N__8559),
            .I(N__8556));
    Span4Mux_v I__1767 (
            .O(N__8556),
            .I(N__8553));
    Odrv4 I__1766 (
            .O(N__8553),
            .I(\U712_CHIP_RAM.N_499 ));
    InMux I__1765 (
            .O(N__8550),
            .I(N__8542));
    InMux I__1764 (
            .O(N__8549),
            .I(N__8542));
    InMux I__1763 (
            .O(N__8548),
            .I(N__8538));
    InMux I__1762 (
            .O(N__8547),
            .I(N__8535));
    LocalMux I__1761 (
            .O(N__8542),
            .I(N__8532));
    InMux I__1760 (
            .O(N__8541),
            .I(N__8529));
    LocalMux I__1759 (
            .O(N__8538),
            .I(N__8526));
    LocalMux I__1758 (
            .O(N__8535),
            .I(N__8523));
    Span4Mux_v I__1757 (
            .O(N__8532),
            .I(N__8516));
    LocalMux I__1756 (
            .O(N__8529),
            .I(N__8516));
    Span4Mux_h I__1755 (
            .O(N__8526),
            .I(N__8511));
    Span4Mux_h I__1754 (
            .O(N__8523),
            .I(N__8511));
    InMux I__1753 (
            .O(N__8522),
            .I(N__8508));
    InMux I__1752 (
            .O(N__8521),
            .I(N__8505));
    Span4Mux_h I__1751 (
            .O(N__8516),
            .I(N__8502));
    Span4Mux_v I__1750 (
            .O(N__8511),
            .I(N__8499));
    LocalMux I__1749 (
            .O(N__8508),
            .I(N__8494));
    LocalMux I__1748 (
            .O(N__8505),
            .I(N__8494));
    Odrv4 I__1747 (
            .O(N__8502),
            .I(DMA_CYCLEm));
    Odrv4 I__1746 (
            .O(N__8499),
            .I(DMA_CYCLEm));
    Odrv12 I__1745 (
            .O(N__8494),
            .I(DMA_CYCLEm));
    InMux I__1744 (
            .O(N__8487),
            .I(N__8477));
    InMux I__1743 (
            .O(N__8486),
            .I(N__8477));
    InMux I__1742 (
            .O(N__8485),
            .I(N__8477));
    InMux I__1741 (
            .O(N__8484),
            .I(N__8474));
    LocalMux I__1740 (
            .O(N__8477),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__1739 (
            .O(N__8474),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    CascadeMux I__1738 (
            .O(N__8469),
            .I(N__8464));
    CascadeMux I__1737 (
            .O(N__8468),
            .I(N__8461));
    InMux I__1736 (
            .O(N__8467),
            .I(N__8458));
    InMux I__1735 (
            .O(N__8464),
            .I(N__8453));
    InMux I__1734 (
            .O(N__8461),
            .I(N__8453));
    LocalMux I__1733 (
            .O(N__8458),
            .I(N__8450));
    LocalMux I__1732 (
            .O(N__8453),
            .I(N__8447));
    Odrv4 I__1731 (
            .O(N__8450),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ));
    Odrv12 I__1730 (
            .O(N__8447),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ));
    InMux I__1729 (
            .O(N__8442),
            .I(N__8431));
    InMux I__1728 (
            .O(N__8441),
            .I(N__8427));
    InMux I__1727 (
            .O(N__8440),
            .I(N__8418));
    InMux I__1726 (
            .O(N__8439),
            .I(N__8418));
    InMux I__1725 (
            .O(N__8438),
            .I(N__8410));
    InMux I__1724 (
            .O(N__8437),
            .I(N__8410));
    InMux I__1723 (
            .O(N__8436),
            .I(N__8410));
    CascadeMux I__1722 (
            .O(N__8435),
            .I(N__8406));
    CascadeMux I__1721 (
            .O(N__8434),
            .I(N__8397));
    LocalMux I__1720 (
            .O(N__8431),
            .I(N__8394));
    InMux I__1719 (
            .O(N__8430),
            .I(N__8391));
    LocalMux I__1718 (
            .O(N__8427),
            .I(N__8388));
    CascadeMux I__1717 (
            .O(N__8426),
            .I(N__8385));
    InMux I__1716 (
            .O(N__8425),
            .I(N__8379));
    InMux I__1715 (
            .O(N__8424),
            .I(N__8379));
    InMux I__1714 (
            .O(N__8423),
            .I(N__8376));
    LocalMux I__1713 (
            .O(N__8418),
            .I(N__8373));
    CascadeMux I__1712 (
            .O(N__8417),
            .I(N__8368));
    LocalMux I__1711 (
            .O(N__8410),
            .I(N__8365));
    InMux I__1710 (
            .O(N__8409),
            .I(N__8358));
    InMux I__1709 (
            .O(N__8406),
            .I(N__8358));
    InMux I__1708 (
            .O(N__8405),
            .I(N__8358));
    InMux I__1707 (
            .O(N__8404),
            .I(N__8351));
    InMux I__1706 (
            .O(N__8403),
            .I(N__8351));
    InMux I__1705 (
            .O(N__8402),
            .I(N__8351));
    CascadeMux I__1704 (
            .O(N__8401),
            .I(N__8348));
    InMux I__1703 (
            .O(N__8400),
            .I(N__8343));
    InMux I__1702 (
            .O(N__8397),
            .I(N__8340));
    Span4Mux_v I__1701 (
            .O(N__8394),
            .I(N__8333));
    LocalMux I__1700 (
            .O(N__8391),
            .I(N__8333));
    Span4Mux_v I__1699 (
            .O(N__8388),
            .I(N__8333));
    InMux I__1698 (
            .O(N__8385),
            .I(N__8328));
    InMux I__1697 (
            .O(N__8384),
            .I(N__8328));
    LocalMux I__1696 (
            .O(N__8379),
            .I(N__8321));
    LocalMux I__1695 (
            .O(N__8376),
            .I(N__8321));
    Span4Mux_h I__1694 (
            .O(N__8373),
            .I(N__8321));
    InMux I__1693 (
            .O(N__8372),
            .I(N__8314));
    InMux I__1692 (
            .O(N__8371),
            .I(N__8314));
    InMux I__1691 (
            .O(N__8368),
            .I(N__8314));
    Span4Mux_h I__1690 (
            .O(N__8365),
            .I(N__8307));
    LocalMux I__1689 (
            .O(N__8358),
            .I(N__8307));
    LocalMux I__1688 (
            .O(N__8351),
            .I(N__8307));
    InMux I__1687 (
            .O(N__8348),
            .I(N__8300));
    InMux I__1686 (
            .O(N__8347),
            .I(N__8300));
    InMux I__1685 (
            .O(N__8346),
            .I(N__8300));
    LocalMux I__1684 (
            .O(N__8343),
            .I(N__8297));
    LocalMux I__1683 (
            .O(N__8340),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1682 (
            .O(N__8333),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1681 (
            .O(N__8328),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1680 (
            .O(N__8321),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1679 (
            .O(N__8314),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1678 (
            .O(N__8307),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1677 (
            .O(N__8300),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1676 (
            .O(N__8297),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    CascadeMux I__1675 (
            .O(N__8280),
            .I(\U712_CHIP_RAM.N_506_cascade_ ));
    InMux I__1674 (
            .O(N__8277),
            .I(N__8274));
    LocalMux I__1673 (
            .O(N__8274),
            .I(\U712_CHIP_RAM.N_147_i_i_a2_0 ));
    InMux I__1672 (
            .O(N__8271),
            .I(N__8268));
    LocalMux I__1671 (
            .O(N__8268),
            .I(N__8265));
    Span4Mux_h I__1670 (
            .O(N__8265),
            .I(N__8261));
    InMux I__1669 (
            .O(N__8264),
            .I(N__8258));
    Odrv4 I__1668 (
            .O(N__8261),
            .I(\U712_CHIP_RAM.N_359 ));
    LocalMux I__1667 (
            .O(N__8258),
            .I(\U712_CHIP_RAM.N_359 ));
    InMux I__1666 (
            .O(N__8253),
            .I(N__8250));
    LocalMux I__1665 (
            .O(N__8250),
            .I(\U712_CHIP_RAM.N_595 ));
    CascadeMux I__1664 (
            .O(N__8247),
            .I(N__8244));
    InMux I__1663 (
            .O(N__8244),
            .I(N__8240));
    InMux I__1662 (
            .O(N__8243),
            .I(N__8236));
    LocalMux I__1661 (
            .O(N__8240),
            .I(N__8232));
    InMux I__1660 (
            .O(N__8239),
            .I(N__8229));
    LocalMux I__1659 (
            .O(N__8236),
            .I(N__8226));
    CascadeMux I__1658 (
            .O(N__8235),
            .I(N__8223));
    Span4Mux_h I__1657 (
            .O(N__8232),
            .I(N__8218));
    LocalMux I__1656 (
            .O(N__8229),
            .I(N__8218));
    Span4Mux_h I__1655 (
            .O(N__8226),
            .I(N__8215));
    InMux I__1654 (
            .O(N__8223),
            .I(N__8212));
    Odrv4 I__1653 (
            .O(N__8218),
            .I(\U712_CHIP_RAM.N_348 ));
    Odrv4 I__1652 (
            .O(N__8215),
            .I(\U712_CHIP_RAM.N_348 ));
    LocalMux I__1651 (
            .O(N__8212),
            .I(\U712_CHIP_RAM.N_348 ));
    CascadeMux I__1650 (
            .O(N__8205),
            .I(\U712_CHIP_RAM.N_595_cascade_ ));
    InMux I__1649 (
            .O(N__8202),
            .I(N__8196));
    InMux I__1648 (
            .O(N__8201),
            .I(N__8191));
    InMux I__1647 (
            .O(N__8200),
            .I(N__8191));
    InMux I__1646 (
            .O(N__8199),
            .I(N__8188));
    LocalMux I__1645 (
            .O(N__8196),
            .I(\U712_CHIP_RAM.N_577 ));
    LocalMux I__1644 (
            .O(N__8191),
            .I(\U712_CHIP_RAM.N_577 ));
    LocalMux I__1643 (
            .O(N__8188),
            .I(\U712_CHIP_RAM.N_577 ));
    InMux I__1642 (
            .O(N__8181),
            .I(N__8178));
    LocalMux I__1641 (
            .O(N__8178),
            .I(N__8175));
    Odrv4 I__1640 (
            .O(N__8175),
            .I(\U712_CHIP_RAM.N_279 ));
    CascadeMux I__1639 (
            .O(N__8172),
            .I(N__8168));
    InMux I__1638 (
            .O(N__8171),
            .I(N__8158));
    InMux I__1637 (
            .O(N__8168),
            .I(N__8153));
    InMux I__1636 (
            .O(N__8167),
            .I(N__8153));
    InMux I__1635 (
            .O(N__8166),
            .I(N__8150));
    InMux I__1634 (
            .O(N__8165),
            .I(N__8147));
    InMux I__1633 (
            .O(N__8164),
            .I(N__8142));
    InMux I__1632 (
            .O(N__8163),
            .I(N__8142));
    InMux I__1631 (
            .O(N__8162),
            .I(N__8137));
    InMux I__1630 (
            .O(N__8161),
            .I(N__8137));
    LocalMux I__1629 (
            .O(N__8158),
            .I(N__8130));
    LocalMux I__1628 (
            .O(N__8153),
            .I(N__8130));
    LocalMux I__1627 (
            .O(N__8150),
            .I(N__8130));
    LocalMux I__1626 (
            .O(N__8147),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1625 (
            .O(N__8142),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1624 (
            .O(N__8137),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1623 (
            .O(N__8130),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    InMux I__1622 (
            .O(N__8121),
            .I(N__8118));
    LocalMux I__1621 (
            .O(N__8118),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_i_a2_0_1 ));
    CascadeMux I__1620 (
            .O(N__8115),
            .I(N__8107));
    InMux I__1619 (
            .O(N__8114),
            .I(N__8100));
    InMux I__1618 (
            .O(N__8113),
            .I(N__8100));
    CascadeMux I__1617 (
            .O(N__8112),
            .I(N__8095));
    InMux I__1616 (
            .O(N__8111),
            .I(N__8085));
    InMux I__1615 (
            .O(N__8110),
            .I(N__8085));
    InMux I__1614 (
            .O(N__8107),
            .I(N__8085));
    InMux I__1613 (
            .O(N__8106),
            .I(N__8085));
    InMux I__1612 (
            .O(N__8105),
            .I(N__8076));
    LocalMux I__1611 (
            .O(N__8100),
            .I(N__8073));
    InMux I__1610 (
            .O(N__8099),
            .I(N__8064));
    InMux I__1609 (
            .O(N__8098),
            .I(N__8064));
    InMux I__1608 (
            .O(N__8095),
            .I(N__8064));
    InMux I__1607 (
            .O(N__8094),
            .I(N__8064));
    LocalMux I__1606 (
            .O(N__8085),
            .I(N__8061));
    InMux I__1605 (
            .O(N__8084),
            .I(N__8056));
    InMux I__1604 (
            .O(N__8083),
            .I(N__8056));
    InMux I__1603 (
            .O(N__8082),
            .I(N__8051));
    InMux I__1602 (
            .O(N__8081),
            .I(N__8051));
    InMux I__1601 (
            .O(N__8080),
            .I(N__8048));
    InMux I__1600 (
            .O(N__8079),
            .I(N__8045));
    LocalMux I__1599 (
            .O(N__8076),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1598 (
            .O(N__8073),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1597 (
            .O(N__8064),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1596 (
            .O(N__8061),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1595 (
            .O(N__8056),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1594 (
            .O(N__8051),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1593 (
            .O(N__8048),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1592 (
            .O(N__8045),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    InMux I__1591 (
            .O(N__8028),
            .I(N__8024));
    InMux I__1590 (
            .O(N__8027),
            .I(N__8021));
    LocalMux I__1589 (
            .O(N__8024),
            .I(N__8018));
    LocalMux I__1588 (
            .O(N__8021),
            .I(N__8015));
    Span4Mux_v I__1587 (
            .O(N__8018),
            .I(N__8010));
    Span4Mux_h I__1586 (
            .O(N__8015),
            .I(N__8010));
    Odrv4 I__1585 (
            .O(N__8010),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_a2_0 ));
    InMux I__1584 (
            .O(N__8007),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__1583 (
            .O(N__8004),
            .I(N__8001));
    LocalMux I__1582 (
            .O(N__8001),
            .I(N__7998));
    Span12Mux_h I__1581 (
            .O(N__7998),
            .I(N__7995));
    Odrv12 I__1580 (
            .O(N__7995),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    InMux I__1579 (
            .O(N__7992),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    CascadeMux I__1578 (
            .O(N__7989),
            .I(N__7985));
    CascadeMux I__1577 (
            .O(N__7988),
            .I(N__7981));
    InMux I__1576 (
            .O(N__7985),
            .I(N__7978));
    InMux I__1575 (
            .O(N__7984),
            .I(N__7975));
    InMux I__1574 (
            .O(N__7981),
            .I(N__7971));
    LocalMux I__1573 (
            .O(N__7978),
            .I(N__7966));
    LocalMux I__1572 (
            .O(N__7975),
            .I(N__7963));
    CascadeMux I__1571 (
            .O(N__7974),
            .I(N__7958));
    LocalMux I__1570 (
            .O(N__7971),
            .I(N__7954));
    InMux I__1569 (
            .O(N__7970),
            .I(N__7951));
    InMux I__1568 (
            .O(N__7969),
            .I(N__7947));
    Span4Mux_h I__1567 (
            .O(N__7966),
            .I(N__7942));
    Span4Mux_v I__1566 (
            .O(N__7963),
            .I(N__7942));
    InMux I__1565 (
            .O(N__7962),
            .I(N__7937));
    InMux I__1564 (
            .O(N__7961),
            .I(N__7937));
    InMux I__1563 (
            .O(N__7958),
            .I(N__7932));
    InMux I__1562 (
            .O(N__7957),
            .I(N__7932));
    Span4Mux_v I__1561 (
            .O(N__7954),
            .I(N__7927));
    LocalMux I__1560 (
            .O(N__7951),
            .I(N__7927));
    InMux I__1559 (
            .O(N__7950),
            .I(N__7924));
    LocalMux I__1558 (
            .O(N__7947),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1557 (
            .O(N__7942),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1556 (
            .O(N__7937),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1555 (
            .O(N__7932),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1554 (
            .O(N__7927),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1553 (
            .O(N__7924),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    InMux I__1552 (
            .O(N__7911),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    InMux I__1551 (
            .O(N__7908),
            .I(N__7904));
    InMux I__1550 (
            .O(N__7907),
            .I(N__7901));
    LocalMux I__1549 (
            .O(N__7904),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1548 (
            .O(N__7901),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    CascadeMux I__1547 (
            .O(N__7896),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0_cascade_ ));
    IoInMux I__1546 (
            .O(N__7893),
            .I(N__7890));
    LocalMux I__1545 (
            .O(N__7890),
            .I(N__7887));
    Span12Mux_s9_v I__1544 (
            .O(N__7887),
            .I(N__7884));
    Span12Mux_h I__1543 (
            .O(N__7884),
            .I(N__7880));
    InMux I__1542 (
            .O(N__7883),
            .I(N__7877));
    Odrv12 I__1541 (
            .O(N__7880),
            .I(LATCH_CLK_c));
    LocalMux I__1540 (
            .O(N__7877),
            .I(LATCH_CLK_c));
    InMux I__1539 (
            .O(N__7872),
            .I(N__7869));
    LocalMux I__1538 (
            .O(N__7869),
            .I(N__7866));
    Span12Mux_h I__1537 (
            .O(N__7866),
            .I(N__7863));
    Odrv12 I__1536 (
            .O(N__7863),
            .I(DBRn_c_i));
    InMux I__1535 (
            .O(N__7860),
            .I(N__7857));
    LocalMux I__1534 (
            .O(N__7857),
            .I(N__7854));
    Span4Mux_h I__1533 (
            .O(N__7854),
            .I(N__7850));
    InMux I__1532 (
            .O(N__7853),
            .I(N__7847));
    Span4Mux_v I__1531 (
            .O(N__7850),
            .I(N__7844));
    LocalMux I__1530 (
            .O(N__7847),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    Odrv4 I__1529 (
            .O(N__7844),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    IoInMux I__1528 (
            .O(N__7839),
            .I(N__7836));
    LocalMux I__1527 (
            .O(N__7836),
            .I(N__7833));
    Span12Mux_s6_v I__1526 (
            .O(N__7833),
            .I(N__7830));
    Odrv12 I__1525 (
            .O(N__7830),
            .I(N_119_i));
    InMux I__1524 (
            .O(N__7827),
            .I(N__7821));
    InMux I__1523 (
            .O(N__7826),
            .I(N__7818));
    InMux I__1522 (
            .O(N__7825),
            .I(N__7813));
    InMux I__1521 (
            .O(N__7824),
            .I(N__7813));
    LocalMux I__1520 (
            .O(N__7821),
            .I(N__7810));
    LocalMux I__1519 (
            .O(N__7818),
            .I(N__7807));
    LocalMux I__1518 (
            .O(N__7813),
            .I(N__7804));
    Span4Mux_v I__1517 (
            .O(N__7810),
            .I(N__7797));
    Span4Mux_h I__1516 (
            .O(N__7807),
            .I(N__7792));
    Span4Mux_v I__1515 (
            .O(N__7804),
            .I(N__7792));
    InMux I__1514 (
            .O(N__7803),
            .I(N__7787));
    InMux I__1513 (
            .O(N__7802),
            .I(N__7787));
    InMux I__1512 (
            .O(N__7801),
            .I(N__7782));
    InMux I__1511 (
            .O(N__7800),
            .I(N__7782));
    Span4Mux_v I__1510 (
            .O(N__7797),
            .I(N__7779));
    Span4Mux_v I__1509 (
            .O(N__7792),
            .I(N__7776));
    LocalMux I__1508 (
            .O(N__7787),
            .I(N__7771));
    LocalMux I__1507 (
            .O(N__7782),
            .I(N__7771));
    Span4Mux_v I__1506 (
            .O(N__7779),
            .I(N__7768));
    Span4Mux_v I__1505 (
            .O(N__7776),
            .I(N__7763));
    Span4Mux_v I__1504 (
            .O(N__7771),
            .I(N__7763));
    Sp12to4 I__1503 (
            .O(N__7768),
            .I(N__7758));
    Sp12to4 I__1502 (
            .O(N__7763),
            .I(N__7758));
    Span12Mux_h I__1501 (
            .O(N__7758),
            .I(N__7755));
    Odrv12 I__1500 (
            .O(N__7755),
            .I(A_c_1));
    CascadeMux I__1499 (
            .O(N__7752),
            .I(N__7745));
    InMux I__1498 (
            .O(N__7751),
            .I(N__7740));
    InMux I__1497 (
            .O(N__7750),
            .I(N__7740));
    CascadeMux I__1496 (
            .O(N__7749),
            .I(N__7737));
    InMux I__1495 (
            .O(N__7748),
            .I(N__7733));
    InMux I__1494 (
            .O(N__7745),
            .I(N__7727));
    LocalMux I__1493 (
            .O(N__7740),
            .I(N__7724));
    InMux I__1492 (
            .O(N__7737),
            .I(N__7719));
    InMux I__1491 (
            .O(N__7736),
            .I(N__7719));
    LocalMux I__1490 (
            .O(N__7733),
            .I(N__7716));
    InMux I__1489 (
            .O(N__7732),
            .I(N__7713));
    InMux I__1488 (
            .O(N__7731),
            .I(N__7710));
    InMux I__1487 (
            .O(N__7730),
            .I(N__7707));
    LocalMux I__1486 (
            .O(N__7727),
            .I(N__7704));
    Span4Mux_v I__1485 (
            .O(N__7724),
            .I(N__7699));
    LocalMux I__1484 (
            .O(N__7719),
            .I(N__7699));
    Span4Mux_v I__1483 (
            .O(N__7716),
            .I(N__7692));
    LocalMux I__1482 (
            .O(N__7713),
            .I(N__7692));
    LocalMux I__1481 (
            .O(N__7710),
            .I(N__7692));
    LocalMux I__1480 (
            .O(N__7707),
            .I(N__7689));
    Span4Mux_v I__1479 (
            .O(N__7704),
            .I(N__7686));
    Span4Mux_h I__1478 (
            .O(N__7699),
            .I(N__7683));
    Span4Mux_h I__1477 (
            .O(N__7692),
            .I(N__7678));
    Span4Mux_v I__1476 (
            .O(N__7689),
            .I(N__7678));
    Span4Mux_v I__1475 (
            .O(N__7686),
            .I(N__7675));
    Span4Mux_v I__1474 (
            .O(N__7683),
            .I(N__7670));
    Span4Mux_v I__1473 (
            .O(N__7678),
            .I(N__7670));
    Sp12to4 I__1472 (
            .O(N__7675),
            .I(N__7665));
    Sp12to4 I__1471 (
            .O(N__7670),
            .I(N__7665));
    Span12Mux_h I__1470 (
            .O(N__7665),
            .I(N__7662));
    Odrv12 I__1469 (
            .O(N__7662),
            .I(A_c_0));
    CascadeMux I__1468 (
            .O(N__7659),
            .I(N__7655));
    CascadeMux I__1467 (
            .O(N__7658),
            .I(N__7652));
    InMux I__1466 (
            .O(N__7655),
            .I(N__7647));
    InMux I__1465 (
            .O(N__7652),
            .I(N__7642));
    InMux I__1464 (
            .O(N__7651),
            .I(N__7642));
    CascadeMux I__1463 (
            .O(N__7650),
            .I(N__7638));
    LocalMux I__1462 (
            .O(N__7647),
            .I(N__7635));
    LocalMux I__1461 (
            .O(N__7642),
            .I(N__7630));
    InMux I__1460 (
            .O(N__7641),
            .I(N__7625));
    InMux I__1459 (
            .O(N__7638),
            .I(N__7625));
    Span4Mux_v I__1458 (
            .O(N__7635),
            .I(N__7622));
    InMux I__1457 (
            .O(N__7634),
            .I(N__7619));
    InMux I__1456 (
            .O(N__7633),
            .I(N__7616));
    Span4Mux_h I__1455 (
            .O(N__7630),
            .I(N__7610));
    LocalMux I__1454 (
            .O(N__7625),
            .I(N__7610));
    Span4Mux_h I__1453 (
            .O(N__7622),
            .I(N__7607));
    LocalMux I__1452 (
            .O(N__7619),
            .I(N__7604));
    LocalMux I__1451 (
            .O(N__7616),
            .I(N__7601));
    InMux I__1450 (
            .O(N__7615),
            .I(N__7598));
    Span4Mux_h I__1449 (
            .O(N__7610),
            .I(N__7595));
    Sp12to4 I__1448 (
            .O(N__7607),
            .I(N__7586));
    Span12Mux_h I__1447 (
            .O(N__7604),
            .I(N__7586));
    Sp12to4 I__1446 (
            .O(N__7601),
            .I(N__7586));
    LocalMux I__1445 (
            .O(N__7598),
            .I(N__7586));
    Span4Mux_v I__1444 (
            .O(N__7595),
            .I(N__7583));
    Span12Mux_h I__1443 (
            .O(N__7586),
            .I(N__7580));
    Span4Mux_h I__1442 (
            .O(N__7583),
            .I(N__7577));
    Span12Mux_v I__1441 (
            .O(N__7580),
            .I(N__7574));
    Sp12to4 I__1440 (
            .O(N__7577),
            .I(N__7571));
    Odrv12 I__1439 (
            .O(N__7574),
            .I(SIZ_c_0));
    Odrv12 I__1438 (
            .O(N__7571),
            .I(SIZ_c_0));
    CascadeMux I__1437 (
            .O(N__7566),
            .I(N__7562));
    InMux I__1436 (
            .O(N__7565),
            .I(N__7554));
    InMux I__1435 (
            .O(N__7562),
            .I(N__7554));
    InMux I__1434 (
            .O(N__7561),
            .I(N__7550));
    CascadeMux I__1433 (
            .O(N__7560),
            .I(N__7547));
    CascadeMux I__1432 (
            .O(N__7559),
            .I(N__7544));
    LocalMux I__1431 (
            .O(N__7554),
            .I(N__7540));
    InMux I__1430 (
            .O(N__7553),
            .I(N__7537));
    LocalMux I__1429 (
            .O(N__7550),
            .I(N__7532));
    InMux I__1428 (
            .O(N__7547),
            .I(N__7529));
    InMux I__1427 (
            .O(N__7544),
            .I(N__7526));
    InMux I__1426 (
            .O(N__7543),
            .I(N__7523));
    Span4Mux_h I__1425 (
            .O(N__7540),
            .I(N__7520));
    LocalMux I__1424 (
            .O(N__7537),
            .I(N__7517));
    InMux I__1423 (
            .O(N__7536),
            .I(N__7512));
    InMux I__1422 (
            .O(N__7535),
            .I(N__7512));
    Sp12to4 I__1421 (
            .O(N__7532),
            .I(N__7509));
    LocalMux I__1420 (
            .O(N__7529),
            .I(N__7502));
    LocalMux I__1419 (
            .O(N__7526),
            .I(N__7502));
    LocalMux I__1418 (
            .O(N__7523),
            .I(N__7502));
    Span4Mux_v I__1417 (
            .O(N__7520),
            .I(N__7499));
    Span12Mux_v I__1416 (
            .O(N__7517),
            .I(N__7494));
    LocalMux I__1415 (
            .O(N__7512),
            .I(N__7494));
    Span12Mux_v I__1414 (
            .O(N__7509),
            .I(N__7491));
    Span12Mux_h I__1413 (
            .O(N__7502),
            .I(N__7488));
    Sp12to4 I__1412 (
            .O(N__7499),
            .I(N__7483));
    Span12Mux_v I__1411 (
            .O(N__7494),
            .I(N__7483));
    Span12Mux_h I__1410 (
            .O(N__7491),
            .I(N__7480));
    Span12Mux_v I__1409 (
            .O(N__7488),
            .I(N__7477));
    Span12Mux_h I__1408 (
            .O(N__7483),
            .I(N__7474));
    Odrv12 I__1407 (
            .O(N__7480),
            .I(SIZ_c_1));
    Odrv12 I__1406 (
            .O(N__7477),
            .I(SIZ_c_1));
    Odrv12 I__1405 (
            .O(N__7474),
            .I(SIZ_c_1));
    IoInMux I__1404 (
            .O(N__7467),
            .I(N__7464));
    LocalMux I__1403 (
            .O(N__7464),
            .I(N__7461));
    Span4Mux_s3_v I__1402 (
            .O(N__7461),
            .I(N__7458));
    Odrv4 I__1401 (
            .O(N__7458),
            .I(N_61_i));
    IoInMux I__1400 (
            .O(N__7455),
            .I(N__7452));
    LocalMux I__1399 (
            .O(N__7452),
            .I(N__7449));
    Span4Mux_s0_v I__1398 (
            .O(N__7449),
            .I(N__7446));
    Span4Mux_v I__1397 (
            .O(N__7446),
            .I(N__7443));
    Span4Mux_v I__1396 (
            .O(N__7443),
            .I(N__7440));
    Span4Mux_h I__1395 (
            .O(N__7440),
            .I(N__7437));
    Odrv4 I__1394 (
            .O(N__7437),
            .I(CMA_c_2));
    InMux I__1393 (
            .O(N__7434),
            .I(N__7431));
    LocalMux I__1392 (
            .O(N__7431),
            .I(N__7428));
    Span4Mux_v I__1391 (
            .O(N__7428),
            .I(N__7425));
    Odrv4 I__1390 (
            .O(N__7425),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ));
    InMux I__1389 (
            .O(N__7422),
            .I(N__7419));
    LocalMux I__1388 (
            .O(N__7419),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ));
    IoInMux I__1387 (
            .O(N__7416),
            .I(N__7412));
    InMux I__1386 (
            .O(N__7415),
            .I(N__7409));
    LocalMux I__1385 (
            .O(N__7412),
            .I(N__7406));
    LocalMux I__1384 (
            .O(N__7409),
            .I(N__7403));
    Span4Mux_s3_v I__1383 (
            .O(N__7406),
            .I(N__7400));
    Span4Mux_v I__1382 (
            .O(N__7403),
            .I(N__7397));
    Odrv4 I__1381 (
            .O(N__7400),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1380 (
            .O(N__7397),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__1379 (
            .O(N__7392),
            .I(N__7389));
    InMux I__1378 (
            .O(N__7389),
            .I(N__7386));
    LocalMux I__1377 (
            .O(N__7386),
            .I(N__7383));
    Span4Mux_h I__1376 (
            .O(N__7383),
            .I(N__7380));
    Odrv4 I__1375 (
            .O(N__7380),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ));
    InMux I__1374 (
            .O(N__7377),
            .I(N__7374));
    LocalMux I__1373 (
            .O(N__7374),
            .I(\U712_CHIP_RAM.N_431 ));
    InMux I__1372 (
            .O(N__7371),
            .I(N__7368));
    LocalMux I__1371 (
            .O(N__7368),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3 ));
    InMux I__1370 (
            .O(N__7365),
            .I(N__7362));
    LocalMux I__1369 (
            .O(N__7362),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ));
    IoInMux I__1368 (
            .O(N__7359),
            .I(N__7356));
    LocalMux I__1367 (
            .O(N__7356),
            .I(N__7353));
    IoSpan4Mux I__1366 (
            .O(N__7353),
            .I(N__7350));
    Span4Mux_s2_v I__1365 (
            .O(N__7350),
            .I(N__7346));
    InMux I__1364 (
            .O(N__7349),
            .I(N__7343));
    Sp12to4 I__1363 (
            .O(N__7346),
            .I(N__7340));
    LocalMux I__1362 (
            .O(N__7343),
            .I(N__7337));
    Span12Mux_s8_v I__1361 (
            .O(N__7340),
            .I(N__7334));
    Sp12to4 I__1360 (
            .O(N__7337),
            .I(N__7331));
    Span12Mux_h I__1359 (
            .O(N__7334),
            .I(N__7328));
    Span12Mux_v I__1358 (
            .O(N__7331),
            .I(N__7325));
    Span12Mux_v I__1357 (
            .O(N__7328),
            .I(N__7322));
    Span12Mux_h I__1356 (
            .O(N__7325),
            .I(N__7319));
    Odrv12 I__1355 (
            .O(N__7322),
            .I(A_c_11));
    Odrv12 I__1354 (
            .O(N__7319),
            .I(A_c_11));
    InMux I__1353 (
            .O(N__7314),
            .I(N__7310));
    InMux I__1352 (
            .O(N__7313),
            .I(N__7307));
    LocalMux I__1351 (
            .O(N__7310),
            .I(\U712_CHIP_RAM.N_350 ));
    LocalMux I__1350 (
            .O(N__7307),
            .I(\U712_CHIP_RAM.N_350 ));
    InMux I__1349 (
            .O(N__7302),
            .I(N__7299));
    LocalMux I__1348 (
            .O(N__7299),
            .I(\U712_CHIP_RAM.N_452 ));
    IoInMux I__1347 (
            .O(N__7296),
            .I(N__7292));
    InMux I__1346 (
            .O(N__7295),
            .I(N__7289));
    LocalMux I__1345 (
            .O(N__7292),
            .I(N__7286));
    LocalMux I__1344 (
            .O(N__7289),
            .I(N__7283));
    Span12Mux_s4_v I__1343 (
            .O(N__7286),
            .I(N__7280));
    Span4Mux_v I__1342 (
            .O(N__7283),
            .I(N__7277));
    Span12Mux_v I__1341 (
            .O(N__7280),
            .I(N__7274));
    Sp12to4 I__1340 (
            .O(N__7277),
            .I(N__7271));
    Span12Mux_h I__1339 (
            .O(N__7274),
            .I(N__7268));
    Span12Mux_h I__1338 (
            .O(N__7271),
            .I(N__7265));
    Odrv12 I__1337 (
            .O(N__7268),
            .I(A_c_9));
    Odrv12 I__1336 (
            .O(N__7265),
            .I(A_c_9));
    InMux I__1335 (
            .O(N__7260),
            .I(N__7257));
    LocalMux I__1334 (
            .O(N__7257),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ));
    CascadeMux I__1333 (
            .O(N__7254),
            .I(\U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a2_1_cascade_ ));
    InMux I__1332 (
            .O(N__7251),
            .I(N__7245));
    InMux I__1331 (
            .O(N__7250),
            .I(N__7242));
    CascadeMux I__1330 (
            .O(N__7249),
            .I(N__7239));
    CascadeMux I__1329 (
            .O(N__7248),
            .I(N__7235));
    LocalMux I__1328 (
            .O(N__7245),
            .I(N__7230));
    LocalMux I__1327 (
            .O(N__7242),
            .I(N__7227));
    InMux I__1326 (
            .O(N__7239),
            .I(N__7222));
    InMux I__1325 (
            .O(N__7238),
            .I(N__7222));
    InMux I__1324 (
            .O(N__7235),
            .I(N__7217));
    InMux I__1323 (
            .O(N__7234),
            .I(N__7217));
    InMux I__1322 (
            .O(N__7233),
            .I(N__7214));
    Odrv12 I__1321 (
            .O(N__7230),
            .I(\U712_CHIP_RAM.N_344 ));
    Odrv4 I__1320 (
            .O(N__7227),
            .I(\U712_CHIP_RAM.N_344 ));
    LocalMux I__1319 (
            .O(N__7222),
            .I(\U712_CHIP_RAM.N_344 ));
    LocalMux I__1318 (
            .O(N__7217),
            .I(\U712_CHIP_RAM.N_344 ));
    LocalMux I__1317 (
            .O(N__7214),
            .I(\U712_CHIP_RAM.N_344 ));
    InMux I__1316 (
            .O(N__7203),
            .I(N__7200));
    LocalMux I__1315 (
            .O(N__7200),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_0 ));
    CascadeMux I__1314 (
            .O(N__7197),
            .I(\U712_CHIP_RAM.N_72_cascade_ ));
    InMux I__1313 (
            .O(N__7194),
            .I(N__7191));
    LocalMux I__1312 (
            .O(N__7191),
            .I(N__7188));
    Span4Mux_h I__1311 (
            .O(N__7188),
            .I(N__7184));
    InMux I__1310 (
            .O(N__7187),
            .I(N__7181));
    Odrv4 I__1309 (
            .O(N__7184),
            .I(CPU_TACKm));
    LocalMux I__1308 (
            .O(N__7181),
            .I(CPU_TACKm));
    InMux I__1307 (
            .O(N__7176),
            .I(N__7173));
    LocalMux I__1306 (
            .O(N__7173),
            .I(\U712_CHIP_RAM.N_462 ));
    InMux I__1305 (
            .O(N__7170),
            .I(N__7164));
    InMux I__1304 (
            .O(N__7169),
            .I(N__7159));
    InMux I__1303 (
            .O(N__7168),
            .I(N__7159));
    InMux I__1302 (
            .O(N__7167),
            .I(N__7155));
    LocalMux I__1301 (
            .O(N__7164),
            .I(N__7152));
    LocalMux I__1300 (
            .O(N__7159),
            .I(N__7149));
    InMux I__1299 (
            .O(N__7158),
            .I(N__7146));
    LocalMux I__1298 (
            .O(N__7155),
            .I(N__7142));
    Span4Mux_v I__1297 (
            .O(N__7152),
            .I(N__7134));
    Span4Mux_v I__1296 (
            .O(N__7149),
            .I(N__7134));
    LocalMux I__1295 (
            .O(N__7146),
            .I(N__7131));
    InMux I__1294 (
            .O(N__7145),
            .I(N__7128));
    Span4Mux_h I__1293 (
            .O(N__7142),
            .I(N__7125));
    InMux I__1292 (
            .O(N__7141),
            .I(N__7118));
    InMux I__1291 (
            .O(N__7140),
            .I(N__7118));
    InMux I__1290 (
            .O(N__7139),
            .I(N__7118));
    Odrv4 I__1289 (
            .O(N__7134),
            .I(\U712_CHIP_RAM.N_503 ));
    Odrv12 I__1288 (
            .O(N__7131),
            .I(\U712_CHIP_RAM.N_503 ));
    LocalMux I__1287 (
            .O(N__7128),
            .I(\U712_CHIP_RAM.N_503 ));
    Odrv4 I__1286 (
            .O(N__7125),
            .I(\U712_CHIP_RAM.N_503 ));
    LocalMux I__1285 (
            .O(N__7118),
            .I(\U712_CHIP_RAM.N_503 ));
    CascadeMux I__1284 (
            .O(N__7107),
            .I(\U712_CHIP_RAM.N_462_cascade_ ));
    InMux I__1283 (
            .O(N__7104),
            .I(N__7095));
    InMux I__1282 (
            .O(N__7103),
            .I(N__7095));
    InMux I__1281 (
            .O(N__7102),
            .I(N__7090));
    InMux I__1280 (
            .O(N__7101),
            .I(N__7090));
    InMux I__1279 (
            .O(N__7100),
            .I(N__7085));
    LocalMux I__1278 (
            .O(N__7095),
            .I(N__7082));
    LocalMux I__1277 (
            .O(N__7090),
            .I(N__7079));
    InMux I__1276 (
            .O(N__7089),
            .I(N__7074));
    InMux I__1275 (
            .O(N__7088),
            .I(N__7074));
    LocalMux I__1274 (
            .O(N__7085),
            .I(\U712_CHIP_RAM.N_510 ));
    Odrv12 I__1273 (
            .O(N__7082),
            .I(\U712_CHIP_RAM.N_510 ));
    Odrv4 I__1272 (
            .O(N__7079),
            .I(\U712_CHIP_RAM.N_510 ));
    LocalMux I__1271 (
            .O(N__7074),
            .I(\U712_CHIP_RAM.N_510 ));
    CascadeMux I__1270 (
            .O(N__7065),
            .I(\U712_CHIP_RAM.N_347_cascade_ ));
    InMux I__1269 (
            .O(N__7062),
            .I(N__7059));
    LocalMux I__1268 (
            .O(N__7059),
            .I(\U712_CHIP_RAM.N_590 ));
    CascadeMux I__1267 (
            .O(N__7056),
            .I(\U712_CHIP_RAM.N_590_cascade_ ));
    InMux I__1266 (
            .O(N__7053),
            .I(N__7050));
    LocalMux I__1265 (
            .O(N__7050),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0 ));
    InMux I__1264 (
            .O(N__7047),
            .I(N__7043));
    InMux I__1263 (
            .O(N__7046),
            .I(N__7040));
    LocalMux I__1262 (
            .O(N__7043),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0 ));
    LocalMux I__1261 (
            .O(N__7040),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0 ));
    CascadeMux I__1260 (
            .O(N__7035),
            .I(\U712_CHIP_RAM.N_509_cascade_ ));
    CascadeMux I__1259 (
            .O(N__7032),
            .I(N__7029));
    InMux I__1258 (
            .O(N__7029),
            .I(N__7026));
    LocalMux I__1257 (
            .O(N__7026),
            .I(N__7023));
    Span4Mux_h I__1256 (
            .O(N__7023),
            .I(N__7020));
    Odrv4 I__1255 (
            .O(N__7020),
            .I(\U712_CHIP_RAM.DBENn_8_0_0 ));
    InMux I__1254 (
            .O(N__7017),
            .I(N__7014));
    LocalMux I__1253 (
            .O(N__7014),
            .I(N__7010));
    InMux I__1252 (
            .O(N__7013),
            .I(N__7007));
    Span4Mux_v I__1251 (
            .O(N__7010),
            .I(N__7004));
    LocalMux I__1250 (
            .O(N__7007),
            .I(N__7001));
    Sp12to4 I__1249 (
            .O(N__7004),
            .I(N__6998));
    Span12Mux_v I__1248 (
            .O(N__7001),
            .I(N__6995));
    Span12Mux_h I__1247 (
            .O(N__6998),
            .I(N__6992));
    Span12Mux_h I__1246 (
            .O(N__6995),
            .I(N__6989));
    Span12Mux_v I__1245 (
            .O(N__6992),
            .I(N__6986));
    Odrv12 I__1244 (
            .O(N__6989),
            .I(TSn_c));
    Odrv12 I__1243 (
            .O(N__6986),
            .I(TSn_c));
    CascadeMux I__1242 (
            .O(N__6981),
            .I(\U712_CHIP_RAM.N_458_cascade_ ));
    InMux I__1241 (
            .O(N__6978),
            .I(N__6975));
    LocalMux I__1240 (
            .O(N__6975),
            .I(N__6972));
    Span4Mux_v I__1239 (
            .O(N__6972),
            .I(N__6969));
    Sp12to4 I__1238 (
            .O(N__6969),
            .I(N__6965));
    IoInMux I__1237 (
            .O(N__6968),
            .I(N__6962));
    Span12Mux_h I__1236 (
            .O(N__6965),
            .I(N__6959));
    LocalMux I__1235 (
            .O(N__6962),
            .I(N__6956));
    Span12Mux_v I__1234 (
            .O(N__6959),
            .I(N__6953));
    IoSpan4Mux I__1233 (
            .O(N__6956),
            .I(N__6950));
    Odrv12 I__1232 (
            .O(N__6953),
            .I(RAMENn_c));
    Odrv4 I__1231 (
            .O(N__6950),
            .I(RAMENn_c));
    CascadeMux I__1230 (
            .O(N__6945),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_1_cascade_ ));
    CascadeMux I__1229 (
            .O(N__6942),
            .I(N__6936));
    InMux I__1228 (
            .O(N__6941),
            .I(N__6933));
    InMux I__1227 (
            .O(N__6940),
            .I(N__6926));
    InMux I__1226 (
            .O(N__6939),
            .I(N__6926));
    InMux I__1225 (
            .O(N__6936),
            .I(N__6926));
    LocalMux I__1224 (
            .O(N__6933),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    LocalMux I__1223 (
            .O(N__6926),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    CascadeMux I__1222 (
            .O(N__6921),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0_0_cascade_ ));
    InMux I__1221 (
            .O(N__6918),
            .I(N__6915));
    LocalMux I__1220 (
            .O(N__6915),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0 ));
    IoInMux I__1219 (
            .O(N__6912),
            .I(N__6909));
    LocalMux I__1218 (
            .O(N__6909),
            .I(N__6906));
    Span4Mux_s1_h I__1217 (
            .O(N__6906),
            .I(N__6903));
    Sp12to4 I__1216 (
            .O(N__6903),
            .I(N__6900));
    Span12Mux_s11_v I__1215 (
            .O(N__6900),
            .I(N__6897));
    Odrv12 I__1214 (
            .O(N__6897),
            .I(CLK_EN_c));
    CEMux I__1213 (
            .O(N__6894),
            .I(N__6891));
    LocalMux I__1212 (
            .O(N__6891),
            .I(N__6888));
    Odrv12 I__1211 (
            .O(N__6888),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0 ));
    CascadeMux I__1210 (
            .O(N__6885),
            .I(\U712_CHIP_RAM.N_344_cascade_ ));
    InMux I__1209 (
            .O(N__6882),
            .I(N__6879));
    LocalMux I__1208 (
            .O(N__6879),
            .I(\U712_CHIP_RAM.N_435 ));
    InMux I__1207 (
            .O(N__6876),
            .I(N__6870));
    InMux I__1206 (
            .O(N__6875),
            .I(N__6870));
    LocalMux I__1205 (
            .O(N__6870),
            .I(N__6867));
    Odrv4 I__1204 (
            .O(N__6867),
            .I(\U712_CHIP_RAM.N_430 ));
    InMux I__1203 (
            .O(N__6864),
            .I(N__6861));
    LocalMux I__1202 (
            .O(N__6861),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1 ));
    CascadeMux I__1201 (
            .O(N__6858),
            .I(N__6855));
    InMux I__1200 (
            .O(N__6855),
            .I(N__6840));
    InMux I__1199 (
            .O(N__6854),
            .I(N__6840));
    InMux I__1198 (
            .O(N__6853),
            .I(N__6840));
    InMux I__1197 (
            .O(N__6852),
            .I(N__6840));
    InMux I__1196 (
            .O(N__6851),
            .I(N__6836));
    InMux I__1195 (
            .O(N__6850),
            .I(N__6831));
    InMux I__1194 (
            .O(N__6849),
            .I(N__6831));
    LocalMux I__1193 (
            .O(N__6840),
            .I(N__6828));
    InMux I__1192 (
            .O(N__6839),
            .I(N__6825));
    LocalMux I__1191 (
            .O(N__6836),
            .I(N__6822));
    LocalMux I__1190 (
            .O(N__6831),
            .I(N__6818));
    Span4Mux_h I__1189 (
            .O(N__6828),
            .I(N__6813));
    LocalMux I__1188 (
            .O(N__6825),
            .I(N__6813));
    Span12Mux_h I__1187 (
            .O(N__6822),
            .I(N__6810));
    InMux I__1186 (
            .O(N__6821),
            .I(N__6807));
    Span4Mux_h I__1185 (
            .O(N__6818),
            .I(N__6802));
    Span4Mux_h I__1184 (
            .O(N__6813),
            .I(N__6802));
    Odrv12 I__1183 (
            .O(N__6810),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__1182 (
            .O(N__6807),
            .I(DBR_SYNCZ0Z_1));
    Odrv4 I__1181 (
            .O(N__6802),
            .I(DBR_SYNCZ0Z_1));
    InMux I__1180 (
            .O(N__6795),
            .I(N__6789));
    InMux I__1179 (
            .O(N__6794),
            .I(N__6789));
    LocalMux I__1178 (
            .O(N__6789),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ0Z_1 ));
    CascadeMux I__1177 (
            .O(N__6786),
            .I(N__6783));
    InMux I__1176 (
            .O(N__6783),
            .I(N__6780));
    LocalMux I__1175 (
            .O(N__6780),
            .I(\U712_CHIP_RAM.N_362 ));
    CascadeMux I__1174 (
            .O(N__6777),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_165_i_i_0_cascade_ ));
    InMux I__1173 (
            .O(N__6774),
            .I(N__6770));
    InMux I__1172 (
            .O(N__6773),
            .I(N__6767));
    LocalMux I__1171 (
            .O(N__6770),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_o2_0_0 ));
    LocalMux I__1170 (
            .O(N__6767),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_o2_0_0 ));
    InMux I__1169 (
            .O(N__6762),
            .I(N__6759));
    LocalMux I__1168 (
            .O(N__6759),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_a2_1_0 ));
    InMux I__1167 (
            .O(N__6756),
            .I(N__6753));
    LocalMux I__1166 (
            .O(N__6753),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER19 ));
    CascadeMux I__1165 (
            .O(N__6750),
            .I(N__6747));
    InMux I__1164 (
            .O(N__6747),
            .I(N__6743));
    InMux I__1163 (
            .O(N__6746),
            .I(N__6740));
    LocalMux I__1162 (
            .O(N__6743),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ));
    LocalMux I__1161 (
            .O(N__6740),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ));
    CascadeMux I__1160 (
            .O(N__6735),
            .I(N__6731));
    InMux I__1159 (
            .O(N__6734),
            .I(N__6728));
    InMux I__1158 (
            .O(N__6731),
            .I(N__6725));
    LocalMux I__1157 (
            .O(N__6728),
            .I(DBR_SYNC_i_1));
    LocalMux I__1156 (
            .O(N__6725),
            .I(DBR_SYNC_i_1));
    CascadeMux I__1155 (
            .O(N__6720),
            .I(N__6717));
    InMux I__1154 (
            .O(N__6717),
            .I(N__6714));
    LocalMux I__1153 (
            .O(N__6714),
            .I(N__6711));
    Odrv4 I__1152 (
            .O(N__6711),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0 ));
    InMux I__1151 (
            .O(N__6708),
            .I(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ));
    InMux I__1150 (
            .O(N__6705),
            .I(N__6701));
    InMux I__1149 (
            .O(N__6704),
            .I(N__6698));
    LocalMux I__1148 (
            .O(N__6701),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ));
    LocalMux I__1147 (
            .O(N__6698),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ));
    InMux I__1146 (
            .O(N__6693),
            .I(N__6690));
    LocalMux I__1145 (
            .O(N__6690),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2 ));
    InMux I__1144 (
            .O(N__6687),
            .I(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ));
    InMux I__1143 (
            .O(N__6684),
            .I(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_2 ));
    CascadeMux I__1142 (
            .O(N__6681),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3_cascade_ ));
    InMux I__1141 (
            .O(N__6678),
            .I(N__6674));
    InMux I__1140 (
            .O(N__6677),
            .I(N__6671));
    LocalMux I__1139 (
            .O(N__6674),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ));
    LocalMux I__1138 (
            .O(N__6671),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ));
    InMux I__1137 (
            .O(N__6666),
            .I(N__6663));
    LocalMux I__1136 (
            .O(N__6663),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3 ));
    CascadeMux I__1135 (
            .O(N__6660),
            .I(\U712_CHIP_RAM.N_451_cascade_ ));
    CEMux I__1134 (
            .O(N__6657),
            .I(N__6654));
    LocalMux I__1133 (
            .O(N__6654),
            .I(\U712_CHIP_RAM.N_452_0 ));
    InMux I__1132 (
            .O(N__6651),
            .I(N__6648));
    LocalMux I__1131 (
            .O(N__6648),
            .I(N__6644));
    InMux I__1130 (
            .O(N__6647),
            .I(N__6641));
    Odrv4 I__1129 (
            .O(N__6644),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_0_2 ));
    LocalMux I__1128 (
            .O(N__6641),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_0_2 ));
    CascadeMux I__1127 (
            .O(N__6636),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_1_cascade_ ));
    InMux I__1126 (
            .O(N__6633),
            .I(N__6630));
    LocalMux I__1125 (
            .O(N__6630),
            .I(N__6626));
    InMux I__1124 (
            .O(N__6629),
            .I(N__6623));
    Span4Mux_h I__1123 (
            .O(N__6626),
            .I(N__6620));
    LocalMux I__1122 (
            .O(N__6623),
            .I(\U712_REG_SM.N_406 ));
    Odrv4 I__1121 (
            .O(N__6620),
            .I(\U712_REG_SM.N_406 ));
    InMux I__1120 (
            .O(N__6615),
            .I(N__6612));
    LocalMux I__1119 (
            .O(N__6612),
            .I(N__6609));
    Span4Mux_h I__1118 (
            .O(N__6609),
            .I(N__6602));
    InMux I__1117 (
            .O(N__6608),
            .I(N__6597));
    InMux I__1116 (
            .O(N__6607),
            .I(N__6597));
    InMux I__1115 (
            .O(N__6606),
            .I(N__6592));
    InMux I__1114 (
            .O(N__6605),
            .I(N__6592));
    Odrv4 I__1113 (
            .O(N__6602),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_8 ));
    LocalMux I__1112 (
            .O(N__6597),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_8 ));
    LocalMux I__1111 (
            .O(N__6592),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_8 ));
    InMux I__1110 (
            .O(N__6585),
            .I(N__6578));
    CascadeMux I__1109 (
            .O(N__6584),
            .I(N__6574));
    InMux I__1108 (
            .O(N__6583),
            .I(N__6571));
    InMux I__1107 (
            .O(N__6582),
            .I(N__6568));
    InMux I__1106 (
            .O(N__6581),
            .I(N__6565));
    LocalMux I__1105 (
            .O(N__6578),
            .I(N__6562));
    InMux I__1104 (
            .O(N__6577),
            .I(N__6553));
    InMux I__1103 (
            .O(N__6574),
            .I(N__6553));
    LocalMux I__1102 (
            .O(N__6571),
            .I(N__6550));
    LocalMux I__1101 (
            .O(N__6568),
            .I(N__6545));
    LocalMux I__1100 (
            .O(N__6565),
            .I(N__6545));
    Span4Mux_h I__1099 (
            .O(N__6562),
            .I(N__6542));
    InMux I__1098 (
            .O(N__6561),
            .I(N__6535));
    InMux I__1097 (
            .O(N__6560),
            .I(N__6535));
    InMux I__1096 (
            .O(N__6559),
            .I(N__6535));
    InMux I__1095 (
            .O(N__6558),
            .I(N__6532));
    LocalMux I__1094 (
            .O(N__6553),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv12 I__1093 (
            .O(N__6550),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__1092 (
            .O(N__6545),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__1091 (
            .O(N__6542),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1090 (
            .O(N__6535),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1089 (
            .O(N__6532),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    CascadeMux I__1088 (
            .O(N__6519),
            .I(\U712_REG_SM.N_445_cascade_ ));
    InMux I__1087 (
            .O(N__6516),
            .I(N__6513));
    LocalMux I__1086 (
            .O(N__6513),
            .I(N__6510));
    Odrv4 I__1085 (
            .O(N__6510),
            .I(\U712_REG_SM.REG_CYCLE_5_iv_0_0 ));
    InMux I__1084 (
            .O(N__6507),
            .I(N__6504));
    LocalMux I__1083 (
            .O(N__6504),
            .I(\U712_BYTE_ENABLE.LMBE_0_i_o3_0_oZ0Z2 ));
    IoInMux I__1082 (
            .O(N__6501),
            .I(N__6498));
    LocalMux I__1081 (
            .O(N__6498),
            .I(N__6495));
    Span4Mux_s2_v I__1080 (
            .O(N__6495),
            .I(N__6492));
    Span4Mux_h I__1079 (
            .O(N__6492),
            .I(N__6489));
    Span4Mux_h I__1078 (
            .O(N__6489),
            .I(N__6486));
    Span4Mux_v I__1077 (
            .O(N__6486),
            .I(N__6483));
    Odrv4 I__1076 (
            .O(N__6483),
            .I(N_282_i));
    IoInMux I__1075 (
            .O(N__6480),
            .I(N__6477));
    LocalMux I__1074 (
            .O(N__6477),
            .I(N__6474));
    Span4Mux_s2_v I__1073 (
            .O(N__6474),
            .I(N__6471));
    Span4Mux_v I__1072 (
            .O(N__6471),
            .I(N__6468));
    Odrv4 I__1071 (
            .O(N__6468),
            .I(N_219));
    IoInMux I__1070 (
            .O(N__6465),
            .I(N__6462));
    LocalMux I__1069 (
            .O(N__6462),
            .I(N__6459));
    Span4Mux_s3_v I__1068 (
            .O(N__6459),
            .I(N__6456));
    Odrv4 I__1067 (
            .O(N__6456),
            .I(N_60_i));
    CascadeMux I__1066 (
            .O(N__6453),
            .I(\U712_CHIP_RAM.N_365_cascade_ ));
    CascadeMux I__1065 (
            .O(N__6450),
            .I(N__6446));
    InMux I__1064 (
            .O(N__6449),
            .I(N__6441));
    InMux I__1063 (
            .O(N__6446),
            .I(N__6441));
    LocalMux I__1062 (
            .O(N__6441),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ));
    CascadeMux I__1061 (
            .O(N__6438),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_ ));
    InMux I__1060 (
            .O(N__6435),
            .I(N__6432));
    LocalMux I__1059 (
            .O(N__6432),
            .I(N__6429));
    Span12Mux_h I__1058 (
            .O(N__6429),
            .I(N__6426));
    Span12Mux_v I__1057 (
            .O(N__6426),
            .I(N__6423));
    Odrv12 I__1056 (
            .O(N__6423),
            .I(A_c_2));
    InMux I__1055 (
            .O(N__6420),
            .I(N__6417));
    LocalMux I__1054 (
            .O(N__6417),
            .I(N__6414));
    Span12Mux_v I__1053 (
            .O(N__6414),
            .I(N__6411));
    Span12Mux_h I__1052 (
            .O(N__6411),
            .I(N__6408));
    Odrv12 I__1051 (
            .O(N__6408),
            .I(A_c_3));
    InMux I__1050 (
            .O(N__6405),
            .I(N__6402));
    LocalMux I__1049 (
            .O(N__6402),
            .I(N__6399));
    Odrv4 I__1048 (
            .O(N__6399),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ));
    InMux I__1047 (
            .O(N__6396),
            .I(N__6393));
    LocalMux I__1046 (
            .O(N__6393),
            .I(N__6390));
    Span12Mux_v I__1045 (
            .O(N__6390),
            .I(N__6387));
    Span12Mux_h I__1044 (
            .O(N__6387),
            .I(N__6384));
    Odrv12 I__1043 (
            .O(N__6384),
            .I(A_c_4));
    InMux I__1042 (
            .O(N__6381),
            .I(N__6378));
    LocalMux I__1041 (
            .O(N__6378),
            .I(N__6375));
    Span4Mux_v I__1040 (
            .O(N__6375),
            .I(N__6372));
    Sp12to4 I__1039 (
            .O(N__6372),
            .I(N__6369));
    Span12Mux_h I__1038 (
            .O(N__6369),
            .I(N__6366));
    Odrv12 I__1037 (
            .O(N__6366),
            .I(A_c_7));
    IoInMux I__1036 (
            .O(N__6363),
            .I(N__6360));
    LocalMux I__1035 (
            .O(N__6360),
            .I(N__6357));
    IoSpan4Mux I__1034 (
            .O(N__6357),
            .I(N__6354));
    Span4Mux_s0_v I__1033 (
            .O(N__6354),
            .I(N__6350));
    CascadeMux I__1032 (
            .O(N__6353),
            .I(N__6345));
    Sp12to4 I__1031 (
            .O(N__6350),
            .I(N__6342));
    InMux I__1030 (
            .O(N__6349),
            .I(N__6339));
    InMux I__1029 (
            .O(N__6348),
            .I(N__6334));
    InMux I__1028 (
            .O(N__6345),
            .I(N__6334));
    Span12Mux_v I__1027 (
            .O(N__6342),
            .I(N__6330));
    LocalMux I__1026 (
            .O(N__6339),
            .I(N__6327));
    LocalMux I__1025 (
            .O(N__6334),
            .I(N__6324));
    InMux I__1024 (
            .O(N__6333),
            .I(N__6321));
    Odrv12 I__1023 (
            .O(N__6330),
            .I(DBENn_c));
    Odrv4 I__1022 (
            .O(N__6327),
            .I(DBENn_c));
    Odrv4 I__1021 (
            .O(N__6324),
            .I(DBENn_c));
    LocalMux I__1020 (
            .O(N__6321),
            .I(DBENn_c));
    InMux I__1019 (
            .O(N__6312),
            .I(N__6309));
    LocalMux I__1018 (
            .O(N__6309),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_1Z0Z_0 ));
    CascadeMux I__1017 (
            .O(N__6306),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_1Z0Z_0_cascade_ ));
    IoInMux I__1016 (
            .O(N__6303),
            .I(N__6300));
    LocalMux I__1015 (
            .O(N__6300),
            .I(N__6297));
    Span4Mux_s2_h I__1014 (
            .O(N__6297),
            .I(N__6294));
    Sp12to4 I__1013 (
            .O(N__6294),
            .I(N__6291));
    Span12Mux_v I__1012 (
            .O(N__6291),
            .I(N__6288));
    Span12Mux_h I__1011 (
            .O(N__6288),
            .I(N__6285));
    Odrv12 I__1010 (
            .O(N__6285),
            .I(N_62_i));
    CascadeMux I__1009 (
            .O(N__6282),
            .I(\U712_CHIP_RAM.N_596_cascade_ ));
    InMux I__1008 (
            .O(N__6279),
            .I(N__6276));
    LocalMux I__1007 (
            .O(N__6276),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_0 ));
    CascadeMux I__1006 (
            .O(N__6273),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_ ));
    InMux I__1005 (
            .O(N__6270),
            .I(N__6266));
    InMux I__1004 (
            .O(N__6269),
            .I(N__6263));
    LocalMux I__1003 (
            .O(N__6266),
            .I(\U712_CHIP_RAM.N_596 ));
    LocalMux I__1002 (
            .O(N__6263),
            .I(\U712_CHIP_RAM.N_596 ));
    CascadeMux I__1001 (
            .O(N__6258),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_0_cascade_ ));
    InMux I__1000 (
            .O(N__6255),
            .I(N__6251));
    InMux I__999 (
            .O(N__6254),
            .I(N__6248));
    LocalMux I__998 (
            .O(N__6251),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0 ));
    LocalMux I__997 (
            .O(N__6248),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0 ));
    InMux I__996 (
            .O(N__6243),
            .I(N__6240));
    LocalMux I__995 (
            .O(N__6240),
            .I(N__6236));
    InMux I__994 (
            .O(N__6239),
            .I(N__6233));
    Span4Mux_v I__993 (
            .O(N__6236),
            .I(N__6229));
    LocalMux I__992 (
            .O(N__6233),
            .I(N__6226));
    InMux I__991 (
            .O(N__6232),
            .I(N__6223));
    Sp12to4 I__990 (
            .O(N__6229),
            .I(N__6220));
    Sp12to4 I__989 (
            .O(N__6226),
            .I(N__6215));
    LocalMux I__988 (
            .O(N__6223),
            .I(N__6215));
    Span12Mux_h I__987 (
            .O(N__6220),
            .I(N__6212));
    Span12Mux_h I__986 (
            .O(N__6215),
            .I(N__6209));
    Span12Mux_v I__985 (
            .O(N__6212),
            .I(N__6206));
    Span12Mux_v I__984 (
            .O(N__6209),
            .I(N__6203));
    Odrv12 I__983 (
            .O(N__6206),
            .I(AWEn_c));
    Odrv12 I__982 (
            .O(N__6203),
            .I(AWEn_c));
    InMux I__981 (
            .O(N__6198),
            .I(N__6194));
    InMux I__980 (
            .O(N__6197),
            .I(N__6191));
    LocalMux I__979 (
            .O(N__6194),
            .I(N__6188));
    LocalMux I__978 (
            .O(N__6191),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ));
    Odrv4 I__977 (
            .O(N__6188),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ));
    CascadeMux I__976 (
            .O(N__6183),
            .I(\U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_i_i_a2_0_cascade_ ));
    InMux I__975 (
            .O(N__6180),
            .I(N__6173));
    InMux I__974 (
            .O(N__6179),
            .I(N__6173));
    InMux I__973 (
            .O(N__6178),
            .I(N__6170));
    LocalMux I__972 (
            .O(N__6173),
            .I(N__6167));
    LocalMux I__971 (
            .O(N__6170),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    Odrv4 I__970 (
            .O(N__6167),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    InMux I__969 (
            .O(N__6162),
            .I(N__6159));
    LocalMux I__968 (
            .O(N__6159),
            .I(\U712_CHIP_RAM.N_365 ));
    SRMux I__967 (
            .O(N__6156),
            .I(N__6153));
    LocalMux I__966 (
            .O(N__6153),
            .I(N__6150));
    Span4Mux_h I__965 (
            .O(N__6150),
            .I(N__6146));
    InMux I__964 (
            .O(N__6149),
            .I(N__6143));
    Span4Mux_h I__963 (
            .O(N__6146),
            .I(N__6140));
    LocalMux I__962 (
            .O(N__6143),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    Odrv4 I__961 (
            .O(N__6140),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    CascadeMux I__960 (
            .O(N__6135),
            .I(\U712_CHIP_RAM.N_362_cascade_ ));
    CascadeMux I__959 (
            .O(N__6132),
            .I(\U712_CHIP_RAM.N_493_cascade_ ));
    CascadeMux I__958 (
            .O(N__6129),
            .I(\U712_CHIP_RAM.N_503_cascade_ ));
    InMux I__957 (
            .O(N__6126),
            .I(N__6123));
    LocalMux I__956 (
            .O(N__6123),
            .I(N__6120));
    Odrv12 I__955 (
            .O(N__6120),
            .I(\U712_REG_SM.N_482 ));
    InMux I__954 (
            .O(N__6117),
            .I(N__6113));
    IoInMux I__953 (
            .O(N__6116),
            .I(N__6110));
    LocalMux I__952 (
            .O(N__6113),
            .I(N__6107));
    LocalMux I__951 (
            .O(N__6110),
            .I(N__6104));
    Span12Mux_h I__950 (
            .O(N__6107),
            .I(N__6101));
    IoSpan4Mux I__949 (
            .O(N__6104),
            .I(N__6098));
    Span12Mux_h I__948 (
            .O(N__6101),
            .I(N__6095));
    IoSpan4Mux I__947 (
            .O(N__6098),
            .I(N__6092));
    Span12Mux_v I__946 (
            .O(N__6095),
            .I(N__6089));
    IoSpan4Mux I__945 (
            .O(N__6092),
            .I(N__6086));
    Odrv12 I__944 (
            .O(N__6089),
            .I(C1_c));
    Odrv4 I__943 (
            .O(N__6086),
            .I(C1_c));
    InMux I__942 (
            .O(N__6081),
            .I(N__6078));
    LocalMux I__941 (
            .O(N__6078),
            .I(N__6075));
    Odrv12 I__940 (
            .O(N__6075),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    InMux I__939 (
            .O(N__6072),
            .I(N__6069));
    LocalMux I__938 (
            .O(N__6069),
            .I(N__6066));
    Odrv4 I__937 (
            .O(N__6066),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ));
    IoInMux I__936 (
            .O(N__6063),
            .I(N__6060));
    LocalMux I__935 (
            .O(N__6060),
            .I(N__6057));
    Span4Mux_s2_h I__934 (
            .O(N__6057),
            .I(N__6054));
    Span4Mux_v I__933 (
            .O(N__6054),
            .I(N__6051));
    Sp12to4 I__932 (
            .O(N__6051),
            .I(N__6048));
    Span12Mux_h I__931 (
            .O(N__6048),
            .I(N__6045));
    Odrv12 I__930 (
            .O(N__6045),
            .I(CMA_c_6));
    InMux I__929 (
            .O(N__6042),
            .I(N__6039));
    LocalMux I__928 (
            .O(N__6039),
            .I(N__6036));
    Odrv4 I__927 (
            .O(N__6036),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ));
    IoInMux I__926 (
            .O(N__6033),
            .I(N__6030));
    LocalMux I__925 (
            .O(N__6030),
            .I(N__6027));
    Span4Mux_s3_h I__924 (
            .O(N__6027),
            .I(N__6024));
    Span4Mux_v I__923 (
            .O(N__6024),
            .I(N__6021));
    Sp12to4 I__922 (
            .O(N__6021),
            .I(N__6018));
    Span12Mux_h I__921 (
            .O(N__6018),
            .I(N__6015));
    Odrv12 I__920 (
            .O(N__6015),
            .I(CMA_c_7));
    InMux I__919 (
            .O(N__6012),
            .I(N__6009));
    LocalMux I__918 (
            .O(N__6009),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8 ));
    IoInMux I__917 (
            .O(N__6006),
            .I(N__6003));
    LocalMux I__916 (
            .O(N__6003),
            .I(N__6000));
    Span4Mux_s2_h I__915 (
            .O(N__6000),
            .I(N__5997));
    Sp12to4 I__914 (
            .O(N__5997),
            .I(N__5994));
    Span12Mux_s9_v I__913 (
            .O(N__5994),
            .I(N__5991));
    Span12Mux_h I__912 (
            .O(N__5991),
            .I(N__5988));
    Odrv12 I__911 (
            .O(N__5988),
            .I(CMA_c_8));
    InMux I__910 (
            .O(N__5985),
            .I(N__5982));
    LocalMux I__909 (
            .O(N__5982),
            .I(N__5979));
    Span4Mux_v I__908 (
            .O(N__5979),
            .I(N__5976));
    Odrv4 I__907 (
            .O(N__5976),
            .I(\U712_REG_SM.N_481 ));
    IoInMux I__906 (
            .O(N__5973),
            .I(N__5970));
    LocalMux I__905 (
            .O(N__5970),
            .I(N__5967));
    Span4Mux_s2_v I__904 (
            .O(N__5967),
            .I(N__5964));
    Sp12to4 I__903 (
            .O(N__5964),
            .I(N__5961));
    Span12Mux_h I__902 (
            .O(N__5961),
            .I(N__5958));
    Span12Mux_v I__901 (
            .O(N__5958),
            .I(N__5954));
    InMux I__900 (
            .O(N__5957),
            .I(N__5951));
    Odrv12 I__899 (
            .O(N__5954),
            .I(LDSn_c));
    LocalMux I__898 (
            .O(N__5951),
            .I(LDSn_c));
    CascadeMux I__897 (
            .O(N__5946),
            .I(N__5942));
    InMux I__896 (
            .O(N__5945),
            .I(N__5937));
    InMux I__895 (
            .O(N__5942),
            .I(N__5937));
    LocalMux I__894 (
            .O(N__5937),
            .I(\U712_REG_SM.N_185 ));
    IoInMux I__893 (
            .O(N__5934),
            .I(N__5931));
    LocalMux I__892 (
            .O(N__5931),
            .I(N__5928));
    IoSpan4Mux I__891 (
            .O(N__5928),
            .I(N__5925));
    Sp12to4 I__890 (
            .O(N__5925),
            .I(N__5922));
    Span12Mux_s6_v I__889 (
            .O(N__5922),
            .I(N__5919));
    Span12Mux_v I__888 (
            .O(N__5919),
            .I(N__5915));
    InMux I__887 (
            .O(N__5918),
            .I(N__5912));
    Odrv12 I__886 (
            .O(N__5915),
            .I(UDSn_c));
    LocalMux I__885 (
            .O(N__5912),
            .I(UDSn_c));
    CascadeMux I__884 (
            .O(N__5907),
            .I(N__5904));
    InMux I__883 (
            .O(N__5904),
            .I(N__5901));
    LocalMux I__882 (
            .O(N__5901),
            .I(N__5898));
    Odrv12 I__881 (
            .O(N__5898),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_0Z0Z_0 ));
    InMux I__880 (
            .O(N__5895),
            .I(N__5892));
    LocalMux I__879 (
            .O(N__5892),
            .I(N__5889));
    Odrv4 I__878 (
            .O(N__5889),
            .I(\U712_BYTE_ENABLE.N_468 ));
    IoInMux I__877 (
            .O(N__5886),
            .I(N__5883));
    LocalMux I__876 (
            .O(N__5883),
            .I(N__5880));
    IoSpan4Mux I__875 (
            .O(N__5880),
            .I(N__5877));
    Span4Mux_s1_h I__874 (
            .O(N__5877),
            .I(N__5874));
    Sp12to4 I__873 (
            .O(N__5874),
            .I(N__5871));
    Span12Mux_h I__872 (
            .O(N__5871),
            .I(N__5868));
    Span12Mux_v I__871 (
            .O(N__5868),
            .I(N__5865));
    Odrv12 I__870 (
            .O(N__5865),
            .I(N_65_i));
    InMux I__869 (
            .O(N__5862),
            .I(N__5855));
    InMux I__868 (
            .O(N__5861),
            .I(N__5855));
    CascadeMux I__867 (
            .O(N__5860),
            .I(N__5852));
    LocalMux I__866 (
            .O(N__5855),
            .I(N__5849));
    InMux I__865 (
            .O(N__5852),
            .I(N__5846));
    Span4Mux_v I__864 (
            .O(N__5849),
            .I(N__5843));
    LocalMux I__863 (
            .O(N__5846),
            .I(N__5840));
    Odrv4 I__862 (
            .O(N__5843),
            .I(\U712_BYTE_ENABLE.N_343_i ));
    Odrv4 I__861 (
            .O(N__5840),
            .I(\U712_BYTE_ENABLE.N_343_i ));
    CascadeMux I__860 (
            .O(N__5835),
            .I(\U712_BYTE_ENABLE.N_466_cascade_ ));
    IoInMux I__859 (
            .O(N__5832),
            .I(N__5829));
    LocalMux I__858 (
            .O(N__5829),
            .I(N__5826));
    Span12Mux_s3_h I__857 (
            .O(N__5826),
            .I(N__5823));
    Span12Mux_h I__856 (
            .O(N__5823),
            .I(N__5820));
    Odrv12 I__855 (
            .O(N__5820),
            .I(N_67_i));
    IoInMux I__854 (
            .O(N__5817),
            .I(N__5814));
    LocalMux I__853 (
            .O(N__5814),
            .I(N__5811));
    Span12Mux_s4_v I__852 (
            .O(N__5811),
            .I(N__5808));
    Span12Mux_h I__851 (
            .O(N__5808),
            .I(N__5805));
    Odrv12 I__850 (
            .O(N__5805),
            .I(ASn_c));
    CEMux I__849 (
            .O(N__5802),
            .I(N__5799));
    LocalMux I__848 (
            .O(N__5799),
            .I(N__5796));
    Odrv4 I__847 (
            .O(N__5796),
            .I(\U712_REG_SM.N_185_0 ));
    InMux I__846 (
            .O(N__5793),
            .I(N__5787));
    InMux I__845 (
            .O(N__5792),
            .I(N__5787));
    LocalMux I__844 (
            .O(N__5787),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_3 ));
    InMux I__843 (
            .O(N__5784),
            .I(N__5781));
    LocalMux I__842 (
            .O(N__5781),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_4 ));
    InMux I__841 (
            .O(N__5778),
            .I(N__5775));
    LocalMux I__840 (
            .O(N__5775),
            .I(N__5772));
    Sp12to4 I__839 (
            .O(N__5772),
            .I(N__5769));
    Span12Mux_v I__838 (
            .O(N__5769),
            .I(N__5766));
    Span12Mux_h I__837 (
            .O(N__5766),
            .I(N__5763));
    Odrv12 I__836 (
            .O(N__5763),
            .I(A_c_8));
    InMux I__835 (
            .O(N__5760),
            .I(N__5757));
    LocalMux I__834 (
            .O(N__5757),
            .I(N__5754));
    Odrv4 I__833 (
            .O(N__5754),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ));
    InMux I__832 (
            .O(N__5751),
            .I(N__5748));
    LocalMux I__831 (
            .O(N__5748),
            .I(N__5745));
    Sp12to4 I__830 (
            .O(N__5745),
            .I(N__5742));
    Span12Mux_v I__829 (
            .O(N__5742),
            .I(N__5739));
    Span12Mux_h I__828 (
            .O(N__5739),
            .I(N__5736));
    Odrv12 I__827 (
            .O(N__5736),
            .I(A_c_18));
    InMux I__826 (
            .O(N__5733),
            .I(N__5730));
    LocalMux I__825 (
            .O(N__5730),
            .I(N__5727));
    Odrv4 I__824 (
            .O(N__5727),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ));
    InMux I__823 (
            .O(N__5724),
            .I(N__5721));
    LocalMux I__822 (
            .O(N__5721),
            .I(N__5718));
    Sp12to4 I__821 (
            .O(N__5718),
            .I(N__5715));
    Span12Mux_v I__820 (
            .O(N__5715),
            .I(N__5712));
    Span12Mux_h I__819 (
            .O(N__5712),
            .I(N__5709));
    Odrv12 I__818 (
            .O(N__5709),
            .I(A_c_20));
    InMux I__817 (
            .O(N__5706),
            .I(N__5702));
    InMux I__816 (
            .O(N__5705),
            .I(N__5699));
    LocalMux I__815 (
            .O(N__5702),
            .I(N__5696));
    LocalMux I__814 (
            .O(N__5699),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ));
    Odrv4 I__813 (
            .O(N__5696),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ));
    InMux I__812 (
            .O(N__5691),
            .I(N__5688));
    LocalMux I__811 (
            .O(N__5688),
            .I(N__5685));
    Span4Mux_v I__810 (
            .O(N__5685),
            .I(N__5682));
    Span4Mux_v I__809 (
            .O(N__5682),
            .I(N__5679));
    Sp12to4 I__808 (
            .O(N__5679),
            .I(N__5676));
    Span12Mux_h I__807 (
            .O(N__5676),
            .I(N__5673));
    Odrv12 I__806 (
            .O(N__5673),
            .I(A_c_15));
    CascadeMux I__805 (
            .O(N__5670),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ));
    InMux I__804 (
            .O(N__5667),
            .I(N__5664));
    LocalMux I__803 (
            .O(N__5664),
            .I(N__5659));
    InMux I__802 (
            .O(N__5663),
            .I(N__5656));
    InMux I__801 (
            .O(N__5662),
            .I(N__5653));
    Span4Mux_h I__800 (
            .O(N__5659),
            .I(N__5645));
    LocalMux I__799 (
            .O(N__5656),
            .I(N__5640));
    LocalMux I__798 (
            .O(N__5653),
            .I(N__5640));
    InMux I__797 (
            .O(N__5652),
            .I(N__5635));
    InMux I__796 (
            .O(N__5651),
            .I(N__5635));
    InMux I__795 (
            .O(N__5650),
            .I(N__5628));
    InMux I__794 (
            .O(N__5649),
            .I(N__5628));
    InMux I__793 (
            .O(N__5648),
            .I(N__5628));
    Odrv4 I__792 (
            .O(N__5645),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__791 (
            .O(N__5640),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__790 (
            .O(N__5635),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__789 (
            .O(N__5628),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    InMux I__788 (
            .O(N__5619),
            .I(N__5616));
    LocalMux I__787 (
            .O(N__5616),
            .I(\U712_REG_SM.N_407 ));
    CascadeMux I__786 (
            .O(N__5613),
            .I(\U712_REG_SM.N_369_cascade_ ));
    InMux I__785 (
            .O(N__5610),
            .I(N__5606));
    InMux I__784 (
            .O(N__5609),
            .I(N__5603));
    LocalMux I__783 (
            .O(N__5606),
            .I(N__5600));
    LocalMux I__782 (
            .O(N__5603),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    Odrv4 I__781 (
            .O(N__5600),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    CEMux I__780 (
            .O(N__5595),
            .I(N__5592));
    LocalMux I__779 (
            .O(N__5592),
            .I(N__5589));
    Span4Mux_v I__778 (
            .O(N__5589),
            .I(N__5586));
    Odrv4 I__777 (
            .O(N__5586),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0 ));
    InMux I__776 (
            .O(N__5583),
            .I(N__5580));
    LocalMux I__775 (
            .O(N__5580),
            .I(N__5577));
    Span4Mux_v I__774 (
            .O(N__5577),
            .I(N__5574));
    Span4Mux_v I__773 (
            .O(N__5574),
            .I(N__5571));
    Sp12to4 I__772 (
            .O(N__5571),
            .I(N__5568));
    Span12Mux_h I__771 (
            .O(N__5568),
            .I(N__5565));
    Odrv12 I__770 (
            .O(N__5565),
            .I(A_c_17));
    InMux I__769 (
            .O(N__5562),
            .I(N__5559));
    LocalMux I__768 (
            .O(N__5559),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8 ));
    CascadeMux I__767 (
            .O(N__5556),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_cascade_ ));
    CascadeMux I__766 (
            .O(N__5553),
            .I(\U712_REG_SM.N_366_cascade_ ));
    InMux I__765 (
            .O(N__5550),
            .I(N__5544));
    InMux I__764 (
            .O(N__5549),
            .I(N__5544));
    LocalMux I__763 (
            .O(N__5544),
            .I(\U712_REG_SM.un1_STATE_COUNT_1_sqmuxa_0 ));
    InMux I__762 (
            .O(N__5541),
            .I(N__5538));
    LocalMux I__761 (
            .O(N__5538),
            .I(N__5534));
    ClkMux I__760 (
            .O(N__5537),
            .I(N__5531));
    Span4Mux_v I__759 (
            .O(N__5534),
            .I(N__5527));
    LocalMux I__758 (
            .O(N__5531),
            .I(N__5524));
    ClkMux I__757 (
            .O(N__5530),
            .I(N__5521));
    Span4Mux_v I__756 (
            .O(N__5527),
            .I(N__5514));
    Span4Mux_h I__755 (
            .O(N__5524),
            .I(N__5514));
    LocalMux I__754 (
            .O(N__5521),
            .I(N__5514));
    Span4Mux_v I__753 (
            .O(N__5514),
            .I(N__5511));
    Span4Mux_v I__752 (
            .O(N__5511),
            .I(N__5508));
    Odrv4 I__751 (
            .O(N__5508),
            .I(CLK40_PLL));
    IoInMux I__750 (
            .O(N__5505),
            .I(N__5501));
    IoInMux I__749 (
            .O(N__5504),
            .I(N__5498));
    LocalMux I__748 (
            .O(N__5501),
            .I(N__5495));
    LocalMux I__747 (
            .O(N__5498),
            .I(N__5492));
    Span4Mux_s0_v I__746 (
            .O(N__5495),
            .I(N__5489));
    Span4Mux_s3_v I__745 (
            .O(N__5492),
            .I(N__5486));
    Span4Mux_v I__744 (
            .O(N__5489),
            .I(N__5483));
    Span4Mux_h I__743 (
            .O(N__5486),
            .I(N__5480));
    Sp12to4 I__742 (
            .O(N__5483),
            .I(N__5476));
    Span4Mux_h I__741 (
            .O(N__5480),
            .I(N__5473));
    IoInMux I__740 (
            .O(N__5479),
            .I(N__5470));
    Span12Mux_s11_h I__739 (
            .O(N__5476),
            .I(N__5465));
    Sp12to4 I__738 (
            .O(N__5473),
            .I(N__5465));
    LocalMux I__737 (
            .O(N__5470),
            .I(N__5462));
    Span12Mux_v I__736 (
            .O(N__5465),
            .I(N__5457));
    Span12Mux_s8_h I__735 (
            .O(N__5462),
            .I(N__5457));
    Odrv12 I__734 (
            .O(N__5457),
            .I(CLK40_PLL_iso_i));
    CascadeMux I__733 (
            .O(N__5454),
            .I(N__5449));
    CascadeMux I__732 (
            .O(N__5453),
            .I(N__5446));
    CascadeMux I__731 (
            .O(N__5452),
            .I(N__5443));
    InMux I__730 (
            .O(N__5449),
            .I(N__5437));
    InMux I__729 (
            .O(N__5446),
            .I(N__5437));
    InMux I__728 (
            .O(N__5443),
            .I(N__5432));
    InMux I__727 (
            .O(N__5442),
            .I(N__5432));
    LocalMux I__726 (
            .O(N__5437),
            .I(\U712_REG_SM.WRITE_CYCLEZ0 ));
    LocalMux I__725 (
            .O(N__5432),
            .I(\U712_REG_SM.WRITE_CYCLEZ0 ));
    CascadeMux I__724 (
            .O(N__5427),
            .I(N__5424));
    InMux I__723 (
            .O(N__5424),
            .I(N__5421));
    LocalMux I__722 (
            .O(N__5421),
            .I(\U712_REG_SM.N_375 ));
    InMux I__721 (
            .O(N__5418),
            .I(N__5412));
    InMux I__720 (
            .O(N__5417),
            .I(N__5409));
    InMux I__719 (
            .O(N__5416),
            .I(N__5404));
    InMux I__718 (
            .O(N__5415),
            .I(N__5404));
    LocalMux I__717 (
            .O(N__5412),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    LocalMux I__716 (
            .O(N__5409),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    LocalMux I__715 (
            .O(N__5404),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    InMux I__714 (
            .O(N__5397),
            .I(N__5390));
    InMux I__713 (
            .O(N__5396),
            .I(N__5390));
    InMux I__712 (
            .O(N__5395),
            .I(N__5387));
    LocalMux I__711 (
            .O(N__5390),
            .I(N__5384));
    LocalMux I__710 (
            .O(N__5387),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    Odrv4 I__709 (
            .O(N__5384),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    InMux I__708 (
            .O(N__5379),
            .I(N__5373));
    InMux I__707 (
            .O(N__5378),
            .I(N__5373));
    LocalMux I__706 (
            .O(N__5373),
            .I(\U712_REG_SM.N_483 ));
    CascadeMux I__705 (
            .O(N__5370),
            .I(\U712_REG_SM.N_483_cascade_ ));
    InMux I__704 (
            .O(N__5367),
            .I(N__5363));
    InMux I__703 (
            .O(N__5366),
            .I(N__5360));
    LocalMux I__702 (
            .O(N__5363),
            .I(N__5356));
    LocalMux I__701 (
            .O(N__5360),
            .I(N__5353));
    InMux I__700 (
            .O(N__5359),
            .I(N__5350));
    Odrv12 I__699 (
            .O(N__5356),
            .I(\U712_REG_SM.N_367 ));
    Odrv4 I__698 (
            .O(N__5353),
            .I(\U712_REG_SM.N_367 ));
    LocalMux I__697 (
            .O(N__5350),
            .I(\U712_REG_SM.N_367 ));
    InMux I__696 (
            .O(N__5343),
            .I(N__5337));
    InMux I__695 (
            .O(N__5342),
            .I(N__5333));
    InMux I__694 (
            .O(N__5341),
            .I(N__5328));
    InMux I__693 (
            .O(N__5340),
            .I(N__5328));
    LocalMux I__692 (
            .O(N__5337),
            .I(N__5325));
    InMux I__691 (
            .O(N__5336),
            .I(N__5322));
    LocalMux I__690 (
            .O(N__5333),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__689 (
            .O(N__5328),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    Odrv12 I__688 (
            .O(N__5325),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__687 (
            .O(N__5322),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    InMux I__686 (
            .O(N__5313),
            .I(N__5307));
    InMux I__685 (
            .O(N__5312),
            .I(N__5304));
    InMux I__684 (
            .O(N__5311),
            .I(N__5299));
    InMux I__683 (
            .O(N__5310),
            .I(N__5299));
    LocalMux I__682 (
            .O(N__5307),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__681 (
            .O(N__5304),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__680 (
            .O(N__5299),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    InMux I__679 (
            .O(N__5292),
            .I(N__5285));
    InMux I__678 (
            .O(N__5291),
            .I(N__5280));
    InMux I__677 (
            .O(N__5290),
            .I(N__5280));
    InMux I__676 (
            .O(N__5289),
            .I(N__5275));
    InMux I__675 (
            .O(N__5288),
            .I(N__5275));
    LocalMux I__674 (
            .O(N__5285),
            .I(\U712_REG_SM.N_358 ));
    LocalMux I__673 (
            .O(N__5280),
            .I(\U712_REG_SM.N_358 ));
    LocalMux I__672 (
            .O(N__5275),
            .I(\U712_REG_SM.N_358 ));
    InMux I__671 (
            .O(N__5268),
            .I(N__5265));
    LocalMux I__670 (
            .O(N__5265),
            .I(\U712_REG_SM.N_592 ));
    IoInMux I__669 (
            .O(N__5262),
            .I(N__5258));
    IoInMux I__668 (
            .O(N__5261),
            .I(N__5254));
    LocalMux I__667 (
            .O(N__5258),
            .I(N__5251));
    IoInMux I__666 (
            .O(N__5257),
            .I(N__5248));
    LocalMux I__665 (
            .O(N__5254),
            .I(N__5245));
    IoSpan4Mux I__664 (
            .O(N__5251),
            .I(N__5242));
    LocalMux I__663 (
            .O(N__5248),
            .I(N__5239));
    Span4Mux_s2_h I__662 (
            .O(N__5245),
            .I(N__5236));
    Span4Mux_s2_v I__661 (
            .O(N__5242),
            .I(N__5233));
    Span4Mux_s2_v I__660 (
            .O(N__5239),
            .I(N__5230));
    Sp12to4 I__659 (
            .O(N__5236),
            .I(N__5226));
    Span4Mux_v I__658 (
            .O(N__5233),
            .I(N__5223));
    Span4Mux_v I__657 (
            .O(N__5230),
            .I(N__5220));
    InMux I__656 (
            .O(N__5229),
            .I(N__5216));
    Span12Mux_v I__655 (
            .O(N__5226),
            .I(N__5213));
    Sp12to4 I__654 (
            .O(N__5223),
            .I(N__5210));
    Sp12to4 I__653 (
            .O(N__5220),
            .I(N__5207));
    CascadeMux I__652 (
            .O(N__5219),
            .I(N__5204));
    LocalMux I__651 (
            .O(N__5216),
            .I(N__5201));
    Span12Mux_h I__650 (
            .O(N__5213),
            .I(N__5194));
    Span12Mux_h I__649 (
            .O(N__5210),
            .I(N__5194));
    Span12Mux_h I__648 (
            .O(N__5207),
            .I(N__5194));
    InMux I__647 (
            .O(N__5204),
            .I(N__5191));
    Span4Mux_v I__646 (
            .O(N__5201),
            .I(N__5188));
    Odrv12 I__645 (
            .O(N__5194),
            .I(TACK_EN));
    LocalMux I__644 (
            .O(N__5191),
            .I(TACK_EN));
    Odrv4 I__643 (
            .O(N__5188),
            .I(TACK_EN));
    SRMux I__642 (
            .O(N__5181),
            .I(N__5178));
    LocalMux I__641 (
            .O(N__5178),
            .I(N__5175));
    Span4Mux_h I__640 (
            .O(N__5175),
            .I(N__5172));
    Span4Mux_h I__639 (
            .O(N__5172),
            .I(N__5169));
    Odrv4 I__638 (
            .O(N__5169),
            .I(\U712_CYCLE_TERM.TACK_RST_0_i ));
    IoInMux I__637 (
            .O(N__5166),
            .I(N__5163));
    LocalMux I__636 (
            .O(N__5163),
            .I(N__5160));
    Span12Mux_s5_v I__635 (
            .O(N__5160),
            .I(N__5157));
    Odrv12 I__634 (
            .O(N__5157),
            .I(RESETn_c_i));
    CascadeMux I__633 (
            .O(N__5154),
            .I(\U712_REG_SM.N_185_cascade_ ));
    InMux I__632 (
            .O(N__5151),
            .I(N__5148));
    LocalMux I__631 (
            .O(N__5148),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_7 ));
    CascadeMux I__630 (
            .O(N__5145),
            .I(\U712_REG_SM.N_368_cascade_ ));
    InMux I__629 (
            .O(N__5142),
            .I(N__5139));
    LocalMux I__628 (
            .O(N__5139),
            .I(N__5136));
    Odrv4 I__627 (
            .O(N__5136),
            .I(\U712_CHIP_RAM.N_378 ));
    InMux I__626 (
            .O(N__5133),
            .I(N__5128));
    InMux I__625 (
            .O(N__5132),
            .I(N__5125));
    InMux I__624 (
            .O(N__5131),
            .I(N__5122));
    LocalMux I__623 (
            .O(N__5128),
            .I(\U712_REG_SM.N_441 ));
    LocalMux I__622 (
            .O(N__5125),
            .I(\U712_REG_SM.N_441 ));
    LocalMux I__621 (
            .O(N__5122),
            .I(\U712_REG_SM.N_441 ));
    CascadeMux I__620 (
            .O(N__5115),
            .I(\U712_REG_SM.N_358_cascade_ ));
    InMux I__619 (
            .O(N__5112),
            .I(N__5109));
    LocalMux I__618 (
            .O(N__5109),
            .I(\U712_REG_SM.N_368 ));
    CascadeMux I__617 (
            .O(N__5106),
            .I(N__5103));
    InMux I__616 (
            .O(N__5103),
            .I(N__5100));
    LocalMux I__615 (
            .O(N__5100),
            .I(\U712_REG_SM.N_366 ));
    IoInMux I__614 (
            .O(N__5097),
            .I(N__5094));
    LocalMux I__613 (
            .O(N__5094),
            .I(N__5091));
    Span12Mux_s7_v I__612 (
            .O(N__5091),
            .I(N__5088));
    Odrv12 I__611 (
            .O(N__5088),
            .I(CMA_c_1));
    InMux I__610 (
            .O(N__5085),
            .I(N__5081));
    InMux I__609 (
            .O(N__5084),
            .I(N__5078));
    LocalMux I__608 (
            .O(N__5081),
            .I(N__5075));
    LocalMux I__607 (
            .O(N__5078),
            .I(\U712_REG_SM.START_RSTZ0 ));
    Odrv4 I__606 (
            .O(N__5075),
            .I(\U712_REG_SM.START_RSTZ0 ));
    InMux I__605 (
            .O(N__5070),
            .I(N__5067));
    LocalMux I__604 (
            .O(N__5067),
            .I(N__5064));
    Span4Mux_v I__603 (
            .O(N__5064),
            .I(N__5061));
    Sp12to4 I__602 (
            .O(N__5061),
            .I(N__5058));
    Span12Mux_h I__601 (
            .O(N__5058),
            .I(N__5055));
    Odrv12 I__600 (
            .O(N__5055),
            .I(REGSPACEn_c));
    CascadeMux I__599 (
            .O(N__5052),
            .I(\U712_REG_SM.N_455_cascade_ ));
    IoInMux I__598 (
            .O(N__5049),
            .I(N__5046));
    LocalMux I__597 (
            .O(N__5046),
            .I(N__5043));
    Span4Mux_s0_v I__596 (
            .O(N__5043),
            .I(N__5040));
    Span4Mux_v I__595 (
            .O(N__5040),
            .I(N__5036));
    InMux I__594 (
            .O(N__5039),
            .I(N__5033));
    Span4Mux_v I__593 (
            .O(N__5036),
            .I(N__5030));
    LocalMux I__592 (
            .O(N__5033),
            .I(N__5027));
    Sp12to4 I__591 (
            .O(N__5030),
            .I(N__5024));
    Span4Mux_v I__590 (
            .O(N__5027),
            .I(N__5021));
    Span12Mux_h I__589 (
            .O(N__5024),
            .I(N__5018));
    Sp12to4 I__588 (
            .O(N__5021),
            .I(N__5015));
    Span12Mux_v I__587 (
            .O(N__5018),
            .I(N__5010));
    Span12Mux_h I__586 (
            .O(N__5015),
            .I(N__5010));
    Odrv12 I__585 (
            .O(N__5010),
            .I(A_c_10));
    InMux I__584 (
            .O(N__5007),
            .I(N__5004));
    LocalMux I__583 (
            .O(N__5004),
            .I(\U712_CHIP_RAM.N_387 ));
    InMux I__582 (
            .O(N__5001),
            .I(N__4997));
    InMux I__581 (
            .O(N__5000),
            .I(N__4994));
    LocalMux I__580 (
            .O(N__4997),
            .I(REG_TACK));
    LocalMux I__579 (
            .O(N__4994),
            .I(REG_TACK));
    IoInMux I__578 (
            .O(N__4989),
            .I(N__4986));
    LocalMux I__577 (
            .O(N__4986),
            .I(N__4983));
    Span4Mux_s2_v I__576 (
            .O(N__4983),
            .I(N__4980));
    Span4Mux_v I__575 (
            .O(N__4980),
            .I(N__4977));
    Span4Mux_h I__574 (
            .O(N__4977),
            .I(N__4974));
    Odrv4 I__573 (
            .O(N__4974),
            .I(VBENn_c));
    InMux I__572 (
            .O(N__4971),
            .I(N__4966));
    InMux I__571 (
            .O(N__4970),
            .I(N__4961));
    InMux I__570 (
            .O(N__4969),
            .I(N__4961));
    LocalMux I__569 (
            .O(N__4966),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__568 (
            .O(N__4961),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    CascadeMux I__567 (
            .O(N__4956),
            .I(N__4952));
    InMux I__566 (
            .O(N__4955),
            .I(N__4948));
    InMux I__565 (
            .O(N__4952),
            .I(N__4943));
    InMux I__564 (
            .O(N__4951),
            .I(N__4943));
    LocalMux I__563 (
            .O(N__4948),
            .I(N__4937));
    LocalMux I__562 (
            .O(N__4943),
            .I(N__4937));
    InMux I__561 (
            .O(N__4942),
            .I(N__4934));
    Span4Mux_v I__560 (
            .O(N__4937),
            .I(N__4931));
    LocalMux I__559 (
            .O(N__4934),
            .I(\U712_CYCLE_TERM.TACK_STARTZ0 ));
    Odrv4 I__558 (
            .O(N__4931),
            .I(\U712_CYCLE_TERM.TACK_STARTZ0 ));
    InMux I__557 (
            .O(N__4926),
            .I(N__4919));
    InMux I__556 (
            .O(N__4925),
            .I(N__4910));
    InMux I__555 (
            .O(N__4924),
            .I(N__4910));
    InMux I__554 (
            .O(N__4923),
            .I(N__4910));
    InMux I__553 (
            .O(N__4922),
            .I(N__4910));
    LocalMux I__552 (
            .O(N__4919),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__551 (
            .O(N__4910),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    CascadeMux I__550 (
            .O(N__4905),
            .I(\U712_CYCLE_TERM.N_36_0_cascade_ ));
    IoInMux I__549 (
            .O(N__4902),
            .I(N__4898));
    IoInMux I__548 (
            .O(N__4901),
            .I(N__4895));
    LocalMux I__547 (
            .O(N__4898),
            .I(N__4891));
    LocalMux I__546 (
            .O(N__4895),
            .I(N__4888));
    IoInMux I__545 (
            .O(N__4894),
            .I(N__4885));
    Span4Mux_s3_h I__544 (
            .O(N__4891),
            .I(N__4882));
    IoSpan4Mux I__543 (
            .O(N__4888),
            .I(N__4879));
    LocalMux I__542 (
            .O(N__4885),
            .I(N__4876));
    Sp12to4 I__541 (
            .O(N__4882),
            .I(N__4873));
    Span4Mux_s3_v I__540 (
            .O(N__4879),
            .I(N__4870));
    Span4Mux_s3_v I__539 (
            .O(N__4876),
            .I(N__4867));
    Span12Mux_v I__538 (
            .O(N__4873),
            .I(N__4864));
    Sp12to4 I__537 (
            .O(N__4870),
            .I(N__4861));
    Sp12to4 I__536 (
            .O(N__4867),
            .I(N__4858));
    Span12Mux_h I__535 (
            .O(N__4864),
            .I(N__4850));
    Span12Mux_h I__534 (
            .O(N__4861),
            .I(N__4850));
    Span12Mux_h I__533 (
            .O(N__4858),
            .I(N__4850));
    InMux I__532 (
            .O(N__4857),
            .I(N__4847));
    Odrv12 I__531 (
            .O(N__4850),
            .I(TACK_OUT));
    LocalMux I__530 (
            .O(N__4847),
            .I(TACK_OUT));
    InMux I__529 (
            .O(N__4842),
            .I(N__4839));
    LocalMux I__528 (
            .O(N__4839),
            .I(N__4836));
    Span4Mux_h I__527 (
            .O(N__4836),
            .I(N__4833));
    Sp12to4 I__526 (
            .O(N__4833),
            .I(N__4830));
    Span12Mux_v I__525 (
            .O(N__4830),
            .I(N__4827));
    Span12Mux_h I__524 (
            .O(N__4827),
            .I(N__4824));
    Odrv12 I__523 (
            .O(N__4824),
            .I(A_c_16));
    CascadeMux I__522 (
            .O(N__4821),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_ ));
    InMux I__521 (
            .O(N__4818),
            .I(N__4815));
    LocalMux I__520 (
            .O(N__4815),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_4 ));
    InMux I__519 (
            .O(N__4812),
            .I(N__4806));
    InMux I__518 (
            .O(N__4811),
            .I(N__4806));
    LocalMux I__517 (
            .O(N__4806),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_5 ));
    InMux I__516 (
            .O(N__4803),
            .I(N__4800));
    LocalMux I__515 (
            .O(N__4800),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_6 ));
    IoInMux I__514 (
            .O(N__4797),
            .I(N__4794));
    LocalMux I__513 (
            .O(N__4794),
            .I(N__4791));
    IoSpan4Mux I__512 (
            .O(N__4791),
            .I(N__4788));
    Span4Mux_s2_v I__511 (
            .O(N__4788),
            .I(N__4785));
    Span4Mux_v I__510 (
            .O(N__4785),
            .I(N__4782));
    Sp12to4 I__509 (
            .O(N__4782),
            .I(N__4779));
    Span12Mux_v I__508 (
            .O(N__4779),
            .I(N__4775));
    InMux I__507 (
            .O(N__4778),
            .I(N__4772));
    Odrv12 I__506 (
            .O(N__4775),
            .I(PRnW_c));
    LocalMux I__505 (
            .O(N__4772),
            .I(PRnW_c));
    InMux I__504 (
            .O(N__4767),
            .I(N__4764));
    LocalMux I__503 (
            .O(N__4764),
            .I(\U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1 ));
    IoInMux I__502 (
            .O(N__4761),
            .I(N__4757));
    IoInMux I__501 (
            .O(N__4760),
            .I(N__4754));
    LocalMux I__500 (
            .O(N__4757),
            .I(N__4751));
    LocalMux I__499 (
            .O(N__4754),
            .I(N__4748));
    IoSpan4Mux I__498 (
            .O(N__4751),
            .I(N__4745));
    Span12Mux_s4_v I__497 (
            .O(N__4748),
            .I(N__4742));
    Span4Mux_s3_v I__496 (
            .O(N__4745),
            .I(N__4739));
    Span12Mux_h I__495 (
            .O(N__4742),
            .I(N__4736));
    Sp12to4 I__494 (
            .O(N__4739),
            .I(N__4733));
    Span12Mux_v I__493 (
            .O(N__4736),
            .I(N__4727));
    Span12Mux_v I__492 (
            .O(N__4733),
            .I(N__4727));
    InMux I__491 (
            .O(N__4732),
            .I(N__4724));
    Odrv12 I__490 (
            .O(N__4727),
            .I(BLSn_c));
    LocalMux I__489 (
            .O(N__4724),
            .I(BLSn_c));
    IoInMux I__488 (
            .O(N__4719),
            .I(N__4716));
    LocalMux I__487 (
            .O(N__4716),
            .I(N__4713));
    IoSpan4Mux I__486 (
            .O(N__4713),
            .I(N__4710));
    Span4Mux_s3_v I__485 (
            .O(N__4710),
            .I(N__4707));
    Sp12to4 I__484 (
            .O(N__4707),
            .I(N__4704));
    Span12Mux_v I__483 (
            .O(N__4704),
            .I(N__4701));
    Odrv12 I__482 (
            .O(N__4701),
            .I(N_58_i));
    InMux I__481 (
            .O(N__4698),
            .I(N__4692));
    InMux I__480 (
            .O(N__4697),
            .I(N__4692));
    LocalMux I__479 (
            .O(N__4692),
            .I(\U712_BYTE_ENABLE.N_352 ));
    InMux I__478 (
            .O(N__4689),
            .I(N__4685));
    InMux I__477 (
            .O(N__4688),
            .I(N__4682));
    LocalMux I__476 (
            .O(N__4685),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__475 (
            .O(N__4682),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__474 (
            .O(N__4677),
            .I(N__4673));
    InMux I__473 (
            .O(N__4676),
            .I(N__4670));
    LocalMux I__472 (
            .O(N__4673),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    LocalMux I__471 (
            .O(N__4670),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    CascadeMux I__470 (
            .O(N__4665),
            .I(N__4661));
    InMux I__469 (
            .O(N__4664),
            .I(N__4658));
    InMux I__468 (
            .O(N__4661),
            .I(N__4655));
    LocalMux I__467 (
            .O(N__4658),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__466 (
            .O(N__4655),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__465 (
            .O(N__4650),
            .I(N__4646));
    InMux I__464 (
            .O(N__4649),
            .I(N__4643));
    LocalMux I__463 (
            .O(N__4646),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    LocalMux I__462 (
            .O(N__4643),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    IoInMux I__461 (
            .O(N__4638),
            .I(N__4635));
    LocalMux I__460 (
            .O(N__4635),
            .I(N__4632));
    Span12Mux_s0_v I__459 (
            .O(N__4632),
            .I(N__4629));
    Span12Mux_v I__458 (
            .O(N__4629),
            .I(N__4625));
    InMux I__457 (
            .O(N__4628),
            .I(N__4622));
    Odrv12 I__456 (
            .O(N__4625),
            .I(DBDIR_c));
    LocalMux I__455 (
            .O(N__4622),
            .I(DBDIR_c));
    InMux I__454 (
            .O(N__4617),
            .I(N__4614));
    LocalMux I__453 (
            .O(N__4614),
            .I(N__4611));
    Odrv4 I__452 (
            .O(N__4611),
            .I(DBR_SYNCZ0Z_0));
    InMux I__451 (
            .O(N__4608),
            .I(N__4605));
    LocalMux I__450 (
            .O(N__4605),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    InMux I__449 (
            .O(N__4602),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__448 (
            .O(N__4599),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    InMux I__447 (
            .O(N__4596),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__446 (
            .O(N__4593),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__445 (
            .O(N__4590),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__444 (
            .O(N__4587),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    ClkMux I__443 (
            .O(N__4584),
            .I(N__4563));
    ClkMux I__442 (
            .O(N__4583),
            .I(N__4563));
    ClkMux I__441 (
            .O(N__4582),
            .I(N__4563));
    ClkMux I__440 (
            .O(N__4581),
            .I(N__4563));
    ClkMux I__439 (
            .O(N__4580),
            .I(N__4563));
    ClkMux I__438 (
            .O(N__4579),
            .I(N__4563));
    ClkMux I__437 (
            .O(N__4578),
            .I(N__4563));
    GlobalMux I__436 (
            .O(N__4563),
            .I(N__4560));
    gio2CtrlBuf I__435 (
            .O(N__4560),
            .I(C1_c_g));
    InMux I__434 (
            .O(N__4557),
            .I(N__4553));
    InMux I__433 (
            .O(N__4556),
            .I(N__4550));
    LocalMux I__432 (
            .O(N__4553),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__431 (
            .O(N__4550),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__430 (
            .O(N__4545),
            .I(N__4541));
    InMux I__429 (
            .O(N__4544),
            .I(N__4538));
    LocalMux I__428 (
            .O(N__4541),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__427 (
            .O(N__4538),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    IoInMux I__426 (
            .O(N__4533),
            .I(N__4530));
    LocalMux I__425 (
            .O(N__4530),
            .I(N__4527));
    IoSpan4Mux I__424 (
            .O(N__4527),
            .I(N__4524));
    Span4Mux_s3_h I__423 (
            .O(N__4524),
            .I(N__4521));
    Span4Mux_h I__422 (
            .O(N__4521),
            .I(N__4517));
    InMux I__421 (
            .O(N__4520),
            .I(N__4514));
    Span4Mux_h I__420 (
            .O(N__4517),
            .I(N__4511));
    LocalMux I__419 (
            .O(N__4514),
            .I(N__4508));
    Span4Mux_h I__418 (
            .O(N__4511),
            .I(N__4505));
    Span4Mux_v I__417 (
            .O(N__4508),
            .I(N__4502));
    Sp12to4 I__416 (
            .O(N__4505),
            .I(N__4497));
    Sp12to4 I__415 (
            .O(N__4502),
            .I(N__4497));
    Span12Mux_h I__414 (
            .O(N__4497),
            .I(N__4494));
    Span12Mux_v I__413 (
            .O(N__4494),
            .I(N__4491));
    Odrv12 I__412 (
            .O(N__4491),
            .I(C3_c));
    InMux I__411 (
            .O(N__4488),
            .I(N__4485));
    LocalMux I__410 (
            .O(N__4485),
            .I(N__4481));
    InMux I__409 (
            .O(N__4484),
            .I(N__4478));
    Span4Mux_v I__408 (
            .O(N__4481),
            .I(N__4475));
    LocalMux I__407 (
            .O(N__4478),
            .I(N__4472));
    Sp12to4 I__406 (
            .O(N__4475),
            .I(N__4469));
    Span12Mux_h I__405 (
            .O(N__4472),
            .I(N__4466));
    Span12Mux_h I__404 (
            .O(N__4469),
            .I(N__4463));
    Span12Mux_v I__403 (
            .O(N__4466),
            .I(N__4460));
    Span12Mux_v I__402 (
            .O(N__4463),
            .I(N__4457));
    Odrv12 I__401 (
            .O(N__4460),
            .I(DBRn_c));
    Odrv12 I__400 (
            .O(N__4457),
            .I(DBRn_c));
    IoInMux I__399 (
            .O(N__4452),
            .I(N__4449));
    LocalMux I__398 (
            .O(N__4449),
            .I(N__4446));
    Span12Mux_s6_v I__397 (
            .O(N__4446),
            .I(N__4443));
    Odrv12 I__396 (
            .O(N__4443),
            .I(CLK80_PLL_i_i));
    CascadeMux I__395 (
            .O(N__4440),
            .I(DBRn_c_i_cascade_));
    IoInMux I__394 (
            .O(N__4437),
            .I(N__4434));
    LocalMux I__393 (
            .O(N__4434),
            .I(N__4431));
    Span12Mux_s3_h I__392 (
            .O(N__4431),
            .I(N__4428));
    Odrv12 I__391 (
            .O(N__4428),
            .I(DBRn_c_i_0));
    InMux I__390 (
            .O(N__4425),
            .I(N__4422));
    LocalMux I__389 (
            .O(N__4422),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__388 (
            .O(N__4419),
            .I(bfn_10_6_0_));
    InMux I__387 (
            .O(N__4416),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    IoInMux I__386 (
            .O(N__4413),
            .I(N__4410));
    LocalMux I__385 (
            .O(N__4410),
            .I(N__4407));
    IoSpan4Mux I__384 (
            .O(N__4407),
            .I(N__4404));
    Span4Mux_s2_v I__383 (
            .O(N__4404),
            .I(N__4401));
    Sp12to4 I__382 (
            .O(N__4401),
            .I(N__4398));
    Span12Mux_v I__381 (
            .O(N__4398),
            .I(N__4395));
    Odrv12 I__380 (
            .O(N__4395),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .I(N__4584));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .I(N__4582));
    INV \INVU712_CHIP_RAM.DMA_A1_nesrC  (
            .O(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .I(N__4580));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .I(N__4581));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .I(N__4579));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ),
            .I(N__4578));
    INV \INVU712_CYCLE_TERM.TACK_STATE_0C  (
            .O(\INVU712_CYCLE_TERM.TACK_STATE_0C_net ),
            .I(N__5530));
    INV \INVU712_CYCLE_TERM.TACK_ENC  (
            .O(\INVU712_CYCLE_TERM.TACK_ENC_net ),
            .I(N__5537));
    defparam IN_MUX_bfv_10_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_6_0_));
    defparam IN_MUX_bfv_16_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_6_0_));
    defparam IN_MUX_bfv_15_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_4_0_));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__6116),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__5166),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB DBRn_c_i_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__4437),
            .GLOBALBUFFEROUTPUT(DBRn_c_i_0_g));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__4533),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_7_1_3.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_7_1_3.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_7_1_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 CLKRAM_obuf_RNO_LC_7_1_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11742),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBRn_ibuf_RNIBAB_LC_7_11_2.C_ON=1'b0;
    defparam DBRn_ibuf_RNIBAB_LC_7_11_2.SEQ_MODE=4'b0000;
    defparam DBRn_ibuf_RNIBAB_LC_7_11_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 DBRn_ibuf_RNIBAB_LC_7_11_2 (
            .in0(N__4488),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DBRn_c_i),
            .ltout(DBRn_c_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_7_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_7_11_3 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_7_11_3  (
            .in0(N__11141),
            .in1(_gnd_net_),
            .in2(N__4440),
            .in3(_gnd_net_),
            .lcout(DBRn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_6_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_6_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_6_0  (
            .in0(_gnd_net_),
            .in1(N__4425),
            .in2(_gnd_net_),
            .in3(N__4419),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_10_6_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__4583),
            .ce(),
            .sr(N__6156));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_6_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_6_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_6_1  (
            .in0(_gnd_net_),
            .in1(N__4677),
            .in2(_gnd_net_),
            .in3(N__4416),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__4583),
            .ce(),
            .sr(N__6156));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_6_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_6_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_6_2  (
            .in0(_gnd_net_),
            .in1(N__4650),
            .in2(_gnd_net_),
            .in3(N__4602),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__4583),
            .ce(),
            .sr(N__6156));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_6_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_6_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_6_3  (
            .in0(_gnd_net_),
            .in1(N__4689),
            .in2(_gnd_net_),
            .in3(N__4599),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__4583),
            .ce(),
            .sr(N__6156));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_6_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_6_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_6_4  (
            .in0(_gnd_net_),
            .in1(N__4664),
            .in2(_gnd_net_),
            .in3(N__4596),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__4583),
            .ce(),
            .sr(N__6156));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_6_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_6_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_6_5  (
            .in0(_gnd_net_),
            .in1(N__4545),
            .in2(_gnd_net_),
            .in3(N__4593),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__4583),
            .ce(),
            .sr(N__6156));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_6_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_6_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_6_6  (
            .in0(_gnd_net_),
            .in1(N__4557),
            .in2(_gnd_net_),
            .in3(N__4590),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__4583),
            .ce(),
            .sr(N__6156));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_6_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_6_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_6_7  (
            .in0(_gnd_net_),
            .in1(N__9149),
            .in2(_gnd_net_),
            .in3(N__4587),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4583),
            .ce(),
            .sr(N__6156));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_7_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_7_2  (
            .in0(_gnd_net_),
            .in1(N__4556),
            .in2(_gnd_net_),
            .in3(N__4544),
            .lcout(\U712_CHIP_RAM.REFRESH5lto7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_0_LC_10_8_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_10_8_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_10_8_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_10_8_2  (
            .in0(N__4520),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11713),
            .ce(),
            .sr(N__11081));
    defparam DBR_SYNC_0_LC_10_9_0.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_10_9_0.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_10_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_0_LC_10_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4484),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11720),
            .ce(),
            .sr(N__11074));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_LC_10_10_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_LC_10_10_1 .LUT_INIT=16'b0100111100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_LC_10_10_1  (
            .in0(N__7825),
            .in1(N__4698),
            .in2(N__5860),
            .in3(N__10516),
            .lcout(\U712_BYTE_ENABLE.N_468 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_58_i_LC_10_10_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_58_i_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_58_i_LC_10_10_3 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U712_BYTE_ENABLE.N_58_i_LC_10_10_3  (
            .in0(N__7824),
            .in1(N__4697),
            .in2(N__5907),
            .in3(N__10515),
            .lcout(N_58_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_o2_LC_10_11_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_o2_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_o2_LC_10_11_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_o2_LC_10_11_3  (
            .in0(N__7730),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7561),
            .lcout(\U712_BYTE_ENABLE.N_352 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_x2_LC_10_12_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_x2_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_x2_LC_10_12_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_x2_LC_10_12_5  (
            .in0(N__7543),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7615),
            .lcout(\U712_BYTE_ENABLE.N_343_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_LC_11_5_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_11_5_0 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_11_5_0 .LUT_INIT=16'b0011000100110000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_LC_11_5_0  (
            .in0(N__4926),
            .in1(N__4971),
            .in2(N__5219),
            .in3(N__4955),
            .lcout(TACK_EN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CYCLE_TERM.TACK_ENC_net ),
            .ce(),
            .sr(N__11096));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_6_0 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_6_0  (
            .in0(N__4688),
            .in1(N__4676),
            .in2(N__4665),
            .in3(N__4649),
            .lcout(\U712_CHIP_RAM.REFRESH5lt7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBDIR_LC_11_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_11_7_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_11_7_0 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_11_7_0  (
            .in0(N__6232),
            .in1(N__4628),
            .in2(_gnd_net_),
            .in3(N__6198),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11701),
            .ce(),
            .sr(N__11082));
    defparam DBR_SYNC_1_LC_11_7_2.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_11_7_2.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_11_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_11_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4617),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11701),
            .ce(),
            .sr(N__11082));
    defparam \U712_REG_SM.C3_SYNC_1_LC_11_8_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_11_8_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_11_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4608),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11707),
            .ce(),
            .sr(N__11075));
    defparam \U712_REG_SM.STATE_COUNT_7_LC_11_9_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_7_LC_11_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_7_LC_11_9_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_7_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__12005),
            .in2(_gnd_net_),
            .in3(N__4803),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11714),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_5_LC_11_9_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_11_9_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_5_LC_11_9_1  (
            .in0(N__12003),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4818),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11714),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_9_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_9_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_11_9_3  (
            .in0(N__12002),
            .in1(N__5312),
            .in2(_gnd_net_),
            .in3(N__5292),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11714),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_2_LC_11_9_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_2_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_2_LC_11_9_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_2_LC_11_9_4  (
            .in0(N__4811),
            .in1(N__5417),
            .in2(_gnd_net_),
            .in3(N__5132),
            .lcout(\U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_6_LC_11_9_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_11_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_11_9_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_6_LC_11_9_5  (
            .in0(N__12004),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4812),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11714),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.PRnW_LC_11_10_0 .C_ON=1'b0;
    defparam \U712_REG_SM.PRnW_LC_11_10_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.PRnW_LC_11_10_0 .LUT_INIT=16'b1110111101000101;
    LogicCell40 \U712_REG_SM.PRnW_LC_11_10_0  (
            .in0(N__5550),
            .in1(N__5663),
            .in2(N__5453),
            .in3(N__4778),
            .lcout(PRnW_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11721),
            .ce(),
            .sr(N__11067));
    defparam \U712_REG_SM.WRITE_CYCLE_LC_11_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.WRITE_CYCLE_LC_11_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.WRITE_CYCLE_LC_11_10_2 .LUT_INIT=16'b0101010111110000;
    LogicCell40 \U712_REG_SM.WRITE_CYCLE_LC_11_10_2  (
            .in0(N__10955),
            .in1(_gnd_net_),
            .in2(N__5454),
            .in3(N__5379),
            .lcout(\U712_REG_SM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11721),
            .ce(),
            .sr(N__11067));
    defparam \U712_REG_SM.REG_TACK_LC_11_10_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_11_10_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_11_10_3  (
            .in0(N__5001),
            .in1(N__4767),
            .in2(N__5427),
            .in3(N__5268),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11721),
            .ce(),
            .sr(N__11067));
    defparam \U712_REG_SM.START_RST_LC_11_10_4 .C_ON=1'b0;
    defparam \U712_REG_SM.START_RST_LC_11_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.START_RST_LC_11_10_4 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \U712_REG_SM.START_RST_LC_11_10_4  (
            .in0(N__5084),
            .in1(N__5342),
            .in2(_gnd_net_),
            .in3(N__5378),
            .lcout(\U712_REG_SM.START_RSTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11721),
            .ce(),
            .sr(N__11067));
    defparam \U712_REG_SM.REGENn_LC_11_10_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_LC_11_10_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_LC_11_10_5 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \U712_REG_SM.REGENn_LC_11_10_5  (
            .in0(N__5291),
            .in1(N__4732),
            .in2(_gnd_net_),
            .in3(N__5549),
            .lcout(BLSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11721),
            .ce(),
            .sr(N__11067));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_11_10_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_11_10_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_11_10_6 .LUT_INIT=16'b1111111110001111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_11_10_6  (
            .in0(N__5418),
            .in1(N__5290),
            .in2(N__5106),
            .in3(N__5133),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11721),
            .ce(),
            .sr(N__11067));
    defparam \U712_CYCLE_TERM.TACK_START_LC_11_11_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_START_LC_11_11_5 .SEQ_MODE=4'b1010;
    defparam \U712_CYCLE_TERM.TACK_START_LC_11_11_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_CYCLE_TERM.TACK_START_LC_11_11_5  (
            .in0(N__5000),
            .in1(N__7194),
            .in2(_gnd_net_),
            .in3(N__4942),
            .lcout(\U712_CYCLE_TERM.TACK_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11726),
            .ce(),
            .sr(N__5181));
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_12_4_1 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_12_4_1 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_12_4_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a2_LC_12_4_1  (
            .in0(N__10499),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9381),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_12_5_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_12_5_1 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_12_5_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_12_5_1  (
            .in0(N__4924),
            .in1(N__11925),
            .in2(N__4956),
            .in3(N__4970),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CYCLE_TERM.TACK_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_12_5_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_12_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_12_5_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_12_5_2  (
            .in0(N__11926),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4923),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CYCLE_TERM.TACK_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_OUT_RNO_0_LC_12_5_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUT_RNO_0_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_OUT_RNO_0_LC_12_5_4 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUT_RNO_0_LC_12_5_4  (
            .in0(N__4969),
            .in1(N__4922),
            .in2(_gnd_net_),
            .in3(N__4951),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_36_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_OUT_LC_12_5_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUT_LC_12_5_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_OUT_LC_12_5_5 .LUT_INIT=16'b1011111110110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUT_LC_12_5_5  (
            .in0(N__4925),
            .in1(N__11924),
            .in2(N__4905),
            .in3(N__4857),
            .lcout(TACK_OUT),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CYCLE_TERM.TACK_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_12_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_12_5_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_12_5_6  (
            .in0(N__5733),
            .in1(N__4842),
            .in2(_gnd_net_),
            .in3(N__9835),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_12_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_12_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_12_5_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_12_5_7  (
            .in0(N__9836),
            .in1(N__10498),
            .in2(N__4821),
            .in3(N__9246),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_12_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_12_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_12_6_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_LC_12_6_0  (
            .in0(N__9026),
            .in1(N__8442),
            .in2(N__9108),
            .in3(N__7170),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11689),
            .ce(N__5595),
            .sr(N__11080));
    defparam \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_12_6_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_12_6_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_12_6_7  (
            .in0(N__5343),
            .in1(N__5609),
            .in2(_gnd_net_),
            .in3(N__5366),
            .lcout(\U712_REG_SM.N_407 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_7_7 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_12_7_7  (
            .in0(N__10305),
            .in1(N__5007),
            .in2(N__9852),
            .in3(N__5142),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11695),
            .ce(N__10084),
            .sr(N__11073));
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_12_8_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_12_8_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(N__5085),
            .in2(_gnd_net_),
            .in3(N__5395),
            .lcout(),
            .ltout(\U712_REG_SM.N_455_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_12_8_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_12_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_12_8_2 .LUT_INIT=16'b1111000100000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_12_8_2  (
            .in0(N__5070),
            .in1(N__7017),
            .in2(N__5052),
            .in3(N__11923),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11700),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_8_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_8_3  (
            .in0(N__5039),
            .in1(N__10476),
            .in2(_gnd_net_),
            .in3(N__9609),
            .lcout(\U712_CHIP_RAM.N_387 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNITI8N_2_LC_12_8_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNITI8N_2_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNITI8N_2_LC_12_8_4 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNITI8N_2_LC_12_8_4  (
            .in0(N__5652),
            .in1(N__5610),
            .in2(_gnd_net_),
            .in3(N__6821),
            .lcout(\U712_REG_SM.N_406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_12_8_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_12_8_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_12_8_7  (
            .in0(_gnd_net_),
            .in1(N__5651),
            .in2(_gnd_net_),
            .in3(N__6558),
            .lcout(\U712_REG_SM.N_367 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNI902R1_1_LC_12_9_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI902R1_1_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI902R1_1_LC_12_9_0 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI902R1_1_LC_12_9_0  (
            .in0(N__5336),
            .in1(N__5131),
            .in2(_gnd_net_),
            .in3(N__5359),
            .lcout(\U712_REG_SM.N_185 ),
            .ltout(\U712_REG_SM.N_185_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_ess_RNO_LC_12_9_1 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_12_9_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_REG_SM.ASn_ess_RNO_LC_12_9_1  (
            .in0(N__11139),
            .in1(_gnd_net_),
            .in2(N__5154),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.N_185_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_0_1_LC_12_9_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_0_1_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_0_1_LC_12_9_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI6FIN_0_1_LC_12_9_2  (
            .in0(N__6560),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5649),
            .lcout(\U712_REG_SM.N_368 ),
            .ltout(\U712_REG_SM.N_368_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_8_LC_12_9_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_8_LC_12_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_8_LC_12_9_3 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_8_LC_12_9_3  (
            .in0(N__11922),
            .in1(N__5151),
            .in2(N__5145),
            .in3(N__6606),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11706),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_9_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_9_4  (
            .in0(N__6405),
            .in1(N__10435),
            .in2(_gnd_net_),
            .in3(N__10689),
            .lcout(\U712_CHIP_RAM.N_378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIO3HT_8_LC_12_9_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIO3HT_8_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIO3HT_8_LC_12_9_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIO3HT_8_LC_12_9_5  (
            .in0(N__5648),
            .in1(N__6605),
            .in2(_gnd_net_),
            .in3(N__6559),
            .lcout(\U712_REG_SM.N_441 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_1_LC_12_9_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_1_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_1_LC_12_9_6 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI6FIN_1_1_LC_12_9_6  (
            .in0(N__6561),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5650),
            .lcout(\U712_REG_SM.N_358 ),
            .ltout(\U712_REG_SM.N_358_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_12_9_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_12_9_7 .LUT_INIT=16'b1000000010100000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_12_9_7  (
            .in0(N__11921),
            .in1(N__5313),
            .in2(N__5115),
            .in3(N__6629),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11706),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_RNO_1_LC_12_10_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_1_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_1_LC_12_10_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_1_LC_12_10_0  (
            .in0(N__5442),
            .in1(N__5112),
            .in2(N__9380),
            .in3(N__6608),
            .lcout(\U712_REG_SM.REG_CYCLE_5_iv_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_RNIT80J_LC_12_10_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNIT80J_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNIT80J_LC_12_10_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNIT80J_LC_12_10_1  (
            .in0(N__5415),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5396),
            .lcout(\U712_REG_SM.N_366 ),
            .ltout(\U712_REG_SM.N_366_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIE5HG1_1_LC_12_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIE5HG1_1_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIE5HG1_1_LC_12_10_2 .LUT_INIT=16'b1111111111010001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIE5HG1_1_LC_12_10_2  (
            .in0(N__5340),
            .in1(N__5662),
            .in2(N__5553),
            .in3(N__6585),
            .lcout(\U712_REG_SM.un1_STATE_COUNT_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLK40_PLL_derived_clock_RNIIOT_LC_12_10_3.C_ON=1'b0;
    defparam CLK40_PLL_derived_clock_RNIIOT_LC_12_10_3.SEQ_MODE=4'b0000;
    defparam CLK40_PLL_derived_clock_RNIIOT_LC_12_10_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLK40_PLL_derived_clock_RNIIOT_LC_12_10_3 (
            .in0(N__5541),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK40_PLL_iso_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_12_10_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_12_10_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_12_10_4  (
            .in0(N__5310),
            .in1(_gnd_net_),
            .in2(N__5452),
            .in3(N__6607),
            .lcout(\U712_REG_SM.N_375 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_RNI3OIA1_LC_12_10_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNI3OIA1_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNI3OIA1_LC_12_10_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNI3OIA1_LC_12_10_5  (
            .in0(N__5416),
            .in1(N__5397),
            .in2(_gnd_net_),
            .in3(N__5288),
            .lcout(\U712_REG_SM.N_483 ),
            .ltout(\U712_REG_SM.N_483_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_12_10_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_12_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_12_10_6 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_12_10_6  (
            .in0(N__5341),
            .in1(N__11920),
            .in2(N__5370),
            .in3(N__5367),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11712),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_12_10_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_12_10_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_1_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(N__5311),
            .in2(_gnd_net_),
            .in3(N__5289),
            .lcout(\U712_REG_SM.N_592 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_START_RNO_0_LC_12_11_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_START_RNO_0_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_START_RNO_0_LC_12_11_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U712_CYCLE_TERM.TACK_START_RNO_0_LC_12_11_7  (
            .in0(N__11846),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5229),
            .lcout(\U712_CYCLE_TERM.TACK_RST_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDSn_RNO_0_LC_12_12_2 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_12_12_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U712_REG_SM.LDSn_RNO_0_LC_12_12_2  (
            .in0(N__10959),
            .in1(N__7731),
            .in2(N__7559),
            .in3(N__7633),
            .lcout(\U712_REG_SM.N_481 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_13_0.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_13_0.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_13_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11975),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_13_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_13_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_13_5_1 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_13_5_1  (
            .in0(N__9770),
            .in1(N__5562),
            .in2(N__10518),
            .in3(N__7860),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_13_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_13_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_13_5_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_13_5_2  (
            .in0(N__5691),
            .in1(N__5760),
            .in2(_gnd_net_),
            .in3(N__9768),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_5_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_5_3  (
            .in0(N__9769),
            .in1(N__10484),
            .in2(N__5670),
            .in3(N__9600),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_13_5_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_13_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_13_5_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_13_5_5  (
            .in0(_gnd_net_),
            .in1(N__5667),
            .in2(_gnd_net_),
            .in3(N__6851),
            .lcout(),
            .ltout(\U712_REG_SM.N_369_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_13_5_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_13_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_13_5_6 .LUT_INIT=16'b0010000000100010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_13_5_6  (
            .in0(N__12001),
            .in1(N__5619),
            .in2(N__5613),
            .in3(N__6583),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11693),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_13_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_13_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_13_6_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_13_6_0  (
            .in0(N__6254),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11143),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_13_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_13_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_13_6_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_13_6_1  (
            .in0(N__5583),
            .in1(N__5706),
            .in2(_gnd_net_),
            .in3(N__9738),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_13_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_13_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_13_6_2 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_13_6_2  (
            .in0(N__9736),
            .in1(N__9970),
            .in2(N__9906),
            .in3(N__6149),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_CMA25_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_13_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_13_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_13_6_3 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_13_6_3  (
            .in0(N__11144),
            .in1(_gnd_net_),
            .in2(N__5556),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_CMA25_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_13_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_13_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_13_6_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_13_6_4  (
            .in0(N__8694),
            .in1(N__5784),
            .in2(_gnd_net_),
            .in3(N__5792),
            .lcout(\U712_CHIP_RAM.N_499 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNI8NM9_LC_13_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNI8NM9_LC_13_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNI8NM9_LC_13_6_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_RNI8NM9_LC_13_6_5  (
            .in0(_gnd_net_),
            .in1(N__10448),
            .in2(_gnd_net_),
            .in3(N__9737),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_13_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_13_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_13_6_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_3_LC_13_6_6  (
            .in0(N__11999),
            .in1(N__12051),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11696),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_13_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_13_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_13_6_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_4_LC_13_6_7  (
            .in0(N__5793),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12000),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11696),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_13_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_13_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_13_7_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_13_7_4  (
            .in0(N__5778),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11702),
            .ce(N__8826),
            .sr(N__11083));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_13_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_13_7_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_13_7_7  (
            .in0(N__5751),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11702),
            .ce(N__8826),
            .sr(N__11083));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_13_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_13_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_13_8_0 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_13_8_0  (
            .in0(N__5724),
            .in1(N__11400),
            .in2(N__6450),
            .in3(N__5705),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11708),
            .ce(),
            .sr(N__11076));
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_13_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_13_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_13_8_1 .LUT_INIT=16'b1101110011111100;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_LC_13_8_1  (
            .in0(N__6162),
            .in1(N__6449),
            .in2(N__10485),
            .in3(N__6270),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11708),
            .ce(),
            .sr(N__11076));
    defparam \U712_CHIP_RAM.DBENn_LC_13_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_13_8_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_13_8_3 .LUT_INIT=16'b0100111011101110;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_13_8_3  (
            .in0(N__6255),
            .in1(N__6333),
            .in2(N__7032),
            .in3(N__9444),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11708),
            .ce(),
            .sr(N__11076));
    defparam \U712_REG_SM.LDSn_LC_13_8_4 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_LC_13_8_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.LDSn_LC_13_8_4 .LUT_INIT=16'b1111101011001100;
    LogicCell40 \U712_REG_SM.LDSn_LC_13_8_4  (
            .in0(N__5985),
            .in1(N__5957),
            .in2(N__6584),
            .in3(N__5945),
            .lcout(LDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11708),
            .ce(),
            .sr(N__11076));
    defparam \U712_REG_SM.UDSn_LC_13_8_5 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_LC_13_8_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.UDSn_LC_13_8_5 .LUT_INIT=16'b1111101011001010;
    LogicCell40 \U712_REG_SM.UDSn_LC_13_8_5  (
            .in0(N__5918),
            .in1(N__6577),
            .in2(N__5946),
            .in3(N__6126),
            .lcout(UDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11708),
            .ce(),
            .sr(N__11076));
    defparam \U712_REG_SM.C1_SYNC_1_LC_13_8_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_13_8_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_13_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_13_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6081),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11708),
            .ce(),
            .sr(N__11076));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_13_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_13_9_0 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_13_9_0  (
            .in0(N__6243),
            .in1(N__10963),
            .in2(_gnd_net_),
            .in3(N__9027),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11715),
            .ce(N__6657),
            .sr(N__11068));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_0_LC_13_10_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_0_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_0_LC_13_10_1 .LUT_INIT=16'b0011101100001010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_0_LC_13_10_1  (
            .in0(N__6312),
            .in1(N__5861),
            .in2(N__10782),
            .in3(N__10466),
            .lcout(\U712_BYTE_ENABLE.un1_CLLBEn_i_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_65_i_LC_13_10_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_65_i_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_65_i_LC_13_10_3 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \U712_BYTE_ENABLE.N_65_i_LC_13_10_3  (
            .in0(N__10778),
            .in1(N__5895),
            .in2(N__6353),
            .in3(N__8549),
            .lcout(N_65_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_13_10_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_13_10_5 .LUT_INIT=16'b0011011100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_13_10_5  (
            .in0(N__7827),
            .in1(N__5862),
            .in2(N__7752),
            .in3(N__10467),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_466_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_67_i_LC_13_10_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_67_i_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_67_i_LC_13_10_6 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \U712_BYTE_ENABLE.N_67_i_LC_13_10_6  (
            .in0(N__8550),
            .in1(N__6348),
            .in2(N__5835),
            .in3(N__10893),
            .lcout(N_67_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_ess_LC_13_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_LC_13_11_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_ess_LC_13_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.ASn_ess_LC_13_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6582),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11727),
            .ce(N__5802),
            .sr(N__11063));
    defparam \U712_REG_SM.UDSn_RNO_0_LC_13_12_1 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_RNO_0_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDSn_RNO_0_LC_13_12_1 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \U712_REG_SM.UDSn_RNO_0_LC_13_12_1  (
            .in0(N__7732),
            .in1(N__7634),
            .in2(N__7560),
            .in3(N__10965),
            .lcout(\U712_REG_SM.N_482 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_0_LC_13_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_13_13_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_13_13_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_13_13_4  (
            .in0(N__6117),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11735),
            .ce(),
            .sr(N__11062));
    defparam \U712_CHIP_RAM.CAS_COUNTER_0_LC_14_4_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_0_LC_14_4_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_0_LC_14_4_0 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_0_LC_14_4_0  (
            .in0(N__6850),
            .in1(N__11995),
            .in2(N__6720),
            .in3(N__8689),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11694),
            .ce(),
            .sr(_gnd_net_));
    defparam DBR_SYNC_RNITKK4_1_LC_14_4_2.C_ON=1'b0;
    defparam DBR_SYNC_RNITKK4_1_LC_14_4_2.SEQ_MODE=4'b0000;
    defparam DBR_SYNC_RNITKK4_1_LC_14_4_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 DBR_SYNC_RNITKK4_1_LC_14_4_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6839),
            .lcout(DBR_SYNC_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_2_LC_14_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_2_LC_14_4_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_2_LC_14_4_5 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_2_LC_14_4_5  (
            .in0(N__8690),
            .in1(N__6849),
            .in2(N__12006),
            .in3(N__6693),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11694),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_14_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_14_4_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_14_4_7 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_14_4_7  (
            .in0(N__8688),
            .in1(N__6704),
            .in2(N__6750),
            .in3(N__6677),
            .lcout(\U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_14_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_14_5_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_14_5_1 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_14_5_1  (
            .in0(N__10292),
            .in1(N__9573),
            .in2(N__10207),
            .in3(N__6072),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11697),
            .ce(N__10080),
            .sr(N__11102));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_14_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_14_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_14_5_2 .LUT_INIT=16'b1100010010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_14_5_2  (
            .in0(N__10194),
            .in1(N__10293),
            .in2(N__9489),
            .in3(N__6042),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11697),
            .ce(N__10080),
            .sr(N__11102));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_14_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_14_5_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_14_5_3 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_14_5_3  (
            .in0(N__10294),
            .in1(N__9261),
            .in2(N__10208),
            .in3(N__6012),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11697),
            .ce(N__10080),
            .sr(N__11102));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_14_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_14_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_14_5_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_14_5_6  (
            .in0(N__9730),
            .in1(N__10590),
            .in2(N__9959),
            .in3(N__9880),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMER12_LC_14_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMER12_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMER12_LC_14_6_0 .LUT_INIT=16'b0001010100110111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMER12_LC_14_6_0  (
            .in0(N__8402),
            .in1(N__8163),
            .in2(N__8235),
            .in3(N__8094),
            .lcout(\U712_CHIP_RAM.N_362 ),
            .ltout(\U712_CHIP_RAM.N_362_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_14_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_14_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_14_6_1 .LUT_INIT=16'b1010101010100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_14_6_1  (
            .in0(N__11991),
            .in1(N__8271),
            .in2(N__6135),
            .in3(N__6774),
            .lcout(\U712_CHIP_RAM.N_435 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_14_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_14_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_14_6_2 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_14_6_2  (
            .in0(N__8404),
            .in1(N__8099),
            .in2(N__7989),
            .in3(N__8965),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_493_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_14_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_14_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_14_6_3 .LUT_INIT=16'b1100110100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_14_6_3  (
            .in0(N__7053),
            .in1(N__6941),
            .in2(N__6132),
            .in3(N__9808),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11703),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_14_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_14_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_14_6_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_14_6_4  (
            .in0(_gnd_net_),
            .in1(N__11145),
            .in2(_gnd_net_),
            .in3(N__6279),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIBERN2_LC_14_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIBERN2_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIBERN2_LC_14_6_5 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNIBERN2_LC_14_6_5  (
            .in0(N__8164),
            .in1(N__8522),
            .in2(N__8112),
            .in3(N__7238),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_o2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_14_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_14_6_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_14_6_6  (
            .in0(N__8403),
            .in1(N__7100),
            .in2(N__7249),
            .in3(N__8098),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_14_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_14_7_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_14_7_0  (
            .in0(_gnd_net_),
            .in1(N__8166),
            .in2(_gnd_net_),
            .in3(N__7233),
            .lcout(\U712_CHIP_RAM.N_503 ),
            .ltout(\U712_CHIP_RAM.N_503_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_LC_14_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_LC_14_7_1 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_LC_14_7_1  (
            .in0(N__7101),
            .in1(_gnd_net_),
            .in2(N__6129),
            .in3(N__8084),
            .lcout(\U712_CHIP_RAM.N_596 ),
            .ltout(\U712_CHIP_RAM.N_596_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_14_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_14_7_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_14_7_2  (
            .in0(N__7141),
            .in1(N__8372),
            .in2(N__6282),
            .in3(N__6647),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_14_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_14_7_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_14_7_3  (
            .in0(N__9085),
            .in1(N__9018),
            .in2(N__8417),
            .in3(N__7139),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNILJ788_LC_14_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNILJ788_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNILJ788_LC_14_7_4 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNILJ788_LC_14_7_4  (
            .in0(N__7140),
            .in1(N__8027),
            .in2(N__6273),
            .in3(N__7102),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIMAOKC_LC_14_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIMAOKC_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIMAOKC_LC_14_7_5 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIMAOKC_LC_14_7_5  (
            .in0(N__8371),
            .in1(N__6269),
            .in2(N__6258),
            .in3(N__6180),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_14_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_14_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_14_7_6 .LUT_INIT=16'b0100010011000000;
    LogicCell40 \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_14_7_6  (
            .in0(N__6239),
            .in1(N__11976),
            .in2(N__10807),
            .in3(N__6197),
            .lcout(DMA_WRITE_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11709),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIVFJO_LC_14_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIVFJO_LC_14_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIVFJO_LC_14_7_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIVFJO_LC_14_7_7  (
            .in0(_gnd_net_),
            .in1(N__6179),
            .in2(_gnd_net_),
            .in3(N__8083),
            .lcout(\U712_CHIP_RAM.N_348 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_14_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_14_8_1 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_14_8_1  (
            .in0(N__7314),
            .in1(_gnd_net_),
            .in2(N__8401),
            .in3(N__9092),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_i_i_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_14_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_14_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_14_8_2 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_14_8_2  (
            .in0(N__8757),
            .in1(N__8004),
            .in2(N__6183),
            .in3(N__8970),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11716),
            .ce(N__9192),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1IJO_LC_14_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1IJO_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1IJO_LC_14_8_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1IJO_LC_14_8_3  (
            .in0(N__8346),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6178),
            .lcout(\U712_CHIP_RAM.N_365 ),
            .ltout(\U712_CHIP_RAM.N_365_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIIFS82_1_LC_14_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIIFS82_1_LC_14_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIIFS82_1_LC_14_8_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIIFS82_1_LC_14_8_4  (
            .in0(N__10389),
            .in1(N__8647),
            .in2(N__6453),
            .in3(N__7047),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIU7TF5_2_LC_14_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIU7TF5_2_LC_14_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIU7TF5_2_LC_14_8_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIU7TF5_2_LC_14_8_6  (
            .in0(N__7371),
            .in1(N__8347),
            .in2(N__9100),
            .in3(N__7145),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_2_LC_14_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_2_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_2_LC_14_8_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_2_LC_14_8_7  (
            .in0(N__11142),
            .in1(_gnd_net_),
            .in2(N__6438),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_14_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_14_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_14_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_14_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6435),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11722),
            .ce(N__8824),
            .sr(N__11077));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_14_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_14_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_14_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6420),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11722),
            .ce(N__8824),
            .sr(N__11077));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_14_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_14_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_14_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_14_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6396),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11722),
            .ce(N__8824),
            .sr(N__11077));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_14_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_14_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_14_9_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_14_9_3  (
            .in0(N__6381),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11722),
            .ce(N__8824),
            .sr(N__11077));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_1_0_LC_14_10_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_1_0_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_1_0_LC_14_10_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_1_0_LC_14_10_0  (
            .in0(N__6349),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8548),
            .lcout(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_1Z0Z_0 ),
            .ltout(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_62_i_LC_14_10_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_62_i_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_62_i_LC_14_10_1 .LUT_INIT=16'b0111011100000111;
    LogicCell40 \U712_BYTE_ENABLE.N_62_i_LC_14_10_1  (
            .in0(N__6507),
            .in1(N__10514),
            .in2(N__6306),
            .in3(N__10889),
            .lcout(N_62_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_14_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_14_10_3 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_14_10_3  (
            .in0(N__11140),
            .in1(N__7302),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_452_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_14_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_14_10_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_14_10_4  (
            .in0(N__8239),
            .in1(N__7984),
            .in2(N__8652),
            .in3(N__8423),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_14_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_14_10_5 .LUT_INIT=16'b1111110000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_14_10_5  (
            .in0(_gnd_net_),
            .in1(N__6651),
            .in2(N__6636),
            .in3(N__7158),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_14_10_6 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_14_10_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_0_LC_14_10_6  (
            .in0(N__6633),
            .in1(N__6615),
            .in2(_gnd_net_),
            .in3(N__6581),
            .lcout(),
            .ltout(\U712_REG_SM.N_445_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_14_10_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_14_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_14_10_7 .LUT_INIT=16'b1110111011100100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_14_10_7  (
            .in0(N__11930),
            .in1(N__9360),
            .in2(N__6519),
            .in3(N__6516),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11728),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LMBE_0_i_o3_0_o2_LC_14_11_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LMBE_0_i_o3_0_o2_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LMBE_0_i_o3_0_o2_LC_14_11_0 .LUT_INIT=16'b1111001000101111;
    LogicCell40 \U712_BYTE_ENABLE.LMBE_0_i_o3_0_o2_LC_14_11_0  (
            .in0(N__7826),
            .in1(N__7748),
            .in2(N__7659),
            .in3(N__7553),
            .lcout(\U712_BYTE_ENABLE.LMBE_0_i_o3_0_oZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.N_282_i_LC_14_20_0 .C_ON=1'b0;
    defparam \U712_BUFFERS.N_282_i_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.N_282_i_LC_14_20_0 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \U712_BUFFERS.N_282_i_LC_14_20_0  (
            .in0(N__10814),
            .in1(N__10869),
            .in2(_gnd_net_),
            .in3(N__10777),
            .lcout(N_282_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LLBE_0_i_o3_i_LC_14_20_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LLBE_0_i_o3_i_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LLBE_0_i_o3_i_LC_14_20_1 .LUT_INIT=16'b0000010101110000;
    LogicCell40 \U712_BYTE_ENABLE.LLBE_0_i_o3_i_LC_14_20_1  (
            .in0(N__7800),
            .in1(N__7736),
            .in2(N__7650),
            .in3(N__7535),
            .lcout(N_219),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_60_i_LC_14_20_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_60_i_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_60_i_LC_14_20_2 .LUT_INIT=16'b0101010010101000;
    LogicCell40 \U712_BYTE_ENABLE.N_60_i_LC_14_20_2  (
            .in0(N__7536),
            .in1(N__7801),
            .in2(N__7749),
            .in3(N__7641),
            .lcout(N_60_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_15_2_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_15_2_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_15_2_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_15_2_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_15_4_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_15_4_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_15_4_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_15_4_0  (
            .in0(_gnd_net_),
            .in1(N__6746),
            .in2(N__6735),
            .in3(N__6734),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_15_4_0_),
            .carryout(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_15_4_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_15_4_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_15_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_15_4_1  (
            .in0(_gnd_net_),
            .in1(N__6794),
            .in2(_gnd_net_),
            .in3(N__6708),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_15_4_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_15_4_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_15_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_15_4_2  (
            .in0(_gnd_net_),
            .in1(N__6705),
            .in2(_gnd_net_),
            .in3(N__6687),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_15_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_15_4_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_15_4_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_15_4_3  (
            .in0(_gnd_net_),
            .in1(N__6678),
            .in2(_gnd_net_),
            .in3(N__6684),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_3_LC_15_4_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_3_LC_15_4_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_3_LC_15_4_4 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_3_LC_15_4_4  (
            .in0(N__11993),
            .in1(N__6853),
            .in2(N__6681),
            .in3(N__8692),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11698),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_15_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_15_4_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_15_4_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_15_4_5  (
            .in0(N__6852),
            .in1(N__6666),
            .in2(_gnd_net_),
            .in3(N__6795),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_451_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_15_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_15_4_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_15_4_6 .LUT_INIT=16'b0000101000000010;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_15_4_6  (
            .in0(N__11994),
            .in1(N__6854),
            .in2(N__6660),
            .in3(N__8693),
            .lcout(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11698),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_1_LC_15_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_1_LC_15_4_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_1_LC_15_4_7 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_1_LC_15_4_7  (
            .in0(N__8691),
            .in1(N__6864),
            .in2(N__6858),
            .in3(N__11992),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11698),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4OVQ3_1_LC_15_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4OVQ3_1_LC_15_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4OVQ3_1_LC_15_5_0 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4OVQ3_1_LC_15_5_0  (
            .in0(N__6762),
            .in1(N__8616),
            .in2(N__6786),
            .in3(N__11990),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_165_i_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0MGF8_1_LC_15_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0MGF8_1_LC_15_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0MGF8_1_LC_15_5_1 .LUT_INIT=16'b0000010100001101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI0MGF8_1_LC_15_5_1  (
            .in0(N__11989),
            .in1(N__8264),
            .in2(N__6777),
            .in3(N__6773),
            .lcout(\U712_CHIP_RAM.N_132_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_15_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_15_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_15_5_2 .LUT_INIT=16'b1111000100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_15_5_2  (
            .in0(N__7377),
            .in1(N__6875),
            .in2(N__6942),
            .in3(N__9893),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11704),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_15_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_15_5_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_15_5_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_15_5_3  (
            .in0(N__8181),
            .in1(N__6940),
            .in2(_gnd_net_),
            .in3(N__10599),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11704),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_15_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_15_5_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_15_5_4 .LUT_INIT=16'b1010000010110001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_15_5_4  (
            .in0(N__6939),
            .in1(N__6876),
            .in2(N__9969),
            .in3(N__8253),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11704),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQ8AQ_LC_15_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQ8AQ_LC_15_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQ8AQ_LC_15_5_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQ8AQ_LC_15_5_5  (
            .in0(N__8400),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8161),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_a2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_15_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_15_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_15_5_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_15_5_6  (
            .in0(_gnd_net_),
            .in1(N__8615),
            .in2(_gnd_net_),
            .in3(N__7950),
            .lcout(\U712_CHIP_RAM.N_510 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_15_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_15_5_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_15_5_7 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_15_5_7  (
            .in0(N__11988),
            .in1(N__6756),
            .in2(_gnd_net_),
            .in3(N__8162),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11704),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI36AQC_2_LC_15_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI36AQC_2_LC_15_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI36AQC_2_LC_15_6_0 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI36AQC_2_LC_15_6_0  (
            .in0(N__8957),
            .in1(N__9101),
            .in2(N__8435),
            .in3(N__6918),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNINN3QI_LC_15_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNINN3QI_LC_15_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNINN3QI_LC_15_6_1 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNINN3QI_LC_15_6_1  (
            .in0(N__9017),
            .in1(N__8277),
            .in2(N__6945),
            .in3(N__8958),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_LC_15_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_LC_15_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_LC_15_6_2 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_LC_15_6_2  (
            .in0(N__8405),
            .in1(N__8626),
            .in2(N__8172),
            .in3(N__7046),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIEVI78_LC_15_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIEVI78_LC_15_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIEVI78_LC_15_6_3 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIEVI78_LC_15_6_3  (
            .in0(N__7088),
            .in1(N__8956),
            .in2(N__6921),
            .in3(N__8199),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_LC_15_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_LC_15_6_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_ess_LC_15_6_4 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_LC_15_6_4  (
            .in0(N__8409),
            .in1(N__7089),
            .in2(N__7248),
            .in3(N__8105),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11710),
            .ce(N__6894),
            .sr(N__11103));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_15_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_15_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_15_6_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_15_6_5  (
            .in0(N__11987),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7234),
            .lcout(\U712_CHIP_RAM.N_577 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_15_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_15_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_15_6_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_15_6_6  (
            .in0(N__8775),
            .in1(N__7907),
            .in2(N__8796),
            .in3(N__8705),
            .lcout(\U712_CHIP_RAM.N_344 ),
            .ltout(\U712_CHIP_RAM.N_344_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIR80N2_LC_15_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIR80N2_LC_15_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIR80N2_LC_15_6_7 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIR80N2_LC_15_6_7  (
            .in0(N__11986),
            .in1(_gnd_net_),
            .in2(N__6885),
            .in3(N__8167),
            .lcout(\U712_CHIP_RAM.N_508 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_15_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_15_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_15_7_2 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_15_7_2  (
            .in0(N__8568),
            .in1(N__6882),
            .in2(N__7392),
            .in3(N__8754),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11717),
            .ce(N__9181),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIF4EE6_2_LC_15_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIF4EE6_2_LC_15_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIF4EE6_2_LC_15_7_3 .LUT_INIT=16'b1010111000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIF4EE6_2_LC_15_7_3  (
            .in0(N__7062),
            .in1(N__9096),
            .in2(N__8426),
            .in3(N__8200),
            .lcout(\U712_CHIP_RAM.N_430 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_15_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_15_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_15_7_4 .LUT_INIT=16'b0000001001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_15_7_4  (
            .in0(N__8082),
            .in1(N__8622),
            .in2(N__7974),
            .in3(N__8384),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_347_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_0_LC_15_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_0_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_0_LC_15_7_5 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_0_LC_15_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7065),
            .in3(N__8171),
            .lcout(\U712_CHIP_RAM.N_590 ),
            .ltout(\U712_CHIP_RAM.N_590_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_15_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_15_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_15_7_6 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_15_7_6  (
            .in0(N__8201),
            .in1(_gnd_net_),
            .in2(N__7056),
            .in3(N__8919),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_3_LC_15_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_3_LC_15_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_3_LC_15_7_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_3_LC_15_7_7  (
            .in0(_gnd_net_),
            .in1(N__7957),
            .in2(_gnd_net_),
            .in3(N__8081),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_15_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_15_8_0 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_15_8_0  (
            .in0(N__9044),
            .in1(N__8485),
            .in2(N__8468),
            .in3(N__9010),
            .lcout(\U712_CHIP_RAM.N_350 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_3_LC_15_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_3_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_3_LC_15_8_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_3_LC_15_8_1  (
            .in0(N__8646),
            .in1(N__7970),
            .in2(_gnd_net_),
            .in3(N__8080),
            .lcout(\U712_CHIP_RAM.N_509 ),
            .ltout(\U712_CHIP_RAM.N_509_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_15_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_15_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_15_8_2 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNO_0_LC_15_8_2  (
            .in0(_gnd_net_),
            .in1(N__8430),
            .in2(N__7035),
            .in3(N__7250),
            .lcout(\U712_CHIP_RAM.DBENn_8_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_15_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_15_8_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_15_8_3  (
            .in0(N__8487),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10483),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_458_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_15_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_15_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_15_8_4 .LUT_INIT=16'b1010000010100010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_15_8_4  (
            .in0(N__11931),
            .in1(N__7013),
            .in2(N__6981),
            .in3(N__6978),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11723),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_0_LC_15_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_0_LC_15_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_0_LC_15_8_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_0_LC_15_8_6  (
            .in0(N__9045),
            .in1(N__8486),
            .in2(N__8469),
            .in3(N__9011),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_15_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_15_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_15_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_15_8_7  (
            .in0(N__7365),
            .in1(N__7349),
            .in2(_gnd_net_),
            .in3(N__9820),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_1_LC_15_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_1_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_1_LC_15_9_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_1_LC_15_9_0  (
            .in0(N__7313),
            .in1(N__9088),
            .in2(N__8434),
            .in3(N__7167),
            .lcout(\U712_CHIP_RAM.N_452 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_15_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_15_9_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_15_9_2  (
            .in0(N__7295),
            .in1(N__7260),
            .in2(_gnd_net_),
            .in3(N__9821),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_15_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_15_10_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_15_10_0  (
            .in0(N__8425),
            .in1(N__8113),
            .in2(N__7988),
            .in3(N__10510),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_15_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_15_10_1 .LUT_INIT=16'b0011001111110011;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(N__8651),
            .in2(N__7254),
            .in3(N__7251),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_72_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_15_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_15_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_15_10_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_15_10_2  (
            .in0(N__7187),
            .in1(N__7203),
            .in2(N__7197),
            .in3(N__7176),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11731),
            .ce(),
            .sr(N__11078));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1NGC4_2_LC_15_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1NGC4_2_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1NGC4_2_LC_15_10_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI1NGC4_2_LC_15_10_5  (
            .in0(N__7103),
            .in1(N__8424),
            .in2(N__8247),
            .in3(N__7168),
            .lcout(\U712_CHIP_RAM.N_462 ),
            .ltout(\U712_CHIP_RAM.N_462_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_15_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_15_10_6 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_15_10_6  (
            .in0(N__7169),
            .in1(N__8028),
            .in2(N__7107),
            .in3(N__7104),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_15_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_15_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_15_10_7 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_LC_15_10_7  (
            .in0(N__8114),
            .in1(N__8547),
            .in2(N__7896),
            .in3(N__7883),
            .lcout(LATCH_CLK_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11731),
            .ce(),
            .sr(N__11078));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_15_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_15_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_15_11_7 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_15_11_7  (
            .in0(N__7872),
            .in1(N__11304),
            .in2(N__10035),
            .in3(N__7853),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ),
            .ce(),
            .sr(N__11069));
    defparam \U712_BYTE_ENABLE.N_119_i_LC_15_20_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_119_i_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_119_i_LC_15_20_2 .LUT_INIT=16'b0000110111000000;
    LogicCell40 \U712_BYTE_ENABLE.N_119_i_LC_15_20_2  (
            .in0(N__7750),
            .in1(N__7802),
            .in2(N__7566),
            .in3(N__7651),
            .lcout(N_119_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_61_i_LC_15_20_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_61_i_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_61_i_LC_15_20_5 .LUT_INIT=16'b0000110111010000;
    LogicCell40 \U712_BYTE_ENABLE.N_61_i_LC_15_20_5  (
            .in0(N__7803),
            .in1(N__7751),
            .in2(N__7658),
            .in3(N__7565),
            .lcout(N_61_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_16_3_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_16_3_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_16_3_3 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_16_3_3  (
            .in0(N__10301),
            .in1(N__11508),
            .in2(N__10227),
            .in3(N__7422),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11699),
            .ce(N__10096),
            .sr(N__11113));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_16_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_16_4_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_16_4_6 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_16_4_6  (
            .in0(N__10529),
            .in1(N__7434),
            .in2(N__9851),
            .in3(N__10680),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_16_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_16_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_16_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_16_5_1  (
            .in0(N__8110),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7415),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_16_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_16_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_16_5_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_16_5_2  (
            .in0(N__8625),
            .in1(N__8438),
            .in2(N__8969),
            .in3(N__8111),
            .lcout(\U712_CHIP_RAM.N_431 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_16_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_16_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_16_5_3 .LUT_INIT=16'b1100110000010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_16_5_3  (
            .in0(N__8106),
            .in1(N__8623),
            .in2(_gnd_net_),
            .in3(N__7961),
            .lcout(\U712_CHIP_RAM.N_359 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIONRK3_1_LC_16_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIONRK3_1_LC_16_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIONRK3_1_LC_16_5_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIONRK3_1_LC_16_5_4  (
            .in0(N__8624),
            .in1(N__8437),
            .in2(_gnd_net_),
            .in3(N__8961),
            .lcout(\U712_CHIP_RAM.N_595 ),
            .ltout(\U712_CHIP_RAM.N_595_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_16_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_16_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_16_5_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_16_5_5  (
            .in0(N__8121),
            .in1(N__8243),
            .in2(N__8205),
            .in3(N__8202),
            .lcout(\U712_CHIP_RAM.N_279 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_16_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_16_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_16_5_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_16_5_7  (
            .in0(N__8436),
            .in1(N__8165),
            .in2(N__8115),
            .in3(N__7962),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_i_a2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI6FNG_LC_16_6_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI6FNG_LC_16_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI6FNG_LC_16_6_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNI6FNG_LC_16_6_0  (
            .in0(_gnd_net_),
            .in1(N__8079),
            .in2(_gnd_net_),
            .in3(N__8521),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_a2_0 ),
            .ltout(),
            .carryin(bfn_16_6_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_16_6_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_16_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_16_6_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_16_6_1  (
            .in0(N__8742),
            .in1(N__8627),
            .in2(_gnd_net_),
            .in3(N__8007),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(N__11718),
            .ce(N__9188),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_16_6_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_16_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_16_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_16_6_2  (
            .in0(_gnd_net_),
            .in1(N__8441),
            .in2(_gnd_net_),
            .in3(N__7992),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_16_6_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_16_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_16_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_16_6_3  (
            .in0(N__8743),
            .in1(N__7969),
            .in2(_gnd_net_),
            .in3(N__7911),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__11718),
            .ce(N__9188),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_16_6_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_16_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_16_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_16_6_4  (
            .in0(N__8755),
            .in1(N__7908),
            .in2(_gnd_net_),
            .in3(N__8799),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__11718),
            .ce(N__9188),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_16_6_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_16_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_16_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_16_6_5  (
            .in0(N__8744),
            .in1(N__8792),
            .in2(_gnd_net_),
            .in3(N__8778),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__11718),
            .ce(N__9188),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_16_6_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_16_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_16_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_16_6_6  (
            .in0(N__8756),
            .in1(N__8774),
            .in2(_gnd_net_),
            .in3(N__8760),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__11718),
            .ce(N__9188),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_16_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_16_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_16_6_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_16_6_7  (
            .in0(N__8745),
            .in1(N__8706),
            .in2(_gnd_net_),
            .in3(N__8709),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11718),
            .ce(N__9188),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_16_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_16_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_16_7_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_16_7_0  (
            .in0(N__11912),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9312),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11724),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_16_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_16_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_16_7_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_16_7_1  (
            .in0(N__8440),
            .in1(N__11919),
            .in2(_gnd_net_),
            .in3(N__8633),
            .lcout(\U712_CHIP_RAM.N_436 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_16_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_16_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_16_7_2 .LUT_INIT=16'b1010000011100000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_16_7_2  (
            .in0(N__8562),
            .in1(N__9016),
            .in2(N__11973),
            .in3(N__8541),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11724),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIHSKQ_LC_16_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIHSKQ_LC_16_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIHSKQ_LC_16_7_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIHSKQ_LC_16_7_3  (
            .in0(_gnd_net_),
            .in1(N__9042),
            .in2(_gnd_net_),
            .in3(N__8484),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_506_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNICG3P2_LC_16_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNICG3P2_LC_16_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNICG3P2_LC_16_7_4 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNICG3P2_LC_16_7_4  (
            .in0(N__8467),
            .in1(N__8439),
            .in2(N__8280),
            .in3(N__9086),
            .lcout(\U712_CHIP_RAM.N_147_i_i_a2_0 ),
            .ltout(\U712_CHIP_RAM.N_147_i_i_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_16_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_16_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_16_7_5 .LUT_INIT=16'b1010111111111111;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_16_7_5  (
            .in0(N__9015),
            .in1(_gnd_net_),
            .in2(N__9195),
            .in3(N__8960),
            .lcout(\U712_CHIP_RAM.N_500_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_16_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_16_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_16_7_6 .LUT_INIT=16'b1111000010110000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_16_7_6  (
            .in0(N__9156),
            .in1(N__9135),
            .in2(N__11974),
            .in3(N__9123),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11724),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_16_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_16_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_16_7_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_16_7_7  (
            .in0(N__9087),
            .in1(N__9043),
            .in2(N__9025),
            .in3(N__8959),
            .lcout(\U712_CHIP_RAM.N_494 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_16_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_16_8_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_16_8_1  (
            .in0(N__8913),
            .in1(N__9823),
            .in2(_gnd_net_),
            .in3(N__8859),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_16_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_16_8_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_16_8_2  (
            .in0(N__9822),
            .in1(N__8892),
            .in2(_gnd_net_),
            .in3(N__8832),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_16_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_16_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_16_8_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_16_8_3  (
            .in0(N__10468),
            .in1(N__9824),
            .in2(N__8877),
            .in3(N__12063),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_16_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_16_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_16_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_16_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8874),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11729),
            .ce(N__8825),
            .sr(N__11097));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_16_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_16_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_16_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_16_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8853),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11729),
            .ce(N__8825),
            .sr(N__11097));
    defparam \U712_BUFFERS.N_207_i_LC_16_9_0 .C_ON=1'b0;
    defparam \U712_BUFFERS.N_207_i_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.N_207_i_LC_16_9_0 .LUT_INIT=16'b0000000011111000;
    LogicCell40 \U712_BUFFERS.N_207_i_LC_16_9_0  (
            .in0(N__10881),
            .in1(N__10770),
            .in2(N__10517),
            .in3(N__9379),
            .lcout(N_207_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_16_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_16_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_16_9_2 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_16_9_2  (
            .in0(N__10882),
            .in1(N__11911),
            .in2(_gnd_net_),
            .in3(N__10771),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11732),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_16_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_16_9_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_16_9_6  (
            .in0(N__9303),
            .in1(_gnd_net_),
            .in2(N__9279),
            .in3(N__9825),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_16_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_16_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_16_9_7 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_16_9_7  (
            .in0(N__9267),
            .in1(N__10494),
            .in2(N__9848),
            .in3(N__10614),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_10_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_10_4  (
            .in0(N__9527),
            .in1(N__10030),
            .in2(_gnd_net_),
            .in3(N__11395),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11207),
            .ce(N__11176),
            .sr(N__11084));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_16_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_16_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_16_11_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_16_11_6  (
            .in0(N__10026),
            .in1(N__9528),
            .in2(_gnd_net_),
            .in3(N__11298),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .ce(N__11174),
            .sr(N__11079));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_17_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_17_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_17_7_7 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_17_7_7  (
            .in0(N__10290),
            .in1(N__9582),
            .in2(N__10228),
            .in3(N__9231),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11730),
            .ce(N__10098),
            .sr(N__11105));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_17_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_17_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_17_8_5 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_17_8_5  (
            .in0(N__10474),
            .in1(N__9207),
            .in2(N__9849),
            .in3(N__9588),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_17_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_17_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_17_8_7 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_17_8_7  (
            .in0(N__10475),
            .in1(N__9201),
            .in2(N__9850),
            .in3(N__10665),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_17_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_17_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_17_9_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_17_9_4  (
            .in0(N__9558),
            .in1(N__11394),
            .in2(_gnd_net_),
            .in3(N__9516),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .ce(N__11178),
            .sr(N__11098));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_17_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_17_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_17_9_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_17_9_6  (
            .in0(N__9557),
            .in1(N__11393),
            .in2(_gnd_net_),
            .in3(N__11448),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .ce(N__11178),
            .sr(N__11098));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_17_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_17_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_17_10_0 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_17_10_0  (
            .in0(N__10654),
            .in1(_gnd_net_),
            .in2(N__9474),
            .in3(N__11385),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11205),
            .ce(N__11177),
            .sr(N__11092));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_17_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_17_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_17_10_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_17_10_6  (
            .in0(N__11439),
            .in1(N__11386),
            .in2(_gnd_net_),
            .in3(N__9547),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11205),
            .ce(N__11177),
            .sr(N__11092));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_10_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_10_7  (
            .in0(N__9548),
            .in1(_gnd_net_),
            .in2(N__11396),
            .in3(N__9526),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11205),
            .ce(N__11177),
            .sr(N__11092));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_17_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_17_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_17_11_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_17_11_0  (
            .in0(N__11297),
            .in1(N__10653),
            .in2(_gnd_net_),
            .in3(N__9473),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__11175),
            .sr(N__11085));
    defparam \U712_CHIP_RAM.RASn_LC_18_2_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_18_2_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_18_2_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_18_2_0  (
            .in0(N__9905),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11705),
            .ce(),
            .sr(N__11118));
    defparam \U712_CHIP_RAM.CRCSn_LC_18_3_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_18_3_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_18_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_18_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9971),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11711),
            .ce(),
            .sr(N__11116));
    defparam \U712_CHIP_RAM.CASn_LC_18_3_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_18_3_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_18_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_18_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9847),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11711),
            .ce(),
            .sr(N__11116));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_18_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_18_4_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_18_4_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_18_4_7  (
            .in0(N__10266),
            .in1(N__9975),
            .in2(_gnd_net_),
            .in3(N__9846),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11719),
            .ce(N__10113),
            .sr(N__11115));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_18_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_18_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_18_5_3 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_18_5_3  (
            .in0(N__10601),
            .in1(N__9898),
            .in2(_gnd_net_),
            .in3(N__9845),
            .lcout(\U712_CHIP_RAM.CMA_5_i_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_18_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_18_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_18_5_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_18_5_6  (
            .in0(_gnd_net_),
            .in1(N__9897),
            .in2(_gnd_net_),
            .in3(N__10600),
            .lcout(\U712_CHIP_RAM.N_354 ),
            .ltout(\U712_CHIP_RAM.N_354_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_18_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_18_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_18_5_7 .LUT_INIT=16'b1110000011111111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_18_5_7  (
            .in0(N__10500),
            .in1(N__11232),
            .in2(N__9855),
            .in3(N__9844),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_18_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_18_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_18_6_7 .LUT_INIT=16'b0000100001010101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_18_6_7  (
            .in0(N__10265),
            .in1(N__11231),
            .in2(N__10528),
            .in3(N__9837),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_18_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_18_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_18_7_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_18_7_5  (
            .in0(N__9681),
            .in1(N__9672),
            .in2(_gnd_net_),
            .in3(N__9666),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11733),
            .ce(N__10108),
            .sr(N__11108));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_18_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_18_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_18_7_7 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_18_7_7  (
            .in0(N__10289),
            .in1(N__9615),
            .in2(N__10230),
            .in3(N__9639),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11733),
            .ce(N__10108),
            .sr(N__11108));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_18_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_18_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_18_8_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_18_8_0  (
            .in0(N__12105),
            .in1(N__11378),
            .in2(_gnd_net_),
            .in3(N__11585),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11208),
            .ce(N__11180),
            .sr(N__11106));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_18_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_18_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_18_8_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_18_8_4  (
            .in0(N__10659),
            .in1(N__11377),
            .in2(_gnd_net_),
            .in3(N__11543),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11208),
            .ce(N__11180),
            .sr(N__11106));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_18_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_18_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_18_9_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_18_9_2  (
            .in0(N__11542),
            .in1(_gnd_net_),
            .in2(N__11383),
            .in3(N__11583),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__11179),
            .sr(N__11104));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_18_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_18_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_18_9_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_18_9_3  (
            .in0(N__11584),
            .in1(N__11356),
            .in2(_gnd_net_),
            .in3(N__12102),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__11179),
            .sr(N__11104));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_18_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_18_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_18_9_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_18_9_4  (
            .in0(N__12103),
            .in1(_gnd_net_),
            .in2(N__11384),
            .in3(N__11495),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__11179),
            .sr(N__11104));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_18_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_18_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_18_9_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_18_9_5  (
            .in0(N__10658),
            .in1(N__11352),
            .in2(_gnd_net_),
            .in3(N__11541),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__11179),
            .sr(N__11104));
    defparam \U712_CHIP_RAM.WEn_LC_19_4_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_19_4_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_19_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_19_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10605),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11725),
            .ce(),
            .sr(N__11117));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_19_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_19_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_19_6_1 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_19_6_1  (
            .in0(N__10554),
            .in1(N__10548),
            .in2(N__10530),
            .in3(N__9984),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11734),
            .ce(N__10097),
            .sr(N__11114));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_19_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_19_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_19_7_7 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_19_7_7  (
            .in0(N__10291),
            .in1(N__12069),
            .in2(N__10229),
            .in3(N__10146),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11736),
            .ce(N__10112),
            .sr(N__11111));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_19_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_19_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_19_8_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_19_8_3  (
            .in0(N__11376),
            .in1(N__12035),
            .in2(_gnd_net_),
            .in3(N__10034),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11206),
            .ce(N__11182),
            .sr(N__11109));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_19_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_19_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_19_8_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_19_8_6  (
            .in0(N__11496),
            .in1(N__11375),
            .in2(_gnd_net_),
            .in3(N__12104),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11206),
            .ce(N__11182),
            .sr(N__11109));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_19_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_19_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_19_9_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_19_9_2  (
            .in0(N__11494),
            .in1(N__11351),
            .in2(_gnd_net_),
            .in3(N__11447),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__11181),
            .sr(N__11107));
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_20_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_20_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_20_6_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_2_LC_20_6_3  (
            .in0(_gnd_net_),
            .in1(N__11834),
            .in2(_gnd_net_),
            .in3(N__11748),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11737),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_20_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_20_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_20_7_3 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_0_LC_20_7_3  (
            .in0(N__12042),
            .in1(N__11832),
            .in2(_gnd_net_),
            .in3(N__12018),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11738),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_20_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_20_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_20_7_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_1_LC_20_7_7  (
            .in0(_gnd_net_),
            .in1(N__11833),
            .in2(_gnd_net_),
            .in3(N__11754),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11738),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_20_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_20_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_20_8_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_20_8_7  (
            .in0(N__11589),
            .in1(N__11379),
            .in2(_gnd_net_),
            .in3(N__11550),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11204),
            .ce(N__11184),
            .sr(N__11112));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_20_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_20_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_20_9_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_20_9_0  (
            .in0(N__11493),
            .in1(N__11440),
            .in2(_gnd_net_),
            .in3(N__11350),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11203),
            .ce(N__11183),
            .sr(N__11110));
    defparam \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_24_20_4 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_24_20_4 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_24_20_4 .LUT_INIT=16'b0100011100001111;
    LogicCell40 \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_24_20_4  (
            .in0(N__10964),
            .in1(N__10857),
            .in2(N__10821),
            .in3(N__10746),
            .lcout(N_409),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U712_TOP

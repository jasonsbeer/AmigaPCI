-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Apr 19 2025 16:01:24

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U111_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U111_TOP
entity U111_TOP is
port (
    D_UU_AMIGA : inout std_logic_vector(7 downto 0);
    D_LL_AMIGA : inout std_logic_vector(7 downto 0);
    D_UM_AMIGA : inout std_logic_vector(7 downto 0);
    D_LM_AMIGA : inout std_logic_vector(7 downto 0);
    D_UU_040 : inout std_logic_vector(7 downto 0);
    D_LM_040 : inout std_logic_vector(7 downto 0);
    D_UM_040 : inout std_logic_vector(7 downto 0);
    D_LL_040 : inout std_logic_vector(7 downto 0);
    A_AMIGA : out std_logic_vector(1 downto 0);
    A_040 : in std_logic_vector(1 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    TEAn : in std_logic;
    TSn : out std_logic;
    RESETn : in std_logic;
    CLKRAMA : out std_logic;
    PORTSIZE : in std_logic;
    TEA_CPUn : out std_logic;
    LBENn : in std_logic;
    CLK40B : out std_logic;
    TBI_CPUn : out std_logic;
    TAn : inout std_logic;
    CPUBGn : out std_logic;
    BUFENn : out std_logic;
    RnW : in std_logic;
    CLK80_CPU : out std_logic;
    BUFDIR : out std_logic;
    TCI_CPUn : out std_logic;
    TS_CPUn : in std_logic;
    CLKRAMB : out std_logic;
    CLK40A : out std_logic;
    TCIn : in std_logic;
    TBIn : in std_logic;
    DMAn : out std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    TACKn : inout std_logic;
    BGn : in std_logic);
end U111_TOP;

-- Architecture of U111_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U111_TOP is

signal \N__13681\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13647\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13618\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13600\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13582\ : std_logic;
signal \N__13575\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13566\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13548\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13528\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13519\ : std_logic;
signal \N__13512\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13501\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13483\ : std_logic;
signal \N__13476\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13458\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13429\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13395\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13377\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13366\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13357\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13321\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13285\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13242\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13240\ : std_logic;
signal \N__13233\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13206\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13204\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13006\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12721\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12714\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12678\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12605\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12382\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12335\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12211\ : std_logic;
signal \N__12208\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12136\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10434\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7972\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7275\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \TCIn_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \TAn_in\ : std_logic;
signal \N_237_i\ : std_logic;
signal \N_240_i\ : std_logic;
signal \N_242_i\ : std_logic;
signal \N_228_i\ : std_logic;
signal \N_241_i\ : std_logic;
signal \N_243_i\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_0\ : std_logic;
signal \N_229_i\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \N_231_i\ : std_logic;
signal \N_220_i\ : std_logic;
signal \N_230_i\ : std_logic;
signal \N_232_i\ : std_logic;
signal \N_222_i\ : std_logic;
signal \N_221_i\ : std_logic;
signal \N_233_i\ : std_logic;
signal \N_234_i\ : std_logic;
signal \N_235_i\ : std_logic;
signal \N_213_i\ : std_logic;
signal \N_223_i\ : std_logic;
signal \N_224_i\ : std_logic;
signal \N_217_i\ : std_logic;
signal \N_227_i\ : std_logic;
signal \N_226_i\ : std_logic;
signal \N_236_i\ : std_logic;
signal \N_239_i\ : std_logic;
signal \N_238_i\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep24_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep25_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep28_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep27_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep26_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep30_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep16_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep29_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep17_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep19_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep18_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep20_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep21_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep22_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep9_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep23_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep11_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep1_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep5_i_ess\ : std_logic;
signal \N_215_i\ : std_logic;
signal \U111_CYCLE_SM_A_AMIGA_0_i_1\ : std_logic;
signal \A_040_c_0\ : std_logic;
signal \A_AMIGA_c_0\ : std_logic;
signal \D_LL_AMIGA_in_7\ : std_logic;
signal \un2_D_LL_AMIGA_7\ : std_logic;
signal \D_LL_040_in_2\ : std_logic;
signal \D_UM_040_in_2\ : std_logic;
signal \un1_D_UM_040_2\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep8_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep10_i_ess\ : std_logic;
signal \D_LM_AMIGA_in_7\ : std_logic;
signal \un2_D_LM_AMIGA_7\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep12_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep14_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep6_i_ess\ : std_logic;
signal \N_218_i\ : std_logic;
signal \D_UU_040_in_7\ : std_logic;
signal \D_LM_040_in_7\ : std_logic;
signal \un1_D_UU_040_7\ : std_logic;
signal \N_219_i\ : std_logic;
signal \D_LL_AMIGA_in_5\ : std_logic;
signal \un2_D_LL_AMIGA_5\ : std_logic;
signal \D_LM_AMIGA_in_1\ : std_logic;
signal \un2_D_LM_AMIGA_1\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep15_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep3_i_ess\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep7_i_ess\ : std_logic;
signal \D_LM_AMIGA_in_3\ : std_logic;
signal \un2_D_LM_AMIGA_3\ : std_logic;
signal \D_LM_AMIGA_in_5\ : std_logic;
signal \un2_D_LM_AMIGA_5\ : std_logic;
signal \N_214_i\ : std_logic;
signal \D_UU_040_in_1\ : std_logic;
signal \D_LM_040_in_1\ : std_logic;
signal \un1_D_UU_040_1\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep0_i_ess\ : std_logic;
signal \N_212_i\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep4_i_ess\ : std_logic;
signal \N_216_i\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep2_i_ess\ : std_logic;
signal \N_225_i\ : std_logic;
signal \LBENn_c_i\ : std_logic;
signal \D_LL_AMIGA_in_0\ : std_logic;
signal \un2_D_LL_AMIGA_0\ : std_logic;
signal \D_LM_AMIGA_in_2\ : std_logic;
signal \un2_D_LM_AMIGA_2\ : std_logic;
signal \WRITE_CYCLE_ACTIVE_rep13_i_ess\ : std_logic;
signal \D_UU_040_in_5\ : std_logic;
signal \D_LM_040_in_5\ : std_logic;
signal \un1_D_UU_040_5\ : std_logic;
signal \D_LL_AMIGA_in_6\ : std_logic;
signal \un2_D_LL_AMIGA_6\ : std_logic;
signal \D_LM_AMIGA_in_0\ : std_logic;
signal \un2_D_LM_AMIGA_0\ : std_logic;
signal \D_LL_AMIGA_in_3\ : std_logic;
signal \un2_D_LL_AMIGA_3\ : std_logic;
signal \D_LL_AMIGA_in_4\ : std_logic;
signal \un2_D_LL_AMIGA_4\ : std_logic;
signal \D_LM_AMIGA_in_4\ : std_logic;
signal \un2_D_LM_AMIGA_4\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \LBENn_c_i_0\ : std_logic;
signal \D_LL_AMIGA_in_1\ : std_logic;
signal \un2_D_LL_AMIGA_1\ : std_logic;
signal \A_040_c_1\ : std_logic;
signal \TSn_c\ : std_logic;
signal \INVU111_CYCLE_SM.TSnC_net\ : std_logic;
signal \U111_CYCLE_SM.TS_ENZ0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_srsts_i_o2_0_5_cascade_\ : std_logic;
signal \U111_CYCLE_SM.N_148_cascade_\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_srsts_0_1_0_cascade_\ : std_logic;
signal \D_UU_AMIGA_in_1\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\ : std_logic;
signal \un1_D_UU_AMIGA_1\ : std_logic;
signal \D_LL_AMIGA_in_2\ : std_logic;
signal \un2_D_LL_AMIGA_2\ : std_logic;
signal \U111_CYCLE_SM.TS_ENZ0Z6\ : std_logic;
signal \U111_CYCLE_SM.N_158_cascade_\ : std_logic;
signal \U111_CYCLE_SM.N_130_0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\ : std_logic;
signal \U111_CYCLE_SM.TS_EN_6\ : std_logic;
signal \U111_CYCLE_SM.N_160_cascade_\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \U111_CYCLE_SM.PORT_MISMATCH_2_cascade_\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\ : std_logic;
signal \U111_CYCLE_SM.N_142_0\ : std_logic;
signal \TBIn_c\ : std_logic;
signal \U111_CYCLE_SM.un7_CYCLE_STATE_0_cascade_\ : std_logic;
signal \U111_CYCLE_SM.N_149\ : std_logic;
signal \U111_CYCLE_SM.BURSTZ0\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\ : std_logic;
signal \U111_CYCLE_SM.BURST_COUNTZ0Z_0\ : std_logic;
signal \U111_CYCLE_SM.N_132_0_cascade_\ : std_logic;
signal \U111_CYCLE_SM.BURST_COUNTZ0Z_1\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_RNIGD6KZ0Z_2_cascade_\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1_cascade_\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_RNIGD6KZ0Z_2\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \TEAn_c\ : std_logic;
signal \U111_CYCLE_SM.un7_CYCLE_STATE_0\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_srsts_i_1_2_cascade_\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\ : std_logic;
signal \D_UM_AMIGA_in_1\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\ : std_logic;
signal \un1_D_UM_AMIGA_1\ : std_logic;
signal \CLK80\ : std_logic;
signal \GB_BUFFER_CLK80_THRU_CO\ : std_logic;
signal \D_LM_AMIGA_in_6\ : std_logic;
signal \un2_D_LM_AMIGA_6\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\ : std_logic;
signal \D_UM_AMIGA_in_5\ : std_logic;
signal \un1_D_UM_AMIGA_5\ : std_logic;
signal \D_UM_AMIGA_in_7\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\ : std_logic;
signal \un1_D_UM_AMIGA_7\ : std_logic;
signal \D_UU_AMIGA_in_0\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\ : std_logic;
signal \un1_D_UU_AMIGA_0\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\ : std_logic;
signal \D_UU_AMIGA_in_7\ : std_logic;
signal \un1_D_UU_AMIGA_7\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\ : std_logic;
signal \D_UU_AMIGA_in_2\ : std_logic;
signal \un1_D_UU_AMIGA_2\ : std_logic;
signal \U111_CYCLE_SM.FLIP_WORD_2\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\ : std_logic;
signal \U111_CYCLE_SM.N_160\ : std_logic;
signal \U111_CYCLE_SM.A2_ENZ0\ : std_logic;
signal \U111_CYCLE_SM.un1_CYCLE_STATE_1_0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\ : std_logic;
signal \un1_D_UM_AMIGA_0\ : std_logic;
signal \U111_CYCLE_SM.LW_TRANSZ0\ : std_logic;
signal \PORTSIZE_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\ : std_logic;
signal \U111_CYCLE_SM.PORT_MISMATCHZ0\ : std_logic;
signal \un1_D_UM_AMIGA_2\ : std_logic;
signal \D_UM_AMIGA_in_6\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\ : std_logic;
signal \un1_D_UM_AMIGA_6\ : std_logic;
signal \D_UM_AMIGA_in_2\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\ : std_logic;
signal \D_UM_AMIGA_in_0\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\ : std_logic;
signal \U111_CYCLE_SM.N_159_0\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1\ : std_logic;
signal \U111_CYCLE_SM.TA_DISZ0\ : std_logic;
signal \TAn_1_i\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\ : std_logic;
signal \D_UU_AMIGA_in_3\ : std_logic;
signal \un1_D_UU_AMIGA_3\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\ : std_logic;
signal \D_UM_AMIGA_in_3\ : std_logic;
signal \un1_D_UM_AMIGA_3\ : std_logic;
signal \D_UM_AMIGA_in_4\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\ : std_logic;
signal \un1_D_UM_AMIGA_4\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\ : std_logic;
signal \D_UU_AMIGA_in_5\ : std_logic;
signal \un1_D_UU_AMIGA_5\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\ : std_logic;
signal \D_UU_AMIGA_in_4\ : std_logic;
signal \un1_D_UU_AMIGA_4\ : std_logic;
signal \D_UU_AMIGA_in_6\ : std_logic;
signal \U111_CYCLE_SM.LATCH_ENZ0\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\ : std_logic;
signal \un1_D_UU_AMIGA_6\ : std_logic;
signal \D_LM_040_in_6\ : std_logic;
signal \D_UU_040_in_6\ : std_logic;
signal \un1_D_UU_040_6\ : std_logic;
signal \D_UM_040_in_6\ : std_logic;
signal \D_LL_040_in_6\ : std_logic;
signal \un1_D_UM_040_6\ : std_logic;
signal \D_LL_040_in_4\ : std_logic;
signal \D_UM_040_in_4\ : std_logic;
signal \un1_D_UM_040_4\ : std_logic;
signal \D_UM_040_in_5\ : std_logic;
signal \D_LL_040_in_5\ : std_logic;
signal \un1_D_UM_040_5\ : std_logic;
signal \D_LL_040_in_1\ : std_logic;
signal \D_UM_040_in_1\ : std_logic;
signal \un1_D_UM_040_1\ : std_logic;
signal \D_LM_040_in_2\ : std_logic;
signal \D_UU_040_in_2\ : std_logic;
signal \un1_D_UU_040_2\ : std_logic;
signal \D_UU_040_in_0\ : std_logic;
signal \D_LM_040_in_0\ : std_logic;
signal \un1_D_UU_040_0\ : std_logic;
signal \D_LM_040_in_3\ : std_logic;
signal \D_UU_040_in_3\ : std_logic;
signal \un1_D_UU_040_3\ : std_logic;
signal \D_UU_040_in_4\ : std_logic;
signal \D_LM_040_in_4\ : std_logic;
signal \un1_D_UU_040_4\ : std_logic;
signal \D_UM_040_in_0\ : std_logic;
signal \D_LL_040_in_0\ : std_logic;
signal \un1_D_UM_040_0\ : std_logic;
signal \D_UM_040_in_3\ : std_logic;
signal \D_LL_040_in_3\ : std_logic;
signal \un1_D_UM_040_3\ : std_logic;
signal \U111_CYCLE_SM.FLIP_WORDZ0\ : std_logic;
signal \D_LL_040_in_7\ : std_logic;
signal \D_UM_040_in_7\ : std_logic;
signal \un1_D_UM_040_7\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep4_i_ess\ : std_logic;
signal \N_184_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep2_i_ess\ : std_logic;
signal \N_182_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep0_i_ess\ : std_logic;
signal \N_180_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep7_i_ess\ : std_logic;
signal \N_187_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep6_i_ess\ : std_logic;
signal \N_186_i\ : std_logic;
signal \N_207_i\ : std_logic;
signal \N_205_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep27_i_ess\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep25_i_ess\ : std_logic;
signal \N_196_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep16_i_ess\ : std_logic;
signal \GB_BUFFER_CLK40_THRU_CO\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep5_i_ess\ : std_logic;
signal \N_185_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep13_i_ess\ : std_logic;
signal \N_193_i\ : std_logic;
signal \N_208_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep28_i_ess\ : std_logic;
signal \N_204_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep30_i_ess\ : std_logic;
signal \N_210_i\ : std_logic;
signal \N_206_i\ : std_logic;
signal \N_209_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep29_i_ess\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep24_i_ess\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep26_i_ess\ : std_logic;
signal \N_197_i\ : std_logic;
signal \N_211_i\ : std_logic;
signal \N_198_i\ : std_logic;
signal \N_199_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep31_i_ess\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep19_i_ess\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep18_i_ess\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep17_i_ess\ : std_logic;
signal \N_200_i\ : std_logic;
signal \N_188_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep21_i_ess\ : std_logic;
signal \N_201_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep20_i_ess\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep8_i_ess\ : std_logic;
signal \N_190_i\ : std_logic;
signal \N_194_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep14_i_ess\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep10_i_ess\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep22_i_ess\ : std_logic;
signal \N_202_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep23_i_ess\ : std_logic;
signal \N_203_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep9_i_ess\ : std_logic;
signal \N_189_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep11_i_ess\ : std_logic;
signal \N_191_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep15_i_ess\ : std_logic;
signal \N_195_i\ : std_logic;
signal \RnW_c\ : std_logic;
signal \TS_CPUn_c\ : std_logic;
signal \LBENn_c\ : std_logic;
signal \BGn_c\ : std_logic;
signal \CLK40\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_g_0\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep1_i_ess\ : std_logic;
signal \N_181_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep12_i_ess\ : std_logic;
signal \N_192_i\ : std_logic;
signal \READ_CYCLE_ACTIVE_rep3_i_ess\ : std_logic;
signal \N_183_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK40_IN_wire\ : std_logic;
signal \LBENn_wire\ : std_logic;
signal \CPUBGn_wire\ : std_logic;
signal \A_040_wire\ : std_logic_vector(1 downto 0);
signal \CLK40B_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \BUFDIR_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \TS_CPUn_wire\ : std_logic;
signal \CLKRAMB_wire\ : std_logic;
signal \TEAn_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \DMAn_wire\ : std_logic;
signal \CLK80_CPU_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \A_AMIGA_wire\ : std_logic_vector(1 downto 0);
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \BGn_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \TBI_CPUn_wire\ : std_logic;
signal \CLK40A_wire\ : std_logic;
signal \CLKRAMA_wire\ : std_logic;
signal \TCI_CPUn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \TEA_CPUn_wire\ : std_logic;
signal \pll_pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK40_IN_wire\ <= CLK40_IN;
    \LBENn_wire\ <= LBENn;
    CPUBGn <= \CPUBGn_wire\;
    \A_040_wire\ <= A_040;
    CLK40B <= \CLK40B_wire\;
    \TBIn_wire\ <= TBIn;
    BUFDIR <= \BUFDIR_wire\;
    \SIZ_wire\ <= SIZ;
    \TS_CPUn_wire\ <= TS_CPUn;
    CLKRAMB <= \CLKRAMB_wire\;
    \TEAn_wire\ <= TEAn;
    BUFENn <= \BUFENn_wire\;
    DMAn <= \DMAn_wire\;
    CLK80_CPU <= \CLK80_CPU_wire\;
    TSn <= \TSn_wire\;
    \PORTSIZE_wire\ <= PORTSIZE;
    A_AMIGA <= \A_AMIGA_wire\;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    \BGn_wire\ <= BGn;
    \TCIn_wire\ <= TCIn;
    TBI_CPUn <= \TBI_CPUn_wire\;
    CLK40A <= \CLK40A_wire\;
    CLKRAMA <= \CLKRAMA_wire\;
    TCI_CPUn <= \TCI_CPUn_wire\;
    \RnW_wire\ <= RnW;
    TEA_CPUn <= \TEA_CPUn_wire\;
    \pll_pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll_pll\ : PLL40_2F
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            SCLK => '0',
            PLLOUTGLOBALA => \CLK80\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALB => \CLK40\,
            SDI => '0',
            PLLOUTCOREA => OPEN,
            BYPASS => '0',
            RESETB => \N__5485\,
            PLLOUTCOREB => OPEN,
            LOCK => OPEN,
            SDO => OPEN,
            EXTFEEDBACK => '0',
            DYNAMICDELAY => \pll_pll_DYNAMICDELAY_wire\,
            PLLIN => \N__13681\
        );

    \pll_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \VCCG0\,
            DIN => '0',
            DOUT => \N__13681\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \LBENn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13665\,
            DIN => \N__13664\,
            DOUT => \N__13663\,
            PACKAGEPIN => \LBENn_wire\
        );

    \LBENn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13665\,
            PADOUT => \N__13664\,
            PADIN => \N__13663\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \LBENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TAn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13656\,
            DIN => \N__13655\,
            DOUT => \N__13654\,
            PACKAGEPIN => TAn
        );

    \TAn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13656\,
            PADOUT => \N__13655\,
            PADIN => \N__13654\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7811\,
            DIN0 => \TAn_in\,
            DOUT0 => \N__6287\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13647\,
            DIN => \N__13646\,
            DOUT => \N__13645\,
            PACKAGEPIN => D_LL_AMIGA(1)
        );

    \D_LL_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13647\,
            PADOUT => \N__13646\,
            PADIN => \N__13645\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4184\,
            DIN0 => \D_LL_AMIGA_in_1\,
            DOUT0 => \N__7988\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13638\,
            DIN => \N__13637\,
            DOUT => \N__13636\,
            PACKAGEPIN => D_UU_040(6)
        );

    \D_UU_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13638\,
            PADOUT => \N__13637\,
            PADIN => \N__13636\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9527\,
            DIN0 => \D_UU_040_in_6\,
            DOUT0 => \N__8333\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CPUBGn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__13629\,
            DIN => \N__13628\,
            DOUT => \N__13627\,
            PACKAGEPIN => \CPUBGn_wire\
        );

    \CPUBGn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13629\,
            PADOUT => \N__13628\,
            PADIN => \N__13627\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13620\,
            DIN => \N__13619\,
            DOUT => \N__13618\,
            PACKAGEPIN => D_UM_AMIGA(3)
        );

    \D_UM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13620\,
            PADOUT => \N__13619\,
            PADIN => \N__13618\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4448\,
            DIN0 => \D_UM_AMIGA_in_3\,
            DOUT0 => \N__9044\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__13611\,
            DIN => \N__13610\,
            DOUT => \N__13609\,
            PACKAGEPIN => \A_040_wire\(1)
        );

    \A_040_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13611\,
            PADOUT => \N__13610\,
            PADIN => \N__13609\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13602\,
            DIN => \N__13601\,
            DOUT => \N__13600\,
            PACKAGEPIN => D_LM_AMIGA(4)
        );

    \D_LM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13602\,
            PADOUT => \N__13601\,
            PADIN => \N__13600\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4280\,
            DIN0 => \D_LM_AMIGA_in_4\,
            DOUT0 => \N__9245\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13593\,
            DIN => \N__13592\,
            DOUT => \N__13591\,
            PACKAGEPIN => D_LM_040(7)
        );

    \D_LM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13593\,
            PADOUT => \N__13592\,
            PADIN => \N__13591\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10082\,
            DIN0 => \D_LM_040_in_7\,
            DOUT0 => \N__5000\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13584\,
            DIN => \N__13583\,
            DOUT => \N__13582\,
            PACKAGEPIN => \CLK40B_wire\
        );

    \CLK40B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13584\,
            PADOUT => \N__13583\,
            PADIN => \N__13582\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9674\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13575\,
            DIN => \N__13574\,
            DOUT => \N__13573\,
            PACKAGEPIN => D_UM_040(1)
        );

    \D_UM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13575\,
            PADOUT => \N__13574\,
            PADIN => \N__13573\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__12776\,
            DIN0 => \D_UM_040_in_1\,
            DOUT0 => \N__6569\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13566\,
            DIN => \N__13565\,
            DOUT => \N__13564\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13566\,
            PADOUT => \N__13565\,
            PADIN => \N__13564\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TBIn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13557\,
            DIN => \N__13556\,
            DOUT => \N__13555\,
            PACKAGEPIN => D_UU_AMIGA(7)
        );

    \D_UU_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13557\,
            PADOUT => \N__13556\,
            PADIN => \N__13555\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4865\,
            DIN0 => \D_UU_AMIGA_in_7\,
            DOUT0 => \N__4883\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13548\,
            DIN => \N__13547\,
            DOUT => \N__13546\,
            PACKAGEPIN => \BUFDIR_wire\
        );

    \BUFDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13548\,
            PADOUT => \N__13547\,
            PADIN => \N__13546\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12718\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13539\,
            DIN => \N__13538\,
            DOUT => \N__13537\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13539\,
            PADOUT => \N__13538\,
            PADIN => \N__13537\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TS_CPUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13530\,
            DIN => \N__13529\,
            DOUT => \N__13528\,
            PACKAGEPIN => \TS_CPUn_wire\
        );

    \TS_CPUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13530\,
            PADOUT => \N__13529\,
            PADIN => \N__13528\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TS_CPUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13521\,
            DIN => \N__13520\,
            DOUT => \N__13519\,
            PACKAGEPIN => D_LL_040(1)
        );

    \D_LL_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13521\,
            PADOUT => \N__13520\,
            PADIN => \N__13519\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9731\,
            DIN0 => \D_LL_040_in_1\,
            DOUT0 => \N__5423\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13512\,
            DIN => \N__13511\,
            DOUT => \N__13510\,
            PACKAGEPIN => D_UU_040(1)
        );

    \D_UU_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13512\,
            PADOUT => \N__13511\,
            PADIN => \N__13510\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10157\,
            DIN0 => \D_UU_040_in_1\,
            DOUT0 => \N__5933\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13503\,
            DIN => \N__13502\,
            DOUT => \N__13501\,
            PACKAGEPIN => D_LM_AMIGA(1)
        );

    \D_LM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13503\,
            PADOUT => \N__13502\,
            PADIN => \N__13501\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4085\,
            DIN0 => \D_LM_AMIGA_in_1\,
            DOUT0 => \N__5062\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13494\,
            DIN => \N__13493\,
            DOUT => \N__13492\,
            PACKAGEPIN => D_LM_040(2)
        );

    \D_LM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13494\,
            PADOUT => \N__13493\,
            PADIN => \N__13492\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9929\,
            DIN0 => \D_LM_040_in_2\,
            DOUT0 => \N__5249\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__13485\,
            DIN => \N__13484\,
            DOUT => \N__13483\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13485\,
            PADOUT => \N__13484\,
            PADIN => \N__13483\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5450\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__4208\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13476\,
            DIN => \N__13475\,
            DOUT => \N__13474\,
            PACKAGEPIN => D_UM_040(2)
        );

    \D_UM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13476\,
            PADOUT => \N__13475\,
            PADIN => \N__13474\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10004\,
            DIN0 => \D_UM_040_in_2\,
            DOUT0 => \N__7418\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMB_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13467\,
            DIN => \N__13466\,
            DOUT => \N__13465\,
            PACKAGEPIN => \CLKRAMB_wire\
        );

    \CLKRAMB_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13467\,
            PADOUT => \N__13466\,
            PADIN => \N__13465\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6536\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13458\,
            DIN => \N__13457\,
            DOUT => \N__13456\,
            PACKAGEPIN => D_LL_AMIGA(2)
        );

    \D_LL_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13458\,
            PADOUT => \N__13457\,
            PADIN => \N__13456\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4334\,
            DIN0 => \D_LL_AMIGA_in_2\,
            DOUT0 => \N__4693\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13449\,
            DIN => \N__13448\,
            DOUT => \N__13447\,
            PACKAGEPIN => D_UU_AMIGA(2)
        );

    \D_UU_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13449\,
            PADOUT => \N__13448\,
            PADIN => \N__13447\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5102\,
            DIN0 => \D_UU_AMIGA_in_2\,
            DOUT0 => \N__9458\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TEAn_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__13440\,
            DIN => \N__13439\,
            DOUT => \N__13438\,
            PACKAGEPIN => \TEAn_wire\
        );

    \TEAn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13440\,
            PADOUT => \N__13439\,
            PADIN => \N__13438\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TEAn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13431\,
            DIN => \N__13430\,
            DOUT => \N__13429\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13431\,
            PADOUT => \N__13430\,
            PADIN => \N__13429\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5318\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMAn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13422\,
            DIN => \N__13421\,
            DOUT => \N__13420\,
            PACKAGEPIN => \DMAn_wire\
        );

    \DMAn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13422\,
            PADOUT => \N__13421\,
            PADIN => \N__13420\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5486\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13413\,
            DIN => \N__13412\,
            DOUT => \N__13411\,
            PACKAGEPIN => D_LL_040(6)
        );

    \D_LL_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13413\,
            PADOUT => \N__13412\,
            PADIN => \N__13411\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9797\,
            DIN0 => \D_LL_040_in_6\,
            DOUT0 => \N__5666\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13404\,
            DIN => \N__13403\,
            DOUT => \N__13402\,
            PACKAGEPIN => D_LL_AMIGA(5)
        );

    \D_LL_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13404\,
            PADOUT => \N__13403\,
            PADIN => \N__13402\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4127\,
            DIN0 => \D_LL_AMIGA_in_5\,
            DOUT0 => \N__8057\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13395\,
            DIN => \N__13394\,
            DOUT => \N__13393\,
            PACKAGEPIN => D_UM_AMIGA(0)
        );

    \D_UM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13395\,
            PADOUT => \N__13394\,
            PADIN => \N__13393\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4298\,
            DIN0 => \D_UM_AMIGA_in_0\,
            DOUT0 => \N__9134\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13386\,
            DIN => \N__13385\,
            DOUT => \N__13384\,
            PACKAGEPIN => D_UU_040(2)
        );

    \D_UU_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13386\,
            PADOUT => \N__13385\,
            PADIN => \N__13384\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9593\,
            DIN0 => \D_UU_040_in_2\,
            DOUT0 => \N__6884\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13377\,
            DIN => \N__13376\,
            DOUT => \N__13375\,
            PACKAGEPIN => D_LM_AMIGA(2)
        );

    \D_LM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13377\,
            PADOUT => \N__13376\,
            PADIN => \N__13375\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4289\,
            DIN0 => \D_LM_AMIGA_in_2\,
            DOUT0 => \N__9511\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK80_CPU_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13368\,
            DIN => \N__13367\,
            DOUT => \N__13366\,
            PACKAGEPIN => \CLK80_CPU_wire\
        );

    \CLK80_CPU_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13368\,
            PADOUT => \N__13367\,
            PADIN => \N__13366\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6529\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13359\,
            DIN => \N__13358\,
            DOUT => \N__13357\,
            PACKAGEPIN => D_LL_040(3)
        );

    \D_LL_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13359\,
            PADOUT => \N__13358\,
            PADIN => \N__13357\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9749\,
            DIN0 => \D_LL_040_in_3\,
            DOUT0 => \N__5585\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13350\,
            DIN => \N__13349\,
            DOUT => \N__13348\,
            PACKAGEPIN => D_LM_040(1)
        );

    \D_LM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13350\,
            PADOUT => \N__13349\,
            PADIN => \N__13348\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9962\,
            DIN0 => \D_LM_040_in_1\,
            DOUT0 => \N__5228\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13341\,
            DIN => \N__13340\,
            DOUT => \N__13339\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13341\,
            PADOUT => \N__13340\,
            PADIN => \N__13339\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5801\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13332\,
            DIN => \N__13331\,
            DOUT => \N__13330\,
            PACKAGEPIN => D_UM_AMIGA(7)
        );

    \D_UM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13332\,
            PADOUT => \N__13331\,
            PADIN => \N__13330\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4400\,
            DIN0 => \D_UM_AMIGA_in_7\,
            DOUT0 => \N__8657\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13323\,
            DIN => \N__13322\,
            DOUT => \N__13321\,
            PACKAGEPIN => D_LM_AMIGA(7)
        );

    \D_LM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13323\,
            PADOUT => \N__13322\,
            PADIN => \N__13321\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4478\,
            DIN0 => \D_LM_AMIGA_in_7\,
            DOUT0 => \N__4919\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13314\,
            DIN => \N__13313\,
            DOUT => \N__13312\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13314\,
            PADOUT => \N__13313\,
            PADIN => \N__13312\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \PORTSIZE_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__13305\,
            DIN => \N__13304\,
            DOUT => \N__13303\,
            PACKAGEPIN => \A_AMIGA_wire\(0)
        );

    \A_AMIGA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13305\,
            PADOUT => \N__13304\,
            PADIN => \N__13303\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4751\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13296\,
            DIN => \N__13295\,
            DOUT => \N__13294\,
            PACKAGEPIN => D_LM_040(4)
        );

    \D_LM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13296\,
            PADOUT => \N__13295\,
            PADIN => \N__13294\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10055\,
            DIN0 => \D_LM_040_in_4\,
            DOUT0 => \N__5510\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13287\,
            DIN => \N__13286\,
            DOUT => \N__13285\,
            PACKAGEPIN => D_UM_040(7)
        );

    \D_UM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13287\,
            PADOUT => \N__13286\,
            PADIN => \N__13285\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__12734\,
            DIN0 => \D_UM_040_in_7\,
            DOUT0 => \N__7097\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13278\,
            DIN => \N__13277\,
            DOUT => \N__13276\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13278\,
            PADOUT => \N__13277\,
            PADIN => \N__13276\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13269\,
            DIN => \N__13268\,
            DOUT => \N__13267\,
            PACKAGEPIN => D_UU_AMIGA(1)
        );

    \D_UU_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13269\,
            PADOUT => \N__13268\,
            PADIN => \N__13267\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4463\,
            DIN0 => \D_UU_AMIGA_in_1\,
            DOUT0 => \N__5399\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13260\,
            DIN => \N__13259\,
            DOUT => \N__13258\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13260\,
            PADOUT => \N__13259\,
            PADIN => \N__13258\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9666\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13251\,
            DIN => \N__13250\,
            DOUT => \N__13249\,
            PACKAGEPIN => D_UM_040(0)
        );

    \D_UM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13251\,
            PADOUT => \N__13250\,
            PADIN => \N__13249\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10040\,
            DIN0 => \D_UM_040_in_0\,
            DOUT0 => \N__7559\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13242\,
            DIN => \N__13241\,
            DOUT => \N__13240\,
            PACKAGEPIN => D_LL_AMIGA(0)
        );

    \D_LL_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13242\,
            PADOUT => \N__13241\,
            PADIN => \N__13240\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4367\,
            DIN0 => \D_LL_AMIGA_in_0\,
            DOUT0 => \N__9173\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13233\,
            DIN => \N__13232\,
            DOUT => \N__13231\,
            PACKAGEPIN => D_UU_AMIGA(4)
        );

    \D_UU_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13233\,
            PADOUT => \N__13232\,
            PADIN => \N__13231\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5351\,
            DIN0 => \D_UU_AMIGA_in_4\,
            DOUT0 => \N__9206\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13224\,
            DIN => \N__13223\,
            DOUT => \N__13222\,
            PACKAGEPIN => D_UU_040(7)
        );

    \D_UU_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13224\,
            PADOUT => \N__13223\,
            PADIN => \N__13222\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9545\,
            DIN0 => \D_UU_040_in_7\,
            DOUT0 => \N__6953\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13215\,
            DIN => \N__13214\,
            DOUT => \N__13213\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13215\,
            PADOUT => \N__13214\,
            PADIN => \N__13213\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BGn_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__13206\,
            DIN => \N__13205\,
            DOUT => \N__13204\,
            PACKAGEPIN => \BGn_wire\
        );

    \BGn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13206\,
            PADOUT => \N__13205\,
            PADIN => \N__13204\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \BGn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13197\,
            DIN => \N__13196\,
            DOUT => \N__13195\,
            PACKAGEPIN => D_LL_040(0)
        );

    \D_LL_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13197\,
            PADOUT => \N__13196\,
            PADIN => \N__13195\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9821\,
            DIN0 => \D_LL_040_in_0\,
            DOUT0 => \N__5282\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13188\,
            DIN => \N__13187\,
            DOUT => \N__13186\,
            PACKAGEPIN => D_UM_AMIGA(2)
        );

    \D_UM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13188\,
            PADOUT => \N__13187\,
            PADIN => \N__13186\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4268\,
            DIN0 => \D_UM_AMIGA_in_2\,
            DOUT0 => \N__4631\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13179\,
            DIN => \N__13178\,
            DOUT => \N__13177\,
            PACKAGEPIN => D_UU_040(0)
        );

    \D_UU_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13179\,
            PADOUT => \N__13178\,
            PADIN => \N__13177\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9572\,
            DIN0 => \D_UU_040_in_0\,
            DOUT0 => \N__7022\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13170\,
            DIN => \N__13169\,
            DOUT => \N__13168\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13170\,
            PADOUT => \N__13169\,
            PADIN => \N__13168\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TCIn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__13161\,
            DIN => \N__13160\,
            DOUT => \N__13159\,
            PACKAGEPIN => \A_040_wire\(0)
        );

    \A_040_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13161\,
            PADOUT => \N__13160\,
            PADIN => \N__13159\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13152\,
            DIN => \N__13151\,
            DOUT => \N__13150\,
            PACKAGEPIN => D_LM_AMIGA(0)
        );

    \D_LM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13152\,
            PADOUT => \N__13151\,
            PADIN => \N__13150\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4142\,
            DIN0 => \D_LM_AMIGA_in_0\,
            DOUT0 => \N__9416\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13143\,
            DIN => \N__13142\,
            DOUT => \N__13141\,
            PACKAGEPIN => \TBI_CPUn_wire\
        );

    \TBI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13143\,
            PADOUT => \N__13142\,
            PADIN => \N__13141\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6010\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13134\,
            DIN => \N__13133\,
            DOUT => \N__13132\,
            PACKAGEPIN => \CLK40A_wire\
        );

    \CLK40A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13134\,
            PADOUT => \N__13133\,
            PADIN => \N__13132\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9642\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13125\,
            DIN => \N__13124\,
            DOUT => \N__13123\,
            PACKAGEPIN => D_LM_040(3)
        );

    \D_LM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13125\,
            PADOUT => \N__13124\,
            PADIN => \N__13123\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9914\,
            DIN0 => \D_LM_040_in_3\,
            DOUT0 => \N__5165\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13116\,
            DIN => \N__13115\,
            DOUT => \N__13114\,
            PACKAGEPIN => D_LM_AMIGA(5)
        );

    \D_LM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13116\,
            PADOUT => \N__13115\,
            PADIN => \N__13114\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4238\,
            DIN0 => \D_LM_AMIGA_in_5\,
            DOUT0 => \N__5744\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13107\,
            DIN => \N__13106\,
            DOUT => \N__13105\,
            PACKAGEPIN => D_LM_040(6)
        );

    \D_LM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13107\,
            PADOUT => \N__13106\,
            PADIN => \N__13105\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10103\,
            DIN0 => \D_LM_040_in_6\,
            DOUT0 => \N__6473\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13098\,
            DIN => \N__13097\,
            DOUT => \N__13096\,
            PACKAGEPIN => D_UM_040(5)
        );

    \D_UM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13098\,
            PADOUT => \N__13097\,
            PADIN => \N__13096\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9857\,
            DIN0 => \D_UM_040_in_5\,
            DOUT0 => \N__7169\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13089\,
            DIN => \N__13088\,
            DOUT => \N__13087\,
            PACKAGEPIN => D_LL_AMIGA(3)
        );

    \D_LL_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13089\,
            PADOUT => \N__13088\,
            PADIN => \N__13087\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4352\,
            DIN0 => \D_LL_AMIGA_in_3\,
            DOUT0 => \N__9092\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13080\,
            DIN => \N__13079\,
            DOUT => \N__13078\,
            PACKAGEPIN => D_UU_AMIGA(3)
        );

    \D_UU_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13080\,
            PADOUT => \N__13079\,
            PADIN => \N__13078\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4790\,
            DIN0 => \D_UU_AMIGA_in_3\,
            DOUT0 => \N__9284\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13071\,
            DIN => \N__13070\,
            DOUT => \N__13069\,
            PACKAGEPIN => D_LL_040(5)
        );

    \D_LL_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13071\,
            PADOUT => \N__13070\,
            PADIN => \N__13069\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9764\,
            DIN0 => \D_LL_040_in_5\,
            DOUT0 => \N__4835\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13062\,
            DIN => \N__13061\,
            DOUT => \N__13060\,
            PACKAGEPIN => D_LL_AMIGA(6)
        );

    \D_LL_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13062\,
            PADOUT => \N__13061\,
            PADIN => \N__13060\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4157\,
            DIN0 => \D_LL_AMIGA_in_6\,
            DOUT0 => \N__8222\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13053\,
            DIN => \N__13052\,
            DOUT => \N__13051\,
            PACKAGEPIN => D_UU_AMIGA(6)
        );

    \D_UU_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13053\,
            PADOUT => \N__13052\,
            PADIN => \N__13051\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4958\,
            DIN0 => \D_UU_AMIGA_in_6\,
            DOUT0 => \N__8261\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13044\,
            DIN => \N__13043\,
            DOUT => \N__13042\,
            PACKAGEPIN => D_UM_AMIGA(1)
        );

    \D_UM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13044\,
            PADOUT => \N__13043\,
            PADIN => \N__13042\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4253\,
            DIN0 => \D_UM_AMIGA_in_1\,
            DOUT0 => \N__7928\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13035\,
            DIN => \N__13034\,
            DOUT => \N__13033\,
            PACKAGEPIN => D_UU_040(5)
        );

    \D_UU_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13035\,
            PADOUT => \N__13034\,
            PADIN => \N__13033\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9878\,
            DIN0 => \D_UU_040_in_5\,
            DOUT0 => \N__8579\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13026\,
            DIN => \N__13025\,
            DOUT => \N__13024\,
            PACKAGEPIN => \CLKRAMA_wire\
        );

    \CLKRAMA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13026\,
            PADOUT => \N__13025\,
            PADIN => \N__13024\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9667\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13017\,
            DIN => \N__13016\,
            DOUT => \N__13015\,
            PACKAGEPIN => D_LL_040(2)
        );

    \D_LL_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13017\,
            PADOUT => \N__13016\,
            PADIN => \N__13015\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9779\,
            DIN0 => \D_LL_040_in_2\,
            DOUT0 => \N__5894\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13008\,
            DIN => \N__13007\,
            DOUT => \N__13006\,
            PACKAGEPIN => \TCI_CPUn_wire\
        );

    \TCI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13008\,
            PADOUT => \N__13007\,
            PADIN => \N__13006\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4076\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12999\,
            DIN => \N__12998\,
            DOUT => \N__12997\,
            PACKAGEPIN => D_UM_AMIGA(4)
        );

    \D_UM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12999\,
            PADOUT => \N__12998\,
            PADIN => \N__12997\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4433\,
            DIN0 => \D_UM_AMIGA_in_4\,
            DOUT0 => \N__8096\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12990\,
            DIN => \N__12989\,
            DOUT => \N__12988\,
            PACKAGEPIN => D_LM_AMIGA(6)
        );

    \D_LM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12990\,
            PADOUT => \N__12989\,
            PADIN => \N__12988\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4223\,
            DIN0 => \D_LM_AMIGA_in_6\,
            DOUT0 => \N__8318\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12981\,
            DIN => \N__12980\,
            DOUT => \N__12979\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12981\,
            PADOUT => \N__12980\,
            PADIN => \N__12979\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12972\,
            DIN => \N__12971\,
            DOUT => \N__12970\,
            PACKAGEPIN => D_LM_040(5)
        );

    \D_LM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12972\,
            PADOUT => \N__12971\,
            PADIN => \N__12970\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10025\,
            DIN0 => \D_LM_040_in_5\,
            DOUT0 => \N__5126\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12963\,
            DIN => \N__12962\,
            DOUT => \N__12961\,
            PACKAGEPIN => D_UM_040(6)
        );

    \D_UM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12963\,
            PADOUT => \N__12962\,
            PADIN => \N__12961\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9992\,
            DIN0 => \D_UM_040_in_6\,
            DOUT0 => \N__7352\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12954\,
            DIN => \N__12953\,
            DOUT => \N__12952\,
            PACKAGEPIN => D_UM_040(3)
        );

    \D_UM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12954\,
            PADOUT => \N__12953\,
            PADIN => \N__12952\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__12755\,
            DIN0 => \D_UM_040_in_3\,
            DOUT0 => \N__7658\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12945\,
            DIN => \N__12944\,
            DOUT => \N__12943\,
            PACKAGEPIN => D_UU_AMIGA(5)
        );

    \D_UU_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12945\,
            PADOUT => \N__12944\,
            PADIN => \N__12943\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4418\,
            DIN0 => \D_UU_AMIGA_in_5\,
            DOUT0 => \N__5699\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12936\,
            DIN => \N__12935\,
            DOUT => \N__12934\,
            PACKAGEPIN => D_LL_040(7)
        );

    \D_LL_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12936\,
            PADOUT => \N__12935\,
            PADIN => \N__12934\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9947\,
            DIN0 => \D_LL_040_in_7\,
            DOUT0 => \N__4718\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12927\,
            DIN => \N__12926\,
            DOUT => \N__12925\,
            PACKAGEPIN => D_LL_AMIGA(4)
        );

    \D_LL_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12927\,
            PADOUT => \N__12926\,
            PADIN => \N__12925\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4172\,
            DIN0 => \D_LL_AMIGA_in_4\,
            DOUT0 => \N__8155\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12918\,
            DIN => \N__12917\,
            DOUT => \N__12916\,
            PACKAGEPIN => D_UU_040(3)
        );

    \D_UU_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12918\,
            PADOUT => \N__12917\,
            PADIN => \N__12916\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__12794\,
            DIN0 => \D_UU_040_in_3\,
            DOUT0 => \N__7733\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TEA_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12909\,
            DIN => \N__12908\,
            DOUT => \N__12907\,
            PACKAGEPIN => \TEA_CPUn_wire\
        );

    \TEA_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12909\,
            PADOUT => \N__12908\,
            PADIN => \N__12907\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6205\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12900\,
            DIN => \N__12899\,
            DOUT => \N__12898\,
            PACKAGEPIN => D_LM_AMIGA(3)
        );

    \D_LM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12900\,
            PADOUT => \N__12899\,
            PADIN => \N__12898\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4307\,
            DIN0 => \D_LM_AMIGA_in_3\,
            DOUT0 => \N__9347\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12891\,
            DIN => \N__12890\,
            DOUT => \N__12889\,
            PACKAGEPIN => D_LM_040(0)
        );

    \D_LM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12891\,
            PADOUT => \N__12890\,
            PADIN => \N__12889\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9698\,
            DIN0 => \D_LM_040_in_0\,
            DOUT0 => \N__5624\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12882\,
            DIN => \N__12881\,
            DOUT => \N__12880\,
            PACKAGEPIN => D_UM_AMIGA(6)
        );

    \D_UM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12882\,
            PADOUT => \N__12881\,
            PADIN => \N__12880\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4385\,
            DIN0 => \D_UM_AMIGA_in_6\,
            DOUT0 => \N__8174\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__12873\,
            DIN => \N__12872\,
            DOUT => \N__12871\,
            PACKAGEPIN => \A_AMIGA_wire\(1)
        );

    \A_AMIGA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12873\,
            PADOUT => \N__12872\,
            PADIN => \N__12871\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4775\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12864\,
            DIN => \N__12863\,
            DOUT => \N__12862\,
            PACKAGEPIN => D_UM_040(4)
        );

    \D_UM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12864\,
            PADOUT => \N__12863\,
            PADIN => \N__12862\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10136\,
            DIN0 => \D_UM_040_in_4\,
            DOUT0 => \N__7583\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12855\,
            DIN => \N__12854\,
            DOUT => \N__12853\,
            PACKAGEPIN => D_UU_AMIGA(0)
        );

    \D_UU_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12855\,
            PADOUT => \N__12854\,
            PADIN => \N__12853\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5375\,
            DIN0 => \D_UU_AMIGA_in_0\,
            DOUT0 => \N__9365\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12846\,
            DIN => \N__12845\,
            DOUT => \N__12844\,
            PACKAGEPIN => D_LL_040(4)
        );

    \D_LL_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12846\,
            PADOUT => \N__12845\,
            PADIN => \N__12844\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9842\,
            DIN0 => \D_LL_040_in_4\,
            DOUT0 => \N__5543\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12837\,
            DIN => \N__12836\,
            DOUT => \N__12835\,
            PACKAGEPIN => D_LL_AMIGA(7)
        );

    \D_LL_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12837\,
            PADOUT => \N__12836\,
            PADIN => \N__12835\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4112\,
            DIN0 => \D_LL_AMIGA_in_7\,
            DOUT0 => \N__8723\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12828\,
            DIN => \N__12827\,
            DOUT => \N__12826\,
            PACKAGEPIN => D_UU_040(4)
        );

    \D_UU_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12828\,
            PADOUT => \N__12827\,
            PADIN => \N__12826\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9614\,
            DIN0 => \D_UU_040_in_4\,
            DOUT0 => \N__8510\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12819\,
            DIN => \N__12818\,
            DOUT => \N__12817\,
            PACKAGEPIN => D_UM_AMIGA(5)
        );

    \D_UM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12819\,
            PADOUT => \N__12818\,
            PADIN => \N__12817\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5330\,
            DIN0 => \D_UM_AMIGA_in_5\,
            DOUT0 => \N__8012\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__3259\ : InMux
    port map (
            O => \N__12800\,
            I => \N__12797\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__12797\,
            I => \READ_CYCLE_ACTIVE_rep3_i_ess\
        );

    \I__3257\ : IoInMux
    port map (
            O => \N__12794\,
            I => \N__12791\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__12791\,
            I => \N__12788\
        );

    \I__3255\ : Span12Mux_s6_v
    port map (
            O => \N__12788\,
            I => \N__12785\
        );

    \I__3254\ : Odrv12
    port map (
            O => \N__12785\,
            I => \N_183_i\
        );

    \I__3253\ : InMux
    port map (
            O => \N__12782\,
            I => \N__12779\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__12779\,
            I => \READ_CYCLE_ACTIVE_rep9_i_ess\
        );

    \I__3251\ : IoInMux
    port map (
            O => \N__12776\,
            I => \N__12773\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__12773\,
            I => \N__12770\
        );

    \I__3249\ : Span4Mux_s3_h
    port map (
            O => \N__12770\,
            I => \N__12767\
        );

    \I__3248\ : Span4Mux_v
    port map (
            O => \N__12767\,
            I => \N__12764\
        );

    \I__3247\ : Odrv4
    port map (
            O => \N__12764\,
            I => \N_189_i\
        );

    \I__3246\ : InMux
    port map (
            O => \N__12761\,
            I => \N__12758\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__12758\,
            I => \READ_CYCLE_ACTIVE_rep11_i_ess\
        );

    \I__3244\ : IoInMux
    port map (
            O => \N__12755\,
            I => \N__12752\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__12752\,
            I => \N__12749\
        );

    \I__3242\ : Span4Mux_s3_h
    port map (
            O => \N__12749\,
            I => \N__12746\
        );

    \I__3241\ : Span4Mux_v
    port map (
            O => \N__12746\,
            I => \N__12743\
        );

    \I__3240\ : Odrv4
    port map (
            O => \N__12743\,
            I => \N_191_i\
        );

    \I__3239\ : InMux
    port map (
            O => \N__12740\,
            I => \N__12737\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__12737\,
            I => \READ_CYCLE_ACTIVE_rep15_i_ess\
        );

    \I__3237\ : IoInMux
    port map (
            O => \N__12734\,
            I => \N__12731\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__12731\,
            I => \N__12728\
        );

    \I__3235\ : Span12Mux_s4_h
    port map (
            O => \N__12728\,
            I => \N__12725\
        );

    \I__3234\ : Odrv12
    port map (
            O => \N__12725\,
            I => \N_195_i\
        );

    \I__3233\ : CascadeMux
    port map (
            O => \N__12722\,
            I => \N__12714\
        );

    \I__3232\ : CascadeMux
    port map (
            O => \N__12721\,
            I => \N__12710\
        );

    \I__3231\ : CascadeMux
    port map (
            O => \N__12720\,
            I => \N__12706\
        );

    \I__3230\ : CascadeMux
    port map (
            O => \N__12719\,
            I => \N__12701\
        );

    \I__3229\ : IoInMux
    port map (
            O => \N__12718\,
            I => \N__12696\
        );

    \I__3228\ : InMux
    port map (
            O => \N__12717\,
            I => \N__12690\
        );

    \I__3227\ : InMux
    port map (
            O => \N__12714\,
            I => \N__12686\
        );

    \I__3226\ : InMux
    port map (
            O => \N__12713\,
            I => \N__12683\
        );

    \I__3225\ : InMux
    port map (
            O => \N__12710\,
            I => \N__12680\
        );

    \I__3224\ : CascadeMux
    port map (
            O => \N__12709\,
            I => \N__12674\
        );

    \I__3223\ : InMux
    port map (
            O => \N__12706\,
            I => \N__12671\
        );

    \I__3222\ : InMux
    port map (
            O => \N__12705\,
            I => \N__12666\
        );

    \I__3221\ : CascadeMux
    port map (
            O => \N__12704\,
            I => \N__12663\
        );

    \I__3220\ : InMux
    port map (
            O => \N__12701\,
            I => \N__12660\
        );

    \I__3219\ : InMux
    port map (
            O => \N__12700\,
            I => \N__12655\
        );

    \I__3218\ : InMux
    port map (
            O => \N__12699\,
            I => \N__12655\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__12696\,
            I => \N__12652\
        );

    \I__3216\ : CascadeMux
    port map (
            O => \N__12695\,
            I => \N__12649\
        );

    \I__3215\ : CascadeMux
    port map (
            O => \N__12694\,
            I => \N__12646\
        );

    \I__3214\ : CascadeMux
    port map (
            O => \N__12693\,
            I => \N__12643\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__12690\,
            I => \N__12637\
        );

    \I__3212\ : InMux
    port map (
            O => \N__12689\,
            I => \N__12634\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__12686\,
            I => \N__12627\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__12683\,
            I => \N__12627\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__12680\,
            I => \N__12627\
        );

    \I__3208\ : InMux
    port map (
            O => \N__12679\,
            I => \N__12624\
        );

    \I__3207\ : InMux
    port map (
            O => \N__12678\,
            I => \N__12621\
        );

    \I__3206\ : CascadeMux
    port map (
            O => \N__12677\,
            I => \N__12617\
        );

    \I__3205\ : InMux
    port map (
            O => \N__12674\,
            I => \N__12614\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__12671\,
            I => \N__12611\
        );

    \I__3203\ : InMux
    port map (
            O => \N__12670\,
            I => \N__12608\
        );

    \I__3202\ : InMux
    port map (
            O => \N__12669\,
            I => \N__12605\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__12666\,
            I => \N__12600\
        );

    \I__3200\ : InMux
    port map (
            O => \N__12663\,
            I => \N__12597\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__12660\,
            I => \N__12586\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__12655\,
            I => \N__12586\
        );

    \I__3197\ : Span4Mux_s3_v
    port map (
            O => \N__12652\,
            I => \N__12583\
        );

    \I__3196\ : InMux
    port map (
            O => \N__12649\,
            I => \N__12580\
        );

    \I__3195\ : InMux
    port map (
            O => \N__12646\,
            I => \N__12575\
        );

    \I__3194\ : InMux
    port map (
            O => \N__12643\,
            I => \N__12575\
        );

    \I__3193\ : InMux
    port map (
            O => \N__12642\,
            I => \N__12570\
        );

    \I__3192\ : InMux
    port map (
            O => \N__12641\,
            I => \N__12570\
        );

    \I__3191\ : InMux
    port map (
            O => \N__12640\,
            I => \N__12567\
        );

    \I__3190\ : Span4Mux_h
    port map (
            O => \N__12637\,
            I => \N__12562\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__12634\,
            I => \N__12562\
        );

    \I__3188\ : Span4Mux_v
    port map (
            O => \N__12627\,
            I => \N__12557\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__12624\,
            I => \N__12557\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__12621\,
            I => \N__12554\
        );

    \I__3185\ : InMux
    port map (
            O => \N__12620\,
            I => \N__12551\
        );

    \I__3184\ : InMux
    port map (
            O => \N__12617\,
            I => \N__12548\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__12614\,
            I => \N__12541\
        );

    \I__3182\ : Span4Mux_h
    port map (
            O => \N__12611\,
            I => \N__12534\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__12608\,
            I => \N__12534\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__12605\,
            I => \N__12534\
        );

    \I__3179\ : InMux
    port map (
            O => \N__12604\,
            I => \N__12529\
        );

    \I__3178\ : InMux
    port map (
            O => \N__12603\,
            I => \N__12529\
        );

    \I__3177\ : Span4Mux_h
    port map (
            O => \N__12600\,
            I => \N__12521\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__12597\,
            I => \N__12521\
        );

    \I__3175\ : InMux
    port map (
            O => \N__12596\,
            I => \N__12516\
        );

    \I__3174\ : InMux
    port map (
            O => \N__12595\,
            I => \N__12516\
        );

    \I__3173\ : InMux
    port map (
            O => \N__12594\,
            I => \N__12509\
        );

    \I__3172\ : InMux
    port map (
            O => \N__12593\,
            I => \N__12509\
        );

    \I__3171\ : InMux
    port map (
            O => \N__12592\,
            I => \N__12509\
        );

    \I__3170\ : InMux
    port map (
            O => \N__12591\,
            I => \N__12506\
        );

    \I__3169\ : Span4Mux_v
    port map (
            O => \N__12586\,
            I => \N__12498\
        );

    \I__3168\ : Span4Mux_v
    port map (
            O => \N__12583\,
            I => \N__12487\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__12580\,
            I => \N__12487\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__12575\,
            I => \N__12487\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__12570\,
            I => \N__12487\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__12567\,
            I => \N__12487\
        );

    \I__3163\ : Span4Mux_v
    port map (
            O => \N__12562\,
            I => \N__12476\
        );

    \I__3162\ : Span4Mux_v
    port map (
            O => \N__12557\,
            I => \N__12476\
        );

    \I__3161\ : Span4Mux_v
    port map (
            O => \N__12554\,
            I => \N__12476\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__12551\,
            I => \N__12476\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__12548\,
            I => \N__12476\
        );

    \I__3158\ : InMux
    port map (
            O => \N__12547\,
            I => \N__12469\
        );

    \I__3157\ : InMux
    port map (
            O => \N__12546\,
            I => \N__12469\
        );

    \I__3156\ : InMux
    port map (
            O => \N__12545\,
            I => \N__12469\
        );

    \I__3155\ : CascadeMux
    port map (
            O => \N__12544\,
            I => \N__12464\
        );

    \I__3154\ : Span4Mux_v
    port map (
            O => \N__12541\,
            I => \N__12459\
        );

    \I__3153\ : Span4Mux_v
    port map (
            O => \N__12534\,
            I => \N__12459\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__12529\,
            I => \N__12456\
        );

    \I__3151\ : InMux
    port map (
            O => \N__12528\,
            I => \N__12453\
        );

    \I__3150\ : InMux
    port map (
            O => \N__12527\,
            I => \N__12449\
        );

    \I__3149\ : InMux
    port map (
            O => \N__12526\,
            I => \N__12446\
        );

    \I__3148\ : Span4Mux_h
    port map (
            O => \N__12521\,
            I => \N__12434\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__12516\,
            I => \N__12434\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__12509\,
            I => \N__12434\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__12506\,
            I => \N__12434\
        );

    \I__3144\ : InMux
    port map (
            O => \N__12505\,
            I => \N__12431\
        );

    \I__3143\ : CascadeMux
    port map (
            O => \N__12504\,
            I => \N__12427\
        );

    \I__3142\ : CascadeMux
    port map (
            O => \N__12503\,
            I => \N__12423\
        );

    \I__3141\ : CascadeMux
    port map (
            O => \N__12502\,
            I => \N__12420\
        );

    \I__3140\ : CascadeMux
    port map (
            O => \N__12501\,
            I => \N__12416\
        );

    \I__3139\ : Span4Mux_v
    port map (
            O => \N__12498\,
            I => \N__12407\
        );

    \I__3138\ : Span4Mux_v
    port map (
            O => \N__12487\,
            I => \N__12402\
        );

    \I__3137\ : Span4Mux_v
    port map (
            O => \N__12476\,
            I => \N__12402\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__12469\,
            I => \N__12399\
        );

    \I__3135\ : InMux
    port map (
            O => \N__12468\,
            I => \N__12392\
        );

    \I__3134\ : InMux
    port map (
            O => \N__12467\,
            I => \N__12392\
        );

    \I__3133\ : InMux
    port map (
            O => \N__12464\,
            I => \N__12392\
        );

    \I__3132\ : Span4Mux_h
    port map (
            O => \N__12459\,
            I => \N__12385\
        );

    \I__3131\ : Span4Mux_h
    port map (
            O => \N__12456\,
            I => \N__12385\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__12453\,
            I => \N__12385\
        );

    \I__3129\ : InMux
    port map (
            O => \N__12452\,
            I => \N__12382\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__12449\,
            I => \N__12379\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__12446\,
            I => \N__12376\
        );

    \I__3126\ : InMux
    port map (
            O => \N__12445\,
            I => \N__12371\
        );

    \I__3125\ : InMux
    port map (
            O => \N__12444\,
            I => \N__12371\
        );

    \I__3124\ : InMux
    port map (
            O => \N__12443\,
            I => \N__12368\
        );

    \I__3123\ : Span4Mux_v
    port map (
            O => \N__12434\,
            I => \N__12365\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__12431\,
            I => \N__12362\
        );

    \I__3121\ : InMux
    port map (
            O => \N__12430\,
            I => \N__12359\
        );

    \I__3120\ : InMux
    port map (
            O => \N__12427\,
            I => \N__12356\
        );

    \I__3119\ : InMux
    port map (
            O => \N__12426\,
            I => \N__12345\
        );

    \I__3118\ : InMux
    port map (
            O => \N__12423\,
            I => \N__12345\
        );

    \I__3117\ : InMux
    port map (
            O => \N__12420\,
            I => \N__12345\
        );

    \I__3116\ : InMux
    port map (
            O => \N__12419\,
            I => \N__12345\
        );

    \I__3115\ : InMux
    port map (
            O => \N__12416\,
            I => \N__12345\
        );

    \I__3114\ : InMux
    port map (
            O => \N__12415\,
            I => \N__12342\
        );

    \I__3113\ : InMux
    port map (
            O => \N__12414\,
            I => \N__12339\
        );

    \I__3112\ : CascadeMux
    port map (
            O => \N__12413\,
            I => \N__12331\
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__12412\,
            I => \N__12328\
        );

    \I__3110\ : CascadeMux
    port map (
            O => \N__12411\,
            I => \N__12324\
        );

    \I__3109\ : CascadeMux
    port map (
            O => \N__12410\,
            I => \N__12321\
        );

    \I__3108\ : Sp12to4
    port map (
            O => \N__12407\,
            I => \N__12316\
        );

    \I__3107\ : Sp12to4
    port map (
            O => \N__12402\,
            I => \N__12316\
        );

    \I__3106\ : Span12Mux_s11_h
    port map (
            O => \N__12399\,
            I => \N__12313\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__12392\,
            I => \N__12310\
        );

    \I__3104\ : Sp12to4
    port map (
            O => \N__12385\,
            I => \N__12305\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__12382\,
            I => \N__12305\
        );

    \I__3102\ : Span4Mux_v
    port map (
            O => \N__12379\,
            I => \N__12302\
        );

    \I__3101\ : Span4Mux_h
    port map (
            O => \N__12376\,
            I => \N__12295\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__12371\,
            I => \N__12295\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__12368\,
            I => \N__12295\
        );

    \I__3098\ : Span4Mux_v
    port map (
            O => \N__12365\,
            I => \N__12292\
        );

    \I__3097\ : Span4Mux_h
    port map (
            O => \N__12362\,
            I => \N__12285\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__12359\,
            I => \N__12285\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__12356\,
            I => \N__12285\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__12345\,
            I => \N__12280\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__12342\,
            I => \N__12280\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__12339\,
            I => \N__12277\
        );

    \I__3091\ : InMux
    port map (
            O => \N__12338\,
            I => \N__12270\
        );

    \I__3090\ : InMux
    port map (
            O => \N__12337\,
            I => \N__12270\
        );

    \I__3089\ : InMux
    port map (
            O => \N__12336\,
            I => \N__12270\
        );

    \I__3088\ : InMux
    port map (
            O => \N__12335\,
            I => \N__12263\
        );

    \I__3087\ : InMux
    port map (
            O => \N__12334\,
            I => \N__12263\
        );

    \I__3086\ : InMux
    port map (
            O => \N__12331\,
            I => \N__12263\
        );

    \I__3085\ : InMux
    port map (
            O => \N__12328\,
            I => \N__12254\
        );

    \I__3084\ : InMux
    port map (
            O => \N__12327\,
            I => \N__12254\
        );

    \I__3083\ : InMux
    port map (
            O => \N__12324\,
            I => \N__12254\
        );

    \I__3082\ : InMux
    port map (
            O => \N__12321\,
            I => \N__12254\
        );

    \I__3081\ : Span12Mux_h
    port map (
            O => \N__12316\,
            I => \N__12251\
        );

    \I__3080\ : Span12Mux_h
    port map (
            O => \N__12313\,
            I => \N__12248\
        );

    \I__3079\ : Span12Mux_s11_h
    port map (
            O => \N__12310\,
            I => \N__12241\
        );

    \I__3078\ : Span12Mux_s11_v
    port map (
            O => \N__12305\,
            I => \N__12241\
        );

    \I__3077\ : Sp12to4
    port map (
            O => \N__12302\,
            I => \N__12241\
        );

    \I__3076\ : Span4Mux_v
    port map (
            O => \N__12295\,
            I => \N__12238\
        );

    \I__3075\ : Span4Mux_v
    port map (
            O => \N__12292\,
            I => \N__12233\
        );

    \I__3074\ : Span4Mux_v
    port map (
            O => \N__12285\,
            I => \N__12233\
        );

    \I__3073\ : Span4Mux_v
    port map (
            O => \N__12280\,
            I => \N__12228\
        );

    \I__3072\ : Span4Mux_v
    port map (
            O => \N__12277\,
            I => \N__12228\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__12270\,
            I => \N__12225\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__12263\,
            I => \N__12222\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__12254\,
            I => \N__12219\
        );

    \I__3068\ : Span12Mux_h
    port map (
            O => \N__12251\,
            I => \N__12216\
        );

    \I__3067\ : Span12Mux_v
    port map (
            O => \N__12248\,
            I => \N__12211\
        );

    \I__3066\ : Span12Mux_h
    port map (
            O => \N__12241\,
            I => \N__12211\
        );

    \I__3065\ : Span4Mux_h
    port map (
            O => \N__12238\,
            I => \N__12208\
        );

    \I__3064\ : Span4Mux_h
    port map (
            O => \N__12233\,
            I => \N__12205\
        );

    \I__3063\ : Span4Mux_v
    port map (
            O => \N__12228\,
            I => \N__12196\
        );

    \I__3062\ : Span4Mux_v
    port map (
            O => \N__12225\,
            I => \N__12196\
        );

    \I__3061\ : Span4Mux_v
    port map (
            O => \N__12222\,
            I => \N__12196\
        );

    \I__3060\ : Span4Mux_v
    port map (
            O => \N__12219\,
            I => \N__12196\
        );

    \I__3059\ : Odrv12
    port map (
            O => \N__12216\,
            I => \RnW_c\
        );

    \I__3058\ : Odrv12
    port map (
            O => \N__12211\,
            I => \RnW_c\
        );

    \I__3057\ : Odrv4
    port map (
            O => \N__12208\,
            I => \RnW_c\
        );

    \I__3056\ : Odrv4
    port map (
            O => \N__12205\,
            I => \RnW_c\
        );

    \I__3055\ : Odrv4
    port map (
            O => \N__12196\,
            I => \RnW_c\
        );

    \I__3054\ : CascadeMux
    port map (
            O => \N__12185\,
            I => \N__12180\
        );

    \I__3053\ : CascadeMux
    port map (
            O => \N__12184\,
            I => \N__12177\
        );

    \I__3052\ : InMux
    port map (
            O => \N__12183\,
            I => \N__12172\
        );

    \I__3051\ : InMux
    port map (
            O => \N__12180\,
            I => \N__12172\
        );

    \I__3050\ : InMux
    port map (
            O => \N__12177\,
            I => \N__12169\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__12172\,
            I => \N__12157\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__12169\,
            I => \N__12157\
        );

    \I__3047\ : InMux
    port map (
            O => \N__12168\,
            I => \N__12154\
        );

    \I__3046\ : InMux
    port map (
            O => \N__12167\,
            I => \N__12151\
        );

    \I__3045\ : InMux
    port map (
            O => \N__12166\,
            I => \N__12148\
        );

    \I__3044\ : InMux
    port map (
            O => \N__12165\,
            I => \N__12145\
        );

    \I__3043\ : CascadeMux
    port map (
            O => \N__12164\,
            I => \N__12141\
        );

    \I__3042\ : CascadeMux
    port map (
            O => \N__12163\,
            I => \N__12138\
        );

    \I__3041\ : CascadeMux
    port map (
            O => \N__12162\,
            I => \N__12128\
        );

    \I__3040\ : Span4Mux_h
    port map (
            O => \N__12157\,
            I => \N__12119\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__12154\,
            I => \N__12119\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__12151\,
            I => \N__12119\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__12148\,
            I => \N__12119\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__12145\,
            I => \N__12116\
        );

    \I__3035\ : InMux
    port map (
            O => \N__12144\,
            I => \N__12113\
        );

    \I__3034\ : InMux
    port map (
            O => \N__12141\,
            I => \N__12110\
        );

    \I__3033\ : InMux
    port map (
            O => \N__12138\,
            I => \N__12107\
        );

    \I__3032\ : InMux
    port map (
            O => \N__12137\,
            I => \N__12103\
        );

    \I__3031\ : CascadeMux
    port map (
            O => \N__12136\,
            I => \N__12100\
        );

    \I__3030\ : InMux
    port map (
            O => \N__12135\,
            I => \N__12089\
        );

    \I__3029\ : InMux
    port map (
            O => \N__12134\,
            I => \N__12089\
        );

    \I__3028\ : InMux
    port map (
            O => \N__12133\,
            I => \N__12085\
        );

    \I__3027\ : InMux
    port map (
            O => \N__12132\,
            I => \N__12082\
        );

    \I__3026\ : InMux
    port map (
            O => \N__12131\,
            I => \N__12077\
        );

    \I__3025\ : InMux
    port map (
            O => \N__12128\,
            I => \N__12077\
        );

    \I__3024\ : Span4Mux_v
    port map (
            O => \N__12119\,
            I => \N__12058\
        );

    \I__3023\ : Span4Mux_h
    port map (
            O => \N__12116\,
            I => \N__12058\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__12113\,
            I => \N__12058\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__12110\,
            I => \N__12058\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__12107\,
            I => \N__12058\
        );

    \I__3019\ : InMux
    port map (
            O => \N__12106\,
            I => \N__12055\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__12103\,
            I => \N__12052\
        );

    \I__3017\ : InMux
    port map (
            O => \N__12100\,
            I => \N__12049\
        );

    \I__3016\ : InMux
    port map (
            O => \N__12099\,
            I => \N__12046\
        );

    \I__3015\ : InMux
    port map (
            O => \N__12098\,
            I => \N__12039\
        );

    \I__3014\ : InMux
    port map (
            O => \N__12097\,
            I => \N__12039\
        );

    \I__3013\ : InMux
    port map (
            O => \N__12096\,
            I => \N__12039\
        );

    \I__3012\ : CascadeMux
    port map (
            O => \N__12095\,
            I => \N__12036\
        );

    \I__3011\ : CascadeMux
    port map (
            O => \N__12094\,
            I => \N__12026\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__12089\,
            I => \N__12023\
        );

    \I__3009\ : InMux
    port map (
            O => \N__12088\,
            I => \N__12020\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__12085\,
            I => \N__12012\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__12082\,
            I => \N__12012\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__12077\,
            I => \N__12012\
        );

    \I__3005\ : InMux
    port map (
            O => \N__12076\,
            I => \N__12009\
        );

    \I__3004\ : InMux
    port map (
            O => \N__12075\,
            I => \N__11998\
        );

    \I__3003\ : InMux
    port map (
            O => \N__12074\,
            I => \N__11998\
        );

    \I__3002\ : InMux
    port map (
            O => \N__12073\,
            I => \N__11998\
        );

    \I__3001\ : InMux
    port map (
            O => \N__12072\,
            I => \N__11998\
        );

    \I__3000\ : InMux
    port map (
            O => \N__12071\,
            I => \N__11998\
        );

    \I__2999\ : CascadeMux
    port map (
            O => \N__12070\,
            I => \N__11995\
        );

    \I__2998\ : CascadeMux
    port map (
            O => \N__12069\,
            I => \N__11992\
        );

    \I__2997\ : Span4Mux_v
    port map (
            O => \N__12058\,
            I => \N__11983\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__12055\,
            I => \N__11983\
        );

    \I__2995\ : Span4Mux_h
    port map (
            O => \N__12052\,
            I => \N__11976\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__12049\,
            I => \N__11976\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__12046\,
            I => \N__11976\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__12039\,
            I => \N__11973\
        );

    \I__2991\ : InMux
    port map (
            O => \N__12036\,
            I => \N__11970\
        );

    \I__2990\ : InMux
    port map (
            O => \N__12035\,
            I => \N__11965\
        );

    \I__2989\ : InMux
    port map (
            O => \N__12034\,
            I => \N__11965\
        );

    \I__2988\ : InMux
    port map (
            O => \N__12033\,
            I => \N__11962\
        );

    \I__2987\ : InMux
    port map (
            O => \N__12032\,
            I => \N__11959\
        );

    \I__2986\ : CascadeMux
    port map (
            O => \N__12031\,
            I => \N__11954\
        );

    \I__2985\ : CascadeMux
    port map (
            O => \N__12030\,
            I => \N__11949\
        );

    \I__2984\ : CascadeMux
    port map (
            O => \N__12029\,
            I => \N__11946\
        );

    \I__2983\ : InMux
    port map (
            O => \N__12026\,
            I => \N__11939\
        );

    \I__2982\ : Span4Mux_h
    port map (
            O => \N__12023\,
            I => \N__11936\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__12020\,
            I => \N__11933\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__12019\,
            I => \N__11929\
        );

    \I__2979\ : Span4Mux_v
    port map (
            O => \N__12012\,
            I => \N__11924\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__12009\,
            I => \N__11924\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__11998\,
            I => \N__11921\
        );

    \I__2976\ : InMux
    port map (
            O => \N__11995\,
            I => \N__11918\
        );

    \I__2975\ : InMux
    port map (
            O => \N__11992\,
            I => \N__11915\
        );

    \I__2974\ : CascadeMux
    port map (
            O => \N__11991\,
            I => \N__11909\
        );

    \I__2973\ : CascadeMux
    port map (
            O => \N__11990\,
            I => \N__11906\
        );

    \I__2972\ : CascadeMux
    port map (
            O => \N__11989\,
            I => \N__11902\
        );

    \I__2971\ : CascadeMux
    port map (
            O => \N__11988\,
            I => \N__11899\
        );

    \I__2970\ : Span4Mux_v
    port map (
            O => \N__11983\,
            I => \N__11884\
        );

    \I__2969\ : Span4Mux_v
    port map (
            O => \N__11976\,
            I => \N__11884\
        );

    \I__2968\ : Span4Mux_h
    port map (
            O => \N__11973\,
            I => \N__11884\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__11970\,
            I => \N__11884\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__11965\,
            I => \N__11884\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__11962\,
            I => \N__11884\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__11959\,
            I => \N__11884\
        );

    \I__2963\ : InMux
    port map (
            O => \N__11958\,
            I => \N__11879\
        );

    \I__2962\ : InMux
    port map (
            O => \N__11957\,
            I => \N__11879\
        );

    \I__2961\ : InMux
    port map (
            O => \N__11954\,
            I => \N__11876\
        );

    \I__2960\ : InMux
    port map (
            O => \N__11953\,
            I => \N__11872\
        );

    \I__2959\ : InMux
    port map (
            O => \N__11952\,
            I => \N__11865\
        );

    \I__2958\ : InMux
    port map (
            O => \N__11949\,
            I => \N__11865\
        );

    \I__2957\ : InMux
    port map (
            O => \N__11946\,
            I => \N__11865\
        );

    \I__2956\ : InMux
    port map (
            O => \N__11945\,
            I => \N__11862\
        );

    \I__2955\ : CascadeMux
    port map (
            O => \N__11944\,
            I => \N__11859\
        );

    \I__2954\ : CascadeMux
    port map (
            O => \N__11943\,
            I => \N__11856\
        );

    \I__2953\ : CascadeMux
    port map (
            O => \N__11942\,
            I => \N__11853\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__11939\,
            I => \N__11850\
        );

    \I__2951\ : Span4Mux_v
    port map (
            O => \N__11936\,
            I => \N__11845\
        );

    \I__2950\ : Span4Mux_h
    port map (
            O => \N__11933\,
            I => \N__11845\
        );

    \I__2949\ : CascadeMux
    port map (
            O => \N__11932\,
            I => \N__11842\
        );

    \I__2948\ : InMux
    port map (
            O => \N__11929\,
            I => \N__11839\
        );

    \I__2947\ : Span4Mux_v
    port map (
            O => \N__11924\,
            I => \N__11830\
        );

    \I__2946\ : Span4Mux_v
    port map (
            O => \N__11921\,
            I => \N__11830\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__11918\,
            I => \N__11830\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__11915\,
            I => \N__11830\
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__11914\,
            I => \N__11826\
        );

    \I__2942\ : CascadeMux
    port map (
            O => \N__11913\,
            I => \N__11821\
        );

    \I__2941\ : CascadeMux
    port map (
            O => \N__11912\,
            I => \N__11818\
        );

    \I__2940\ : InMux
    port map (
            O => \N__11909\,
            I => \N__11811\
        );

    \I__2939\ : InMux
    port map (
            O => \N__11906\,
            I => \N__11811\
        );

    \I__2938\ : InMux
    port map (
            O => \N__11905\,
            I => \N__11804\
        );

    \I__2937\ : InMux
    port map (
            O => \N__11902\,
            I => \N__11804\
        );

    \I__2936\ : InMux
    port map (
            O => \N__11899\,
            I => \N__11804\
        );

    \I__2935\ : Span4Mux_v
    port map (
            O => \N__11884\,
            I => \N__11799\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__11879\,
            I => \N__11799\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__11876\,
            I => \N__11796\
        );

    \I__2932\ : InMux
    port map (
            O => \N__11875\,
            I => \N__11793\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__11872\,
            I => \N__11790\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__11865\,
            I => \N__11785\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__11862\,
            I => \N__11785\
        );

    \I__2928\ : InMux
    port map (
            O => \N__11859\,
            I => \N__11780\
        );

    \I__2927\ : InMux
    port map (
            O => \N__11856\,
            I => \N__11780\
        );

    \I__2926\ : InMux
    port map (
            O => \N__11853\,
            I => \N__11777\
        );

    \I__2925\ : Span4Mux_h
    port map (
            O => \N__11850\,
            I => \N__11772\
        );

    \I__2924\ : Span4Mux_v
    port map (
            O => \N__11845\,
            I => \N__11772\
        );

    \I__2923\ : InMux
    port map (
            O => \N__11842\,
            I => \N__11769\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__11839\,
            I => \N__11766\
        );

    \I__2921\ : Span4Mux_v
    port map (
            O => \N__11830\,
            I => \N__11763\
        );

    \I__2920\ : InMux
    port map (
            O => \N__11829\,
            I => \N__11754\
        );

    \I__2919\ : InMux
    port map (
            O => \N__11826\,
            I => \N__11754\
        );

    \I__2918\ : InMux
    port map (
            O => \N__11825\,
            I => \N__11754\
        );

    \I__2917\ : InMux
    port map (
            O => \N__11824\,
            I => \N__11754\
        );

    \I__2916\ : InMux
    port map (
            O => \N__11821\,
            I => \N__11747\
        );

    \I__2915\ : InMux
    port map (
            O => \N__11818\,
            I => \N__11747\
        );

    \I__2914\ : InMux
    port map (
            O => \N__11817\,
            I => \N__11747\
        );

    \I__2913\ : CascadeMux
    port map (
            O => \N__11816\,
            I => \N__11743\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__11811\,
            I => \N__11737\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__11804\,
            I => \N__11737\
        );

    \I__2910\ : Span4Mux_h
    port map (
            O => \N__11799\,
            I => \N__11730\
        );

    \I__2909\ : Span4Mux_v
    port map (
            O => \N__11796\,
            I => \N__11730\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__11793\,
            I => \N__11730\
        );

    \I__2907\ : Span4Mux_v
    port map (
            O => \N__11790\,
            I => \N__11721\
        );

    \I__2906\ : Span4Mux_h
    port map (
            O => \N__11785\,
            I => \N__11721\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__11780\,
            I => \N__11721\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__11777\,
            I => \N__11721\
        );

    \I__2903\ : Span4Mux_h
    port map (
            O => \N__11772\,
            I => \N__11716\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__11769\,
            I => \N__11716\
        );

    \I__2901\ : Span12Mux_h
    port map (
            O => \N__11766\,
            I => \N__11709\
        );

    \I__2900\ : Sp12to4
    port map (
            O => \N__11763\,
            I => \N__11709\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__11754\,
            I => \N__11709\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__11747\,
            I => \N__11706\
        );

    \I__2897\ : InMux
    port map (
            O => \N__11746\,
            I => \N__11703\
        );

    \I__2896\ : InMux
    port map (
            O => \N__11743\,
            I => \N__11698\
        );

    \I__2895\ : InMux
    port map (
            O => \N__11742\,
            I => \N__11698\
        );

    \I__2894\ : Span4Mux_v
    port map (
            O => \N__11737\,
            I => \N__11695\
        );

    \I__2893\ : Span4Mux_h
    port map (
            O => \N__11730\,
            I => \N__11692\
        );

    \I__2892\ : Span4Mux_h
    port map (
            O => \N__11721\,
            I => \N__11689\
        );

    \I__2891\ : Span4Mux_v
    port map (
            O => \N__11716\,
            I => \N__11686\
        );

    \I__2890\ : Span12Mux_h
    port map (
            O => \N__11709\,
            I => \N__11683\
        );

    \I__2889\ : Span12Mux_h
    port map (
            O => \N__11706\,
            I => \N__11680\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__11703\,
            I => \N__11675\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__11698\,
            I => \N__11675\
        );

    \I__2886\ : Sp12to4
    port map (
            O => \N__11695\,
            I => \N__11672\
        );

    \I__2885\ : Span4Mux_v
    port map (
            O => \N__11692\,
            I => \N__11669\
        );

    \I__2884\ : Span4Mux_v
    port map (
            O => \N__11689\,
            I => \N__11666\
        );

    \I__2883\ : Span4Mux_v
    port map (
            O => \N__11686\,
            I => \N__11663\
        );

    \I__2882\ : Span12Mux_v
    port map (
            O => \N__11683\,
            I => \N__11660\
        );

    \I__2881\ : Span12Mux_v
    port map (
            O => \N__11680\,
            I => \N__11655\
        );

    \I__2880\ : Span12Mux_h
    port map (
            O => \N__11675\,
            I => \N__11655\
        );

    \I__2879\ : Span12Mux_h
    port map (
            O => \N__11672\,
            I => \N__11652\
        );

    \I__2878\ : Span4Mux_h
    port map (
            O => \N__11669\,
            I => \N__11647\
        );

    \I__2877\ : Span4Mux_h
    port map (
            O => \N__11666\,
            I => \N__11647\
        );

    \I__2876\ : IoSpan4Mux
    port map (
            O => \N__11663\,
            I => \N__11644\
        );

    \I__2875\ : Odrv12
    port map (
            O => \N__11660\,
            I => \TS_CPUn_c\
        );

    \I__2874\ : Odrv12
    port map (
            O => \N__11655\,
            I => \TS_CPUn_c\
        );

    \I__2873\ : Odrv12
    port map (
            O => \N__11652\,
            I => \TS_CPUn_c\
        );

    \I__2872\ : Odrv4
    port map (
            O => \N__11647\,
            I => \TS_CPUn_c\
        );

    \I__2871\ : Odrv4
    port map (
            O => \N__11644\,
            I => \TS_CPUn_c\
        );

    \I__2870\ : InMux
    port map (
            O => \N__11633\,
            I => \N__11626\
        );

    \I__2869\ : InMux
    port map (
            O => \N__11632\,
            I => \N__11621\
        );

    \I__2868\ : InMux
    port map (
            O => \N__11631\,
            I => \N__11621\
        );

    \I__2867\ : CascadeMux
    port map (
            O => \N__11630\,
            I => \N__11612\
        );

    \I__2866\ : CascadeMux
    port map (
            O => \N__11629\,
            I => \N__11609\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__11626\,
            I => \N__11601\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__11621\,
            I => \N__11601\
        );

    \I__2863\ : InMux
    port map (
            O => \N__11620\,
            I => \N__11596\
        );

    \I__2862\ : InMux
    port map (
            O => \N__11619\,
            I => \N__11596\
        );

    \I__2861\ : CascadeMux
    port map (
            O => \N__11618\,
            I => \N__11593\
        );

    \I__2860\ : InMux
    port map (
            O => \N__11617\,
            I => \N__11590\
        );

    \I__2859\ : InMux
    port map (
            O => \N__11616\,
            I => \N__11585\
        );

    \I__2858\ : InMux
    port map (
            O => \N__11615\,
            I => \N__11585\
        );

    \I__2857\ : InMux
    port map (
            O => \N__11612\,
            I => \N__11580\
        );

    \I__2856\ : InMux
    port map (
            O => \N__11609\,
            I => \N__11580\
        );

    \I__2855\ : InMux
    port map (
            O => \N__11608\,
            I => \N__11577\
        );

    \I__2854\ : InMux
    port map (
            O => \N__11607\,
            I => \N__11574\
        );

    \I__2853\ : CascadeMux
    port map (
            O => \N__11606\,
            I => \N__11567\
        );

    \I__2852\ : Span4Mux_v
    port map (
            O => \N__11601\,
            I => \N__11558\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__11596\,
            I => \N__11558\
        );

    \I__2850\ : InMux
    port map (
            O => \N__11593\,
            I => \N__11555\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__11590\,
            I => \N__11545\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__11585\,
            I => \N__11536\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__11580\,
            I => \N__11536\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__11577\,
            I => \N__11536\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__11574\,
            I => \N__11536\
        );

    \I__2844\ : InMux
    port map (
            O => \N__11573\,
            I => \N__11529\
        );

    \I__2843\ : InMux
    port map (
            O => \N__11572\,
            I => \N__11529\
        );

    \I__2842\ : InMux
    port map (
            O => \N__11571\,
            I => \N__11529\
        );

    \I__2841\ : InMux
    port map (
            O => \N__11570\,
            I => \N__11526\
        );

    \I__2840\ : InMux
    port map (
            O => \N__11567\,
            I => \N__11523\
        );

    \I__2839\ : InMux
    port map (
            O => \N__11566\,
            I => \N__11520\
        );

    \I__2838\ : InMux
    port map (
            O => \N__11565\,
            I => \N__11517\
        );

    \I__2837\ : CascadeMux
    port map (
            O => \N__11564\,
            I => \N__11511\
        );

    \I__2836\ : InMux
    port map (
            O => \N__11563\,
            I => \N__11506\
        );

    \I__2835\ : Span4Mux_h
    port map (
            O => \N__11558\,
            I => \N__11498\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__11555\,
            I => \N__11498\
        );

    \I__2833\ : InMux
    port map (
            O => \N__11554\,
            I => \N__11495\
        );

    \I__2832\ : CascadeMux
    port map (
            O => \N__11553\,
            I => \N__11492\
        );

    \I__2831\ : CascadeMux
    port map (
            O => \N__11552\,
            I => \N__11489\
        );

    \I__2830\ : CascadeMux
    port map (
            O => \N__11551\,
            I => \N__11484\
        );

    \I__2829\ : CascadeMux
    port map (
            O => \N__11550\,
            I => \N__11479\
        );

    \I__2828\ : CascadeMux
    port map (
            O => \N__11549\,
            I => \N__11469\
        );

    \I__2827\ : CascadeMux
    port map (
            O => \N__11548\,
            I => \N__11466\
        );

    \I__2826\ : Span4Mux_v
    port map (
            O => \N__11545\,
            I => \N__11450\
        );

    \I__2825\ : Span4Mux_v
    port map (
            O => \N__11536\,
            I => \N__11450\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__11529\,
            I => \N__11450\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__11526\,
            I => \N__11450\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__11523\,
            I => \N__11450\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__11520\,
            I => \N__11450\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__11517\,
            I => \N__11450\
        );

    \I__2819\ : InMux
    port map (
            O => \N__11516\,
            I => \N__11447\
        );

    \I__2818\ : InMux
    port map (
            O => \N__11515\,
            I => \N__11444\
        );

    \I__2817\ : InMux
    port map (
            O => \N__11514\,
            I => \N__11441\
        );

    \I__2816\ : InMux
    port map (
            O => \N__11511\,
            I => \N__11438\
        );

    \I__2815\ : CascadeMux
    port map (
            O => \N__11510\,
            I => \N__11435\
        );

    \I__2814\ : CascadeMux
    port map (
            O => \N__11509\,
            I => \N__11431\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__11506\,
            I => \N__11427\
        );

    \I__2812\ : InMux
    port map (
            O => \N__11505\,
            I => \N__11424\
        );

    \I__2811\ : InMux
    port map (
            O => \N__11504\,
            I => \N__11421\
        );

    \I__2810\ : InMux
    port map (
            O => \N__11503\,
            I => \N__11418\
        );

    \I__2809\ : Span4Mux_v
    port map (
            O => \N__11498\,
            I => \N__11415\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__11495\,
            I => \N__11412\
        );

    \I__2807\ : InMux
    port map (
            O => \N__11492\,
            I => \N__11409\
        );

    \I__2806\ : InMux
    port map (
            O => \N__11489\,
            I => \N__11401\
        );

    \I__2805\ : InMux
    port map (
            O => \N__11488\,
            I => \N__11401\
        );

    \I__2804\ : InMux
    port map (
            O => \N__11487\,
            I => \N__11401\
        );

    \I__2803\ : InMux
    port map (
            O => \N__11484\,
            I => \N__11398\
        );

    \I__2802\ : InMux
    port map (
            O => \N__11483\,
            I => \N__11393\
        );

    \I__2801\ : InMux
    port map (
            O => \N__11482\,
            I => \N__11393\
        );

    \I__2800\ : InMux
    port map (
            O => \N__11479\,
            I => \N__11390\
        );

    \I__2799\ : InMux
    port map (
            O => \N__11478\,
            I => \N__11385\
        );

    \I__2798\ : InMux
    port map (
            O => \N__11477\,
            I => \N__11385\
        );

    \I__2797\ : InMux
    port map (
            O => \N__11476\,
            I => \N__11382\
        );

    \I__2796\ : InMux
    port map (
            O => \N__11475\,
            I => \N__11379\
        );

    \I__2795\ : CascadeMux
    port map (
            O => \N__11474\,
            I => \N__11370\
        );

    \I__2794\ : CascadeMux
    port map (
            O => \N__11473\,
            I => \N__11365\
        );

    \I__2793\ : CascadeMux
    port map (
            O => \N__11472\,
            I => \N__11359\
        );

    \I__2792\ : InMux
    port map (
            O => \N__11469\,
            I => \N__11355\
        );

    \I__2791\ : InMux
    port map (
            O => \N__11466\,
            I => \N__11350\
        );

    \I__2790\ : InMux
    port map (
            O => \N__11465\,
            I => \N__11350\
        );

    \I__2789\ : Span4Mux_v
    port map (
            O => \N__11450\,
            I => \N__11338\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__11447\,
            I => \N__11338\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__11444\,
            I => \N__11338\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__11441\,
            I => \N__11338\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__11438\,
            I => \N__11338\
        );

    \I__2784\ : InMux
    port map (
            O => \N__11435\,
            I => \N__11335\
        );

    \I__2783\ : InMux
    port map (
            O => \N__11434\,
            I => \N__11332\
        );

    \I__2782\ : InMux
    port map (
            O => \N__11431\,
            I => \N__11329\
        );

    \I__2781\ : InMux
    port map (
            O => \N__11430\,
            I => \N__11326\
        );

    \I__2780\ : Span4Mux_v
    port map (
            O => \N__11427\,
            I => \N__11321\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__11424\,
            I => \N__11321\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__11421\,
            I => \N__11316\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__11418\,
            I => \N__11316\
        );

    \I__2776\ : Span4Mux_h
    port map (
            O => \N__11415\,
            I => \N__11309\
        );

    \I__2775\ : Span4Mux_v
    port map (
            O => \N__11412\,
            I => \N__11309\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__11409\,
            I => \N__11309\
        );

    \I__2773\ : CascadeMux
    port map (
            O => \N__11408\,
            I => \N__11305\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__11401\,
            I => \N__11298\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__11398\,
            I => \N__11298\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__11393\,
            I => \N__11298\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__11390\,
            I => \N__11289\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__11385\,
            I => \N__11289\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__11382\,
            I => \N__11289\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__11379\,
            I => \N__11289\
        );

    \I__2765\ : InMux
    port map (
            O => \N__11378\,
            I => \N__11280\
        );

    \I__2764\ : InMux
    port map (
            O => \N__11377\,
            I => \N__11280\
        );

    \I__2763\ : InMux
    port map (
            O => \N__11376\,
            I => \N__11280\
        );

    \I__2762\ : InMux
    port map (
            O => \N__11375\,
            I => \N__11280\
        );

    \I__2761\ : InMux
    port map (
            O => \N__11374\,
            I => \N__11275\
        );

    \I__2760\ : InMux
    port map (
            O => \N__11373\,
            I => \N__11275\
        );

    \I__2759\ : InMux
    port map (
            O => \N__11370\,
            I => \N__11264\
        );

    \I__2758\ : InMux
    port map (
            O => \N__11369\,
            I => \N__11264\
        );

    \I__2757\ : InMux
    port map (
            O => \N__11368\,
            I => \N__11264\
        );

    \I__2756\ : InMux
    port map (
            O => \N__11365\,
            I => \N__11264\
        );

    \I__2755\ : InMux
    port map (
            O => \N__11364\,
            I => \N__11264\
        );

    \I__2754\ : InMux
    port map (
            O => \N__11363\,
            I => \N__11257\
        );

    \I__2753\ : InMux
    port map (
            O => \N__11362\,
            I => \N__11257\
        );

    \I__2752\ : InMux
    port map (
            O => \N__11359\,
            I => \N__11257\
        );

    \I__2751\ : InMux
    port map (
            O => \N__11358\,
            I => \N__11254\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__11355\,
            I => \N__11249\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__11350\,
            I => \N__11249\
        );

    \I__2748\ : CascadeMux
    port map (
            O => \N__11349\,
            I => \N__11246\
        );

    \I__2747\ : Span4Mux_v
    port map (
            O => \N__11338\,
            I => \N__11241\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__11335\,
            I => \N__11241\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__11332\,
            I => \N__11234\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__11329\,
            I => \N__11234\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__11326\,
            I => \N__11234\
        );

    \I__2742\ : Span4Mux_v
    port map (
            O => \N__11321\,
            I => \N__11228\
        );

    \I__2741\ : Span4Mux_v
    port map (
            O => \N__11316\,
            I => \N__11225\
        );

    \I__2740\ : Span4Mux_v
    port map (
            O => \N__11309\,
            I => \N__11222\
        );

    \I__2739\ : InMux
    port map (
            O => \N__11308\,
            I => \N__11217\
        );

    \I__2738\ : InMux
    port map (
            O => \N__11305\,
            I => \N__11217\
        );

    \I__2737\ : Span12Mux_v
    port map (
            O => \N__11298\,
            I => \N__11213\
        );

    \I__2736\ : Span12Mux_h
    port map (
            O => \N__11289\,
            I => \N__11210\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__11280\,
            I => \N__11201\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__11275\,
            I => \N__11201\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__11264\,
            I => \N__11201\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__11257\,
            I => \N__11201\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__11254\,
            I => \N__11198\
        );

    \I__2730\ : Span4Mux_v
    port map (
            O => \N__11249\,
            I => \N__11195\
        );

    \I__2729\ : InMux
    port map (
            O => \N__11246\,
            I => \N__11192\
        );

    \I__2728\ : Span4Mux_v
    port map (
            O => \N__11241\,
            I => \N__11187\
        );

    \I__2727\ : Span4Mux_v
    port map (
            O => \N__11234\,
            I => \N__11187\
        );

    \I__2726\ : InMux
    port map (
            O => \N__11233\,
            I => \N__11180\
        );

    \I__2725\ : InMux
    port map (
            O => \N__11232\,
            I => \N__11180\
        );

    \I__2724\ : InMux
    port map (
            O => \N__11231\,
            I => \N__11180\
        );

    \I__2723\ : Span4Mux_h
    port map (
            O => \N__11228\,
            I => \N__11177\
        );

    \I__2722\ : Sp12to4
    port map (
            O => \N__11225\,
            I => \N__11172\
        );

    \I__2721\ : Sp12to4
    port map (
            O => \N__11222\,
            I => \N__11172\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__11217\,
            I => \N__11169\
        );

    \I__2719\ : InMux
    port map (
            O => \N__11216\,
            I => \N__11166\
        );

    \I__2718\ : Span12Mux_h
    port map (
            O => \N__11213\,
            I => \N__11161\
        );

    \I__2717\ : Span12Mux_v
    port map (
            O => \N__11210\,
            I => \N__11161\
        );

    \I__2716\ : Span12Mux_v
    port map (
            O => \N__11201\,
            I => \N__11152\
        );

    \I__2715\ : Span12Mux_s8_v
    port map (
            O => \N__11198\,
            I => \N__11152\
        );

    \I__2714\ : Sp12to4
    port map (
            O => \N__11195\,
            I => \N__11152\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__11192\,
            I => \N__11152\
        );

    \I__2712\ : Sp12to4
    port map (
            O => \N__11187\,
            I => \N__11147\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__11180\,
            I => \N__11147\
        );

    \I__2710\ : Sp12to4
    port map (
            O => \N__11177\,
            I => \N__11140\
        );

    \I__2709\ : Span12Mux_h
    port map (
            O => \N__11172\,
            I => \N__11140\
        );

    \I__2708\ : Sp12to4
    port map (
            O => \N__11169\,
            I => \N__11140\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__11166\,
            I => \N__11137\
        );

    \I__2706\ : Span12Mux_v
    port map (
            O => \N__11161\,
            I => \N__11134\
        );

    \I__2705\ : Span12Mux_h
    port map (
            O => \N__11152\,
            I => \N__11127\
        );

    \I__2704\ : Span12Mux_h
    port map (
            O => \N__11147\,
            I => \N__11127\
        );

    \I__2703\ : Span12Mux_v
    port map (
            O => \N__11140\,
            I => \N__11127\
        );

    \I__2702\ : Span4Mux_v
    port map (
            O => \N__11137\,
            I => \N__11124\
        );

    \I__2701\ : Odrv12
    port map (
            O => \N__11134\,
            I => \LBENn_c\
        );

    \I__2700\ : Odrv12
    port map (
            O => \N__11127\,
            I => \LBENn_c\
        );

    \I__2699\ : Odrv4
    port map (
            O => \N__11124\,
            I => \LBENn_c\
        );

    \I__2698\ : InMux
    port map (
            O => \N__11117\,
            I => \N__11103\
        );

    \I__2697\ : InMux
    port map (
            O => \N__11116\,
            I => \N__11100\
        );

    \I__2696\ : InMux
    port map (
            O => \N__11115\,
            I => \N__11097\
        );

    \I__2695\ : InMux
    port map (
            O => \N__11114\,
            I => \N__11094\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__11113\,
            I => \N__11080\
        );

    \I__2693\ : InMux
    port map (
            O => \N__11112\,
            I => \N__11076\
        );

    \I__2692\ : InMux
    port map (
            O => \N__11111\,
            I => \N__11071\
        );

    \I__2691\ : InMux
    port map (
            O => \N__11110\,
            I => \N__11071\
        );

    \I__2690\ : InMux
    port map (
            O => \N__11109\,
            I => \N__11066\
        );

    \I__2689\ : InMux
    port map (
            O => \N__11108\,
            I => \N__11066\
        );

    \I__2688\ : CascadeMux
    port map (
            O => \N__11107\,
            I => \N__11061\
        );

    \I__2687\ : CascadeMux
    port map (
            O => \N__11106\,
            I => \N__11058\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__11103\,
            I => \N__11054\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__11100\,
            I => \N__11049\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__11097\,
            I => \N__11049\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__11094\,
            I => \N__11046\
        );

    \I__2682\ : InMux
    port map (
            O => \N__11093\,
            I => \N__11043\
        );

    \I__2681\ : InMux
    port map (
            O => \N__11092\,
            I => \N__11040\
        );

    \I__2680\ : InMux
    port map (
            O => \N__11091\,
            I => \N__11037\
        );

    \I__2679\ : InMux
    port map (
            O => \N__11090\,
            I => \N__11034\
        );

    \I__2678\ : InMux
    port map (
            O => \N__11089\,
            I => \N__11022\
        );

    \I__2677\ : InMux
    port map (
            O => \N__11088\,
            I => \N__11022\
        );

    \I__2676\ : InMux
    port map (
            O => \N__11087\,
            I => \N__11022\
        );

    \I__2675\ : InMux
    port map (
            O => \N__11086\,
            I => \N__11017\
        );

    \I__2674\ : InMux
    port map (
            O => \N__11085\,
            I => \N__11017\
        );

    \I__2673\ : InMux
    port map (
            O => \N__11084\,
            I => \N__11008\
        );

    \I__2672\ : InMux
    port map (
            O => \N__11083\,
            I => \N__11008\
        );

    \I__2671\ : InMux
    port map (
            O => \N__11080\,
            I => \N__11003\
        );

    \I__2670\ : InMux
    port map (
            O => \N__11079\,
            I => \N__11003\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__11076\,
            I => \N__10996\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__11071\,
            I => \N__10996\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__11066\,
            I => \N__10993\
        );

    \I__2666\ : InMux
    port map (
            O => \N__11065\,
            I => \N__10990\
        );

    \I__2665\ : InMux
    port map (
            O => \N__11064\,
            I => \N__10987\
        );

    \I__2664\ : InMux
    port map (
            O => \N__11061\,
            I => \N__10980\
        );

    \I__2663\ : InMux
    port map (
            O => \N__11058\,
            I => \N__10980\
        );

    \I__2662\ : InMux
    port map (
            O => \N__11057\,
            I => \N__10980\
        );

    \I__2661\ : Span4Mux_v
    port map (
            O => \N__11054\,
            I => \N__10967\
        );

    \I__2660\ : Span4Mux_v
    port map (
            O => \N__11049\,
            I => \N__10967\
        );

    \I__2659\ : Span4Mux_h
    port map (
            O => \N__11046\,
            I => \N__10967\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__11043\,
            I => \N__10967\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__11040\,
            I => \N__10967\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__11037\,
            I => \N__10967\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__11034\,
            I => \N__10964\
        );

    \I__2654\ : InMux
    port map (
            O => \N__11033\,
            I => \N__10961\
        );

    \I__2653\ : InMux
    port map (
            O => \N__11032\,
            I => \N__10958\
        );

    \I__2652\ : InMux
    port map (
            O => \N__11031\,
            I => \N__10955\
        );

    \I__2651\ : InMux
    port map (
            O => \N__11030\,
            I => \N__10952\
        );

    \I__2650\ : InMux
    port map (
            O => \N__11029\,
            I => \N__10949\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__11022\,
            I => \N__10944\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__11017\,
            I => \N__10944\
        );

    \I__2647\ : InMux
    port map (
            O => \N__11016\,
            I => \N__10941\
        );

    \I__2646\ : InMux
    port map (
            O => \N__11015\,
            I => \N__10938\
        );

    \I__2645\ : InMux
    port map (
            O => \N__11014\,
            I => \N__10935\
        );

    \I__2644\ : InMux
    port map (
            O => \N__11013\,
            I => \N__10932\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__11008\,
            I => \N__10922\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__11003\,
            I => \N__10919\
        );

    \I__2641\ : InMux
    port map (
            O => \N__11002\,
            I => \N__10914\
        );

    \I__2640\ : InMux
    port map (
            O => \N__11001\,
            I => \N__10914\
        );

    \I__2639\ : Span4Mux_v
    port map (
            O => \N__10996\,
            I => \N__10903\
        );

    \I__2638\ : Span4Mux_h
    port map (
            O => \N__10993\,
            I => \N__10903\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__10990\,
            I => \N__10903\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__10987\,
            I => \N__10903\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__10980\,
            I => \N__10903\
        );

    \I__2634\ : Span4Mux_v
    port map (
            O => \N__10967\,
            I => \N__10888\
        );

    \I__2633\ : Span4Mux_h
    port map (
            O => \N__10964\,
            I => \N__10888\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__10961\,
            I => \N__10888\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__10958\,
            I => \N__10888\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__10955\,
            I => \N__10888\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__10952\,
            I => \N__10888\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__10949\,
            I => \N__10888\
        );

    \I__2627\ : Span4Mux_v
    port map (
            O => \N__10944\,
            I => \N__10883\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__10941\,
            I => \N__10883\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__10938\,
            I => \N__10880\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__10935\,
            I => \N__10877\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__10932\,
            I => \N__10874\
        );

    \I__2622\ : InMux
    port map (
            O => \N__10931\,
            I => \N__10871\
        );

    \I__2621\ : InMux
    port map (
            O => \N__10930\,
            I => \N__10868\
        );

    \I__2620\ : InMux
    port map (
            O => \N__10929\,
            I => \N__10860\
        );

    \I__2619\ : InMux
    port map (
            O => \N__10928\,
            I => \N__10853\
        );

    \I__2618\ : InMux
    port map (
            O => \N__10927\,
            I => \N__10853\
        );

    \I__2617\ : InMux
    port map (
            O => \N__10926\,
            I => \N__10853\
        );

    \I__2616\ : InMux
    port map (
            O => \N__10925\,
            I => \N__10850\
        );

    \I__2615\ : Span4Mux_h
    port map (
            O => \N__10922\,
            I => \N__10842\
        );

    \I__2614\ : Span12Mux_v
    port map (
            O => \N__10919\,
            I => \N__10837\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__10914\,
            I => \N__10834\
        );

    \I__2612\ : Span4Mux_v
    port map (
            O => \N__10903\,
            I => \N__10829\
        );

    \I__2611\ : Span4Mux_v
    port map (
            O => \N__10888\,
            I => \N__10829\
        );

    \I__2610\ : Span4Mux_h
    port map (
            O => \N__10883\,
            I => \N__10824\
        );

    \I__2609\ : Span4Mux_v
    port map (
            O => \N__10880\,
            I => \N__10824\
        );

    \I__2608\ : Span4Mux_v
    port map (
            O => \N__10877\,
            I => \N__10818\
        );

    \I__2607\ : Span4Mux_v
    port map (
            O => \N__10874\,
            I => \N__10815\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__10871\,
            I => \N__10812\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__10868\,
            I => \N__10809\
        );

    \I__2604\ : InMux
    port map (
            O => \N__10867\,
            I => \N__10806\
        );

    \I__2603\ : InMux
    port map (
            O => \N__10866\,
            I => \N__10803\
        );

    \I__2602\ : InMux
    port map (
            O => \N__10865\,
            I => \N__10796\
        );

    \I__2601\ : InMux
    port map (
            O => \N__10864\,
            I => \N__10796\
        );

    \I__2600\ : InMux
    port map (
            O => \N__10863\,
            I => \N__10796\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__10860\,
            I => \N__10788\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__10853\,
            I => \N__10788\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__10850\,
            I => \N__10785\
        );

    \I__2596\ : InMux
    port map (
            O => \N__10849\,
            I => \N__10774\
        );

    \I__2595\ : InMux
    port map (
            O => \N__10848\,
            I => \N__10774\
        );

    \I__2594\ : InMux
    port map (
            O => \N__10847\,
            I => \N__10774\
        );

    \I__2593\ : InMux
    port map (
            O => \N__10846\,
            I => \N__10774\
        );

    \I__2592\ : InMux
    port map (
            O => \N__10845\,
            I => \N__10774\
        );

    \I__2591\ : Span4Mux_h
    port map (
            O => \N__10842\,
            I => \N__10771\
        );

    \I__2590\ : InMux
    port map (
            O => \N__10841\,
            I => \N__10766\
        );

    \I__2589\ : InMux
    port map (
            O => \N__10840\,
            I => \N__10766\
        );

    \I__2588\ : Span12Mux_h
    port map (
            O => \N__10837\,
            I => \N__10759\
        );

    \I__2587\ : Span4Mux_h
    port map (
            O => \N__10834\,
            I => \N__10756\
        );

    \I__2586\ : Sp12to4
    port map (
            O => \N__10829\,
            I => \N__10753\
        );

    \I__2585\ : Span4Mux_v
    port map (
            O => \N__10824\,
            I => \N__10750\
        );

    \I__2584\ : InMux
    port map (
            O => \N__10823\,
            I => \N__10747\
        );

    \I__2583\ : InMux
    port map (
            O => \N__10822\,
            I => \N__10742\
        );

    \I__2582\ : InMux
    port map (
            O => \N__10821\,
            I => \N__10742\
        );

    \I__2581\ : Span4Mux_v
    port map (
            O => \N__10818\,
            I => \N__10739\
        );

    \I__2580\ : Span4Mux_h
    port map (
            O => \N__10815\,
            I => \N__10734\
        );

    \I__2579\ : Span4Mux_v
    port map (
            O => \N__10812\,
            I => \N__10734\
        );

    \I__2578\ : Span4Mux_v
    port map (
            O => \N__10809\,
            I => \N__10727\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__10806\,
            I => \N__10727\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__10803\,
            I => \N__10727\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__10796\,
            I => \N__10724\
        );

    \I__2574\ : InMux
    port map (
            O => \N__10795\,
            I => \N__10717\
        );

    \I__2573\ : InMux
    port map (
            O => \N__10794\,
            I => \N__10717\
        );

    \I__2572\ : InMux
    port map (
            O => \N__10793\,
            I => \N__10717\
        );

    \I__2571\ : Span4Mux_v
    port map (
            O => \N__10788\,
            I => \N__10710\
        );

    \I__2570\ : Span4Mux_h
    port map (
            O => \N__10785\,
            I => \N__10710\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__10774\,
            I => \N__10710\
        );

    \I__2568\ : Span4Mux_h
    port map (
            O => \N__10771\,
            I => \N__10705\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__10766\,
            I => \N__10705\
        );

    \I__2566\ : InMux
    port map (
            O => \N__10765\,
            I => \N__10696\
        );

    \I__2565\ : InMux
    port map (
            O => \N__10764\,
            I => \N__10696\
        );

    \I__2564\ : InMux
    port map (
            O => \N__10763\,
            I => \N__10696\
        );

    \I__2563\ : InMux
    port map (
            O => \N__10762\,
            I => \N__10696\
        );

    \I__2562\ : Span12Mux_h
    port map (
            O => \N__10759\,
            I => \N__10693\
        );

    \I__2561\ : Sp12to4
    port map (
            O => \N__10756\,
            I => \N__10690\
        );

    \I__2560\ : Span12Mux_h
    port map (
            O => \N__10753\,
            I => \N__10683\
        );

    \I__2559\ : Sp12to4
    port map (
            O => \N__10750\,
            I => \N__10683\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__10747\,
            I => \N__10683\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__10742\,
            I => \N__10680\
        );

    \I__2556\ : Span4Mux_v
    port map (
            O => \N__10739\,
            I => \N__10677\
        );

    \I__2555\ : Span4Mux_h
    port map (
            O => \N__10734\,
            I => \N__10674\
        );

    \I__2554\ : Span4Mux_h
    port map (
            O => \N__10727\,
            I => \N__10667\
        );

    \I__2553\ : Span4Mux_v
    port map (
            O => \N__10724\,
            I => \N__10667\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__10717\,
            I => \N__10667\
        );

    \I__2551\ : Span4Mux_v
    port map (
            O => \N__10710\,
            I => \N__10660\
        );

    \I__2550\ : Span4Mux_h
    port map (
            O => \N__10705\,
            I => \N__10660\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__10696\,
            I => \N__10660\
        );

    \I__2548\ : Span12Mux_v
    port map (
            O => \N__10693\,
            I => \N__10657\
        );

    \I__2547\ : Span12Mux_v
    port map (
            O => \N__10690\,
            I => \N__10650\
        );

    \I__2546\ : Span12Mux_h
    port map (
            O => \N__10683\,
            I => \N__10650\
        );

    \I__2545\ : Span12Mux_v
    port map (
            O => \N__10680\,
            I => \N__10650\
        );

    \I__2544\ : Span4Mux_h
    port map (
            O => \N__10677\,
            I => \N__10645\
        );

    \I__2543\ : Span4Mux_v
    port map (
            O => \N__10674\,
            I => \N__10645\
        );

    \I__2542\ : Span4Mux_v
    port map (
            O => \N__10667\,
            I => \N__10640\
        );

    \I__2541\ : Span4Mux_v
    port map (
            O => \N__10660\,
            I => \N__10640\
        );

    \I__2540\ : Odrv12
    port map (
            O => \N__10657\,
            I => \BGn_c\
        );

    \I__2539\ : Odrv12
    port map (
            O => \N__10650\,
            I => \BGn_c\
        );

    \I__2538\ : Odrv4
    port map (
            O => \N__10645\,
            I => \BGn_c\
        );

    \I__2537\ : Odrv4
    port map (
            O => \N__10640\,
            I => \BGn_c\
        );

    \I__2536\ : InMux
    port map (
            O => \N__10631\,
            I => \N__10628\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__10628\,
            I => \N__10611\
        );

    \I__2534\ : ClkMux
    port map (
            O => \N__10627\,
            I => \N__10448\
        );

    \I__2533\ : ClkMux
    port map (
            O => \N__10626\,
            I => \N__10448\
        );

    \I__2532\ : ClkMux
    port map (
            O => \N__10625\,
            I => \N__10448\
        );

    \I__2531\ : ClkMux
    port map (
            O => \N__10624\,
            I => \N__10448\
        );

    \I__2530\ : ClkMux
    port map (
            O => \N__10623\,
            I => \N__10448\
        );

    \I__2529\ : ClkMux
    port map (
            O => \N__10622\,
            I => \N__10448\
        );

    \I__2528\ : ClkMux
    port map (
            O => \N__10621\,
            I => \N__10448\
        );

    \I__2527\ : ClkMux
    port map (
            O => \N__10620\,
            I => \N__10448\
        );

    \I__2526\ : ClkMux
    port map (
            O => \N__10619\,
            I => \N__10448\
        );

    \I__2525\ : ClkMux
    port map (
            O => \N__10618\,
            I => \N__10448\
        );

    \I__2524\ : ClkMux
    port map (
            O => \N__10617\,
            I => \N__10448\
        );

    \I__2523\ : ClkMux
    port map (
            O => \N__10616\,
            I => \N__10448\
        );

    \I__2522\ : ClkMux
    port map (
            O => \N__10615\,
            I => \N__10448\
        );

    \I__2521\ : ClkMux
    port map (
            O => \N__10614\,
            I => \N__10448\
        );

    \I__2520\ : Glb2LocalMux
    port map (
            O => \N__10611\,
            I => \N__10448\
        );

    \I__2519\ : ClkMux
    port map (
            O => \N__10610\,
            I => \N__10448\
        );

    \I__2518\ : ClkMux
    port map (
            O => \N__10609\,
            I => \N__10448\
        );

    \I__2517\ : ClkMux
    port map (
            O => \N__10608\,
            I => \N__10448\
        );

    \I__2516\ : ClkMux
    port map (
            O => \N__10607\,
            I => \N__10448\
        );

    \I__2515\ : ClkMux
    port map (
            O => \N__10606\,
            I => \N__10448\
        );

    \I__2514\ : ClkMux
    port map (
            O => \N__10605\,
            I => \N__10448\
        );

    \I__2513\ : ClkMux
    port map (
            O => \N__10604\,
            I => \N__10448\
        );

    \I__2512\ : ClkMux
    port map (
            O => \N__10603\,
            I => \N__10448\
        );

    \I__2511\ : ClkMux
    port map (
            O => \N__10602\,
            I => \N__10448\
        );

    \I__2510\ : ClkMux
    port map (
            O => \N__10601\,
            I => \N__10448\
        );

    \I__2509\ : ClkMux
    port map (
            O => \N__10600\,
            I => \N__10448\
        );

    \I__2508\ : ClkMux
    port map (
            O => \N__10599\,
            I => \N__10448\
        );

    \I__2507\ : ClkMux
    port map (
            O => \N__10598\,
            I => \N__10448\
        );

    \I__2506\ : ClkMux
    port map (
            O => \N__10597\,
            I => \N__10448\
        );

    \I__2505\ : ClkMux
    port map (
            O => \N__10596\,
            I => \N__10448\
        );

    \I__2504\ : ClkMux
    port map (
            O => \N__10595\,
            I => \N__10448\
        );

    \I__2503\ : ClkMux
    port map (
            O => \N__10594\,
            I => \N__10448\
        );

    \I__2502\ : ClkMux
    port map (
            O => \N__10593\,
            I => \N__10448\
        );

    \I__2501\ : ClkMux
    port map (
            O => \N__10592\,
            I => \N__10448\
        );

    \I__2500\ : ClkMux
    port map (
            O => \N__10591\,
            I => \N__10448\
        );

    \I__2499\ : ClkMux
    port map (
            O => \N__10590\,
            I => \N__10448\
        );

    \I__2498\ : ClkMux
    port map (
            O => \N__10589\,
            I => \N__10448\
        );

    \I__2497\ : ClkMux
    port map (
            O => \N__10588\,
            I => \N__10448\
        );

    \I__2496\ : ClkMux
    port map (
            O => \N__10587\,
            I => \N__10448\
        );

    \I__2495\ : ClkMux
    port map (
            O => \N__10586\,
            I => \N__10448\
        );

    \I__2494\ : ClkMux
    port map (
            O => \N__10585\,
            I => \N__10448\
        );

    \I__2493\ : ClkMux
    port map (
            O => \N__10584\,
            I => \N__10448\
        );

    \I__2492\ : ClkMux
    port map (
            O => \N__10583\,
            I => \N__10448\
        );

    \I__2491\ : ClkMux
    port map (
            O => \N__10582\,
            I => \N__10448\
        );

    \I__2490\ : ClkMux
    port map (
            O => \N__10581\,
            I => \N__10448\
        );

    \I__2489\ : ClkMux
    port map (
            O => \N__10580\,
            I => \N__10448\
        );

    \I__2488\ : ClkMux
    port map (
            O => \N__10579\,
            I => \N__10448\
        );

    \I__2487\ : ClkMux
    port map (
            O => \N__10578\,
            I => \N__10448\
        );

    \I__2486\ : ClkMux
    port map (
            O => \N__10577\,
            I => \N__10448\
        );

    \I__2485\ : ClkMux
    port map (
            O => \N__10576\,
            I => \N__10448\
        );

    \I__2484\ : ClkMux
    port map (
            O => \N__10575\,
            I => \N__10448\
        );

    \I__2483\ : ClkMux
    port map (
            O => \N__10574\,
            I => \N__10448\
        );

    \I__2482\ : ClkMux
    port map (
            O => \N__10573\,
            I => \N__10448\
        );

    \I__2481\ : ClkMux
    port map (
            O => \N__10572\,
            I => \N__10448\
        );

    \I__2480\ : ClkMux
    port map (
            O => \N__10571\,
            I => \N__10448\
        );

    \I__2479\ : ClkMux
    port map (
            O => \N__10570\,
            I => \N__10448\
        );

    \I__2478\ : ClkMux
    port map (
            O => \N__10569\,
            I => \N__10448\
        );

    \I__2477\ : ClkMux
    port map (
            O => \N__10568\,
            I => \N__10448\
        );

    \I__2476\ : ClkMux
    port map (
            O => \N__10567\,
            I => \N__10448\
        );

    \I__2475\ : GlobalMux
    port map (
            O => \N__10448\,
            I => \CLK40\
        );

    \I__2474\ : CEMux
    port map (
            O => \N__10445\,
            I => \N__10325\
        );

    \I__2473\ : CEMux
    port map (
            O => \N__10444\,
            I => \N__10325\
        );

    \I__2472\ : CEMux
    port map (
            O => \N__10443\,
            I => \N__10325\
        );

    \I__2471\ : CEMux
    port map (
            O => \N__10442\,
            I => \N__10325\
        );

    \I__2470\ : CEMux
    port map (
            O => \N__10441\,
            I => \N__10325\
        );

    \I__2469\ : CEMux
    port map (
            O => \N__10440\,
            I => \N__10325\
        );

    \I__2468\ : CEMux
    port map (
            O => \N__10439\,
            I => \N__10325\
        );

    \I__2467\ : CEMux
    port map (
            O => \N__10438\,
            I => \N__10325\
        );

    \I__2466\ : CEMux
    port map (
            O => \N__10437\,
            I => \N__10325\
        );

    \I__2465\ : CEMux
    port map (
            O => \N__10436\,
            I => \N__10325\
        );

    \I__2464\ : CEMux
    port map (
            O => \N__10435\,
            I => \N__10325\
        );

    \I__2463\ : CEMux
    port map (
            O => \N__10434\,
            I => \N__10325\
        );

    \I__2462\ : CEMux
    port map (
            O => \N__10433\,
            I => \N__10325\
        );

    \I__2461\ : CEMux
    port map (
            O => \N__10432\,
            I => \N__10325\
        );

    \I__2460\ : CEMux
    port map (
            O => \N__10431\,
            I => \N__10325\
        );

    \I__2459\ : CEMux
    port map (
            O => \N__10430\,
            I => \N__10325\
        );

    \I__2458\ : CEMux
    port map (
            O => \N__10429\,
            I => \N__10325\
        );

    \I__2457\ : CEMux
    port map (
            O => \N__10428\,
            I => \N__10325\
        );

    \I__2456\ : CEMux
    port map (
            O => \N__10427\,
            I => \N__10325\
        );

    \I__2455\ : CEMux
    port map (
            O => \N__10426\,
            I => \N__10325\
        );

    \I__2454\ : CEMux
    port map (
            O => \N__10425\,
            I => \N__10325\
        );

    \I__2453\ : CEMux
    port map (
            O => \N__10424\,
            I => \N__10325\
        );

    \I__2452\ : CEMux
    port map (
            O => \N__10423\,
            I => \N__10325\
        );

    \I__2451\ : CEMux
    port map (
            O => \N__10422\,
            I => \N__10325\
        );

    \I__2450\ : CEMux
    port map (
            O => \N__10421\,
            I => \N__10325\
        );

    \I__2449\ : CEMux
    port map (
            O => \N__10420\,
            I => \N__10325\
        );

    \I__2448\ : CEMux
    port map (
            O => \N__10419\,
            I => \N__10325\
        );

    \I__2447\ : CEMux
    port map (
            O => \N__10418\,
            I => \N__10325\
        );

    \I__2446\ : CEMux
    port map (
            O => \N__10417\,
            I => \N__10325\
        );

    \I__2445\ : CEMux
    port map (
            O => \N__10416\,
            I => \N__10325\
        );

    \I__2444\ : CEMux
    port map (
            O => \N__10415\,
            I => \N__10325\
        );

    \I__2443\ : CEMux
    port map (
            O => \N__10414\,
            I => \N__10325\
        );

    \I__2442\ : CEMux
    port map (
            O => \N__10413\,
            I => \N__10325\
        );

    \I__2441\ : CEMux
    port map (
            O => \N__10412\,
            I => \N__10325\
        );

    \I__2440\ : CEMux
    port map (
            O => \N__10411\,
            I => \N__10325\
        );

    \I__2439\ : CEMux
    port map (
            O => \N__10410\,
            I => \N__10325\
        );

    \I__2438\ : CEMux
    port map (
            O => \N__10409\,
            I => \N__10325\
        );

    \I__2437\ : CEMux
    port map (
            O => \N__10408\,
            I => \N__10325\
        );

    \I__2436\ : CEMux
    port map (
            O => \N__10407\,
            I => \N__10325\
        );

    \I__2435\ : CEMux
    port map (
            O => \N__10406\,
            I => \N__10325\
        );

    \I__2434\ : GlobalMux
    port map (
            O => \N__10325\,
            I => \N__10322\
        );

    \I__2433\ : gio2CtrlBuf
    port map (
            O => \N__10322\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_g_0\
        );

    \I__2432\ : InMux
    port map (
            O => \N__10319\,
            I => \N__10316\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__10316\,
            I => \N__10266\
        );

    \I__2430\ : SRMux
    port map (
            O => \N__10315\,
            I => \N__10169\
        );

    \I__2429\ : SRMux
    port map (
            O => \N__10314\,
            I => \N__10169\
        );

    \I__2428\ : SRMux
    port map (
            O => \N__10313\,
            I => \N__10169\
        );

    \I__2427\ : SRMux
    port map (
            O => \N__10312\,
            I => \N__10169\
        );

    \I__2426\ : SRMux
    port map (
            O => \N__10311\,
            I => \N__10169\
        );

    \I__2425\ : SRMux
    port map (
            O => \N__10310\,
            I => \N__10169\
        );

    \I__2424\ : SRMux
    port map (
            O => \N__10309\,
            I => \N__10169\
        );

    \I__2423\ : SRMux
    port map (
            O => \N__10308\,
            I => \N__10169\
        );

    \I__2422\ : SRMux
    port map (
            O => \N__10307\,
            I => \N__10169\
        );

    \I__2421\ : SRMux
    port map (
            O => \N__10306\,
            I => \N__10169\
        );

    \I__2420\ : SRMux
    port map (
            O => \N__10305\,
            I => \N__10169\
        );

    \I__2419\ : SRMux
    port map (
            O => \N__10304\,
            I => \N__10169\
        );

    \I__2418\ : SRMux
    port map (
            O => \N__10303\,
            I => \N__10169\
        );

    \I__2417\ : SRMux
    port map (
            O => \N__10302\,
            I => \N__10169\
        );

    \I__2416\ : SRMux
    port map (
            O => \N__10301\,
            I => \N__10169\
        );

    \I__2415\ : SRMux
    port map (
            O => \N__10300\,
            I => \N__10169\
        );

    \I__2414\ : SRMux
    port map (
            O => \N__10299\,
            I => \N__10169\
        );

    \I__2413\ : SRMux
    port map (
            O => \N__10298\,
            I => \N__10169\
        );

    \I__2412\ : SRMux
    port map (
            O => \N__10297\,
            I => \N__10169\
        );

    \I__2411\ : SRMux
    port map (
            O => \N__10296\,
            I => \N__10169\
        );

    \I__2410\ : SRMux
    port map (
            O => \N__10295\,
            I => \N__10169\
        );

    \I__2409\ : SRMux
    port map (
            O => \N__10294\,
            I => \N__10169\
        );

    \I__2408\ : SRMux
    port map (
            O => \N__10293\,
            I => \N__10169\
        );

    \I__2407\ : SRMux
    port map (
            O => \N__10292\,
            I => \N__10169\
        );

    \I__2406\ : SRMux
    port map (
            O => \N__10291\,
            I => \N__10169\
        );

    \I__2405\ : SRMux
    port map (
            O => \N__10290\,
            I => \N__10169\
        );

    \I__2404\ : SRMux
    port map (
            O => \N__10289\,
            I => \N__10169\
        );

    \I__2403\ : SRMux
    port map (
            O => \N__10288\,
            I => \N__10169\
        );

    \I__2402\ : SRMux
    port map (
            O => \N__10287\,
            I => \N__10169\
        );

    \I__2401\ : SRMux
    port map (
            O => \N__10286\,
            I => \N__10169\
        );

    \I__2400\ : SRMux
    port map (
            O => \N__10285\,
            I => \N__10169\
        );

    \I__2399\ : SRMux
    port map (
            O => \N__10284\,
            I => \N__10169\
        );

    \I__2398\ : SRMux
    port map (
            O => \N__10283\,
            I => \N__10169\
        );

    \I__2397\ : SRMux
    port map (
            O => \N__10282\,
            I => \N__10169\
        );

    \I__2396\ : SRMux
    port map (
            O => \N__10281\,
            I => \N__10169\
        );

    \I__2395\ : SRMux
    port map (
            O => \N__10280\,
            I => \N__10169\
        );

    \I__2394\ : SRMux
    port map (
            O => \N__10279\,
            I => \N__10169\
        );

    \I__2393\ : SRMux
    port map (
            O => \N__10278\,
            I => \N__10169\
        );

    \I__2392\ : SRMux
    port map (
            O => \N__10277\,
            I => \N__10169\
        );

    \I__2391\ : SRMux
    port map (
            O => \N__10276\,
            I => \N__10169\
        );

    \I__2390\ : SRMux
    port map (
            O => \N__10275\,
            I => \N__10169\
        );

    \I__2389\ : SRMux
    port map (
            O => \N__10274\,
            I => \N__10169\
        );

    \I__2388\ : SRMux
    port map (
            O => \N__10273\,
            I => \N__10169\
        );

    \I__2387\ : SRMux
    port map (
            O => \N__10272\,
            I => \N__10169\
        );

    \I__2386\ : SRMux
    port map (
            O => \N__10271\,
            I => \N__10169\
        );

    \I__2385\ : SRMux
    port map (
            O => \N__10270\,
            I => \N__10169\
        );

    \I__2384\ : SRMux
    port map (
            O => \N__10269\,
            I => \N__10169\
        );

    \I__2383\ : Glb2LocalMux
    port map (
            O => \N__10266\,
            I => \N__10169\
        );

    \I__2382\ : GlobalMux
    port map (
            O => \N__10169\,
            I => \N__10166\
        );

    \I__2381\ : gio2CtrlBuf
    port map (
            O => \N__10166\,
            I => \RESETn_c_i_g\
        );

    \I__2380\ : InMux
    port map (
            O => \N__10163\,
            I => \N__10160\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__10160\,
            I => \READ_CYCLE_ACTIVE_rep1_i_ess\
        );

    \I__2378\ : IoInMux
    port map (
            O => \N__10157\,
            I => \N__10154\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__10154\,
            I => \N__10151\
        );

    \I__2376\ : IoSpan4Mux
    port map (
            O => \N__10151\,
            I => \N__10148\
        );

    \I__2375\ : Span4Mux_s3_h
    port map (
            O => \N__10148\,
            I => \N__10145\
        );

    \I__2374\ : Odrv4
    port map (
            O => \N__10145\,
            I => \N_181_i\
        );

    \I__2373\ : InMux
    port map (
            O => \N__10142\,
            I => \N__10139\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__10139\,
            I => \READ_CYCLE_ACTIVE_rep12_i_ess\
        );

    \I__2371\ : IoInMux
    port map (
            O => \N__10136\,
            I => \N__10133\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__10133\,
            I => \N__10130\
        );

    \I__2369\ : Span4Mux_s2_v
    port map (
            O => \N__10130\,
            I => \N__10127\
        );

    \I__2368\ : Span4Mux_v
    port map (
            O => \N__10127\,
            I => \N__10124\
        );

    \I__2367\ : Odrv4
    port map (
            O => \N__10124\,
            I => \N_192_i\
        );

    \I__2366\ : InMux
    port map (
            O => \N__10121\,
            I => \N__10118\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__10118\,
            I => \READ_CYCLE_ACTIVE_rep14_i_ess\
        );

    \I__2364\ : InMux
    port map (
            O => \N__10115\,
            I => \N__10112\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__10112\,
            I => \READ_CYCLE_ACTIVE_rep10_i_ess\
        );

    \I__2362\ : InMux
    port map (
            O => \N__10109\,
            I => \N__10106\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__10106\,
            I => \READ_CYCLE_ACTIVE_rep22_i_ess\
        );

    \I__2360\ : IoInMux
    port map (
            O => \N__10103\,
            I => \N__10100\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__10100\,
            I => \N__10097\
        );

    \I__2358\ : Span4Mux_s3_h
    port map (
            O => \N__10097\,
            I => \N__10094\
        );

    \I__2357\ : Odrv4
    port map (
            O => \N__10094\,
            I => \N_202_i\
        );

    \I__2356\ : InMux
    port map (
            O => \N__10091\,
            I => \N__10088\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__10088\,
            I => \N__10085\
        );

    \I__2354\ : Odrv4
    port map (
            O => \N__10085\,
            I => \READ_CYCLE_ACTIVE_rep23_i_ess\
        );

    \I__2353\ : IoInMux
    port map (
            O => \N__10082\,
            I => \N__10079\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__10079\,
            I => \N__10076\
        );

    \I__2351\ : Span4Mux_s3_h
    port map (
            O => \N__10076\,
            I => \N__10073\
        );

    \I__2350\ : Odrv4
    port map (
            O => \N__10073\,
            I => \N_203_i\
        );

    \I__2349\ : InMux
    port map (
            O => \N__10070\,
            I => \N__10067\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__10067\,
            I => \READ_CYCLE_ACTIVE_rep18_i_ess\
        );

    \I__2347\ : InMux
    port map (
            O => \N__10064\,
            I => \N__10061\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__10061\,
            I => \N__10058\
        );

    \I__2345\ : Odrv4
    port map (
            O => \N__10058\,
            I => \READ_CYCLE_ACTIVE_rep17_i_ess\
        );

    \I__2344\ : IoInMux
    port map (
            O => \N__10055\,
            I => \N__10052\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__10052\,
            I => \N__10049\
        );

    \I__2342\ : IoSpan4Mux
    port map (
            O => \N__10049\,
            I => \N__10046\
        );

    \I__2341\ : Span4Mux_s2_h
    port map (
            O => \N__10046\,
            I => \N__10043\
        );

    \I__2340\ : Odrv4
    port map (
            O => \N__10043\,
            I => \N_200_i\
        );

    \I__2339\ : IoInMux
    port map (
            O => \N__10040\,
            I => \N__10037\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__10037\,
            I => \N__10034\
        );

    \I__2337\ : Odrv12
    port map (
            O => \N__10034\,
            I => \N_188_i\
        );

    \I__2336\ : InMux
    port map (
            O => \N__10031\,
            I => \N__10028\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__10028\,
            I => \READ_CYCLE_ACTIVE_rep21_i_ess\
        );

    \I__2334\ : IoInMux
    port map (
            O => \N__10025\,
            I => \N__10022\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__10022\,
            I => \N__10019\
        );

    \I__2332\ : Odrv12
    port map (
            O => \N__10019\,
            I => \N_201_i\
        );

    \I__2331\ : InMux
    port map (
            O => \N__10016\,
            I => \N__10013\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__10013\,
            I => \READ_CYCLE_ACTIVE_rep20_i_ess\
        );

    \I__2329\ : InMux
    port map (
            O => \N__10010\,
            I => \N__10007\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__10007\,
            I => \READ_CYCLE_ACTIVE_rep8_i_ess\
        );

    \I__2327\ : IoInMux
    port map (
            O => \N__10004\,
            I => \N__10001\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__10001\,
            I => \N__9998\
        );

    \I__2325\ : Span4Mux_s3_h
    port map (
            O => \N__9998\,
            I => \N__9995\
        );

    \I__2324\ : Odrv4
    port map (
            O => \N__9995\,
            I => \N_190_i\
        );

    \I__2323\ : IoInMux
    port map (
            O => \N__9992\,
            I => \N__9989\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__9989\,
            I => \N__9986\
        );

    \I__2321\ : Span4Mux_s3_h
    port map (
            O => \N__9986\,
            I => \N__9983\
        );

    \I__2320\ : Odrv4
    port map (
            O => \N__9983\,
            I => \N_194_i\
        );

    \I__2319\ : InMux
    port map (
            O => \N__9980\,
            I => \N__9977\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__9977\,
            I => \READ_CYCLE_ACTIVE_rep29_i_ess\
        );

    \I__2317\ : InMux
    port map (
            O => \N__9974\,
            I => \N__9971\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__9971\,
            I => \READ_CYCLE_ACTIVE_rep24_i_ess\
        );

    \I__2315\ : InMux
    port map (
            O => \N__9968\,
            I => \N__9965\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__9965\,
            I => \READ_CYCLE_ACTIVE_rep26_i_ess\
        );

    \I__2313\ : IoInMux
    port map (
            O => \N__9962\,
            I => \N__9959\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__9959\,
            I => \N__9956\
        );

    \I__2311\ : Span4Mux_s3_h
    port map (
            O => \N__9956\,
            I => \N__9953\
        );

    \I__2310\ : Span4Mux_v
    port map (
            O => \N__9953\,
            I => \N__9950\
        );

    \I__2309\ : Odrv4
    port map (
            O => \N__9950\,
            I => \N_197_i\
        );

    \I__2308\ : IoInMux
    port map (
            O => \N__9947\,
            I => \N__9944\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__9944\,
            I => \N__9941\
        );

    \I__2306\ : IoSpan4Mux
    port map (
            O => \N__9941\,
            I => \N__9938\
        );

    \I__2305\ : Span4Mux_s0_h
    port map (
            O => \N__9938\,
            I => \N__9935\
        );

    \I__2304\ : Span4Mux_v
    port map (
            O => \N__9935\,
            I => \N__9932\
        );

    \I__2303\ : Odrv4
    port map (
            O => \N__9932\,
            I => \N_211_i\
        );

    \I__2302\ : IoInMux
    port map (
            O => \N__9929\,
            I => \N__9926\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__9926\,
            I => \N__9923\
        );

    \I__2300\ : Span4Mux_s3_h
    port map (
            O => \N__9923\,
            I => \N__9920\
        );

    \I__2299\ : Span4Mux_v
    port map (
            O => \N__9920\,
            I => \N__9917\
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__9917\,
            I => \N_198_i\
        );

    \I__2297\ : IoInMux
    port map (
            O => \N__9914\,
            I => \N__9911\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__9911\,
            I => \N__9908\
        );

    \I__2295\ : Span4Mux_s3_h
    port map (
            O => \N__9908\,
            I => \N__9905\
        );

    \I__2294\ : Odrv4
    port map (
            O => \N__9905\,
            I => \N_199_i\
        );

    \I__2293\ : InMux
    port map (
            O => \N__9902\,
            I => \N__9899\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__9899\,
            I => \N__9896\
        );

    \I__2291\ : Odrv4
    port map (
            O => \N__9896\,
            I => \READ_CYCLE_ACTIVE_rep31_i_ess\
        );

    \I__2290\ : InMux
    port map (
            O => \N__9893\,
            I => \N__9890\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__9890\,
            I => \READ_CYCLE_ACTIVE_rep19_i_ess\
        );

    \I__2288\ : InMux
    port map (
            O => \N__9887\,
            I => \N__9884\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__9884\,
            I => \N__9881\
        );

    \I__2286\ : Odrv12
    port map (
            O => \N__9881\,
            I => \READ_CYCLE_ACTIVE_rep5_i_ess\
        );

    \I__2285\ : IoInMux
    port map (
            O => \N__9878\,
            I => \N__9875\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__9875\,
            I => \N__9872\
        );

    \I__2283\ : Span4Mux_s2_v
    port map (
            O => \N__9872\,
            I => \N__9869\
        );

    \I__2282\ : Span4Mux_v
    port map (
            O => \N__9869\,
            I => \N__9866\
        );

    \I__2281\ : Odrv4
    port map (
            O => \N__9866\,
            I => \N_185_i\
        );

    \I__2280\ : InMux
    port map (
            O => \N__9863\,
            I => \N__9860\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__9860\,
            I => \READ_CYCLE_ACTIVE_rep13_i_ess\
        );

    \I__2278\ : IoInMux
    port map (
            O => \N__9857\,
            I => \N__9854\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__9854\,
            I => \N__9851\
        );

    \I__2276\ : Span4Mux_s2_v
    port map (
            O => \N__9851\,
            I => \N__9848\
        );

    \I__2275\ : Span4Mux_v
    port map (
            O => \N__9848\,
            I => \N__9845\
        );

    \I__2274\ : Odrv4
    port map (
            O => \N__9845\,
            I => \N_193_i\
        );

    \I__2273\ : IoInMux
    port map (
            O => \N__9842\,
            I => \N__9839\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__9839\,
            I => \N__9836\
        );

    \I__2271\ : Span4Mux_s3_h
    port map (
            O => \N__9836\,
            I => \N__9833\
        );

    \I__2270\ : Span4Mux_v
    port map (
            O => \N__9833\,
            I => \N__9830\
        );

    \I__2269\ : Odrv4
    port map (
            O => \N__9830\,
            I => \N_208_i\
        );

    \I__2268\ : InMux
    port map (
            O => \N__9827\,
            I => \N__9824\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__9824\,
            I => \READ_CYCLE_ACTIVE_rep28_i_ess\
        );

    \I__2266\ : IoInMux
    port map (
            O => \N__9821\,
            I => \N__9818\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__9818\,
            I => \N__9815\
        );

    \I__2264\ : IoSpan4Mux
    port map (
            O => \N__9815\,
            I => \N__9812\
        );

    \I__2263\ : Span4Mux_s3_h
    port map (
            O => \N__9812\,
            I => \N__9809\
        );

    \I__2262\ : Span4Mux_v
    port map (
            O => \N__9809\,
            I => \N__9806\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__9806\,
            I => \N_204_i\
        );

    \I__2260\ : InMux
    port map (
            O => \N__9803\,
            I => \N__9800\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__9800\,
            I => \READ_CYCLE_ACTIVE_rep30_i_ess\
        );

    \I__2258\ : IoInMux
    port map (
            O => \N__9797\,
            I => \N__9794\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__9794\,
            I => \N__9791\
        );

    \I__2256\ : IoSpan4Mux
    port map (
            O => \N__9791\,
            I => \N__9788\
        );

    \I__2255\ : IoSpan4Mux
    port map (
            O => \N__9788\,
            I => \N__9785\
        );

    \I__2254\ : Span4Mux_s1_h
    port map (
            O => \N__9785\,
            I => \N__9782\
        );

    \I__2253\ : Odrv4
    port map (
            O => \N__9782\,
            I => \N_210_i\
        );

    \I__2252\ : IoInMux
    port map (
            O => \N__9779\,
            I => \N__9776\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__9776\,
            I => \N__9773\
        );

    \I__2250\ : Span4Mux_s3_h
    port map (
            O => \N__9773\,
            I => \N__9770\
        );

    \I__2249\ : Span4Mux_v
    port map (
            O => \N__9770\,
            I => \N__9767\
        );

    \I__2248\ : Odrv4
    port map (
            O => \N__9767\,
            I => \N_206_i\
        );

    \I__2247\ : IoInMux
    port map (
            O => \N__9764\,
            I => \N__9761\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__9761\,
            I => \N__9758\
        );

    \I__2245\ : Span4Mux_s3_h
    port map (
            O => \N__9758\,
            I => \N__9755\
        );

    \I__2244\ : Span4Mux_v
    port map (
            O => \N__9755\,
            I => \N__9752\
        );

    \I__2243\ : Odrv4
    port map (
            O => \N__9752\,
            I => \N_209_i\
        );

    \I__2242\ : IoInMux
    port map (
            O => \N__9749\,
            I => \N__9746\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__9746\,
            I => \N__9743\
        );

    \I__2240\ : IoSpan4Mux
    port map (
            O => \N__9743\,
            I => \N__9740\
        );

    \I__2239\ : Span4Mux_s3_v
    port map (
            O => \N__9740\,
            I => \N__9737\
        );

    \I__2238\ : Span4Mux_v
    port map (
            O => \N__9737\,
            I => \N__9734\
        );

    \I__2237\ : Odrv4
    port map (
            O => \N__9734\,
            I => \N_207_i\
        );

    \I__2236\ : IoInMux
    port map (
            O => \N__9731\,
            I => \N__9728\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__9728\,
            I => \N__9725\
        );

    \I__2234\ : IoSpan4Mux
    port map (
            O => \N__9725\,
            I => \N__9722\
        );

    \I__2233\ : Span4Mux_s3_v
    port map (
            O => \N__9722\,
            I => \N__9719\
        );

    \I__2232\ : Span4Mux_v
    port map (
            O => \N__9719\,
            I => \N__9716\
        );

    \I__2231\ : Odrv4
    port map (
            O => \N__9716\,
            I => \N_205_i\
        );

    \I__2230\ : InMux
    port map (
            O => \N__9713\,
            I => \N__9710\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__9710\,
            I => \READ_CYCLE_ACTIVE_rep27_i_ess\
        );

    \I__2228\ : InMux
    port map (
            O => \N__9707\,
            I => \N__9704\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__9704\,
            I => \N__9701\
        );

    \I__2226\ : Odrv4
    port map (
            O => \N__9701\,
            I => \READ_CYCLE_ACTIVE_rep25_i_ess\
        );

    \I__2225\ : IoInMux
    port map (
            O => \N__9698\,
            I => \N__9695\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__9695\,
            I => \N__9692\
        );

    \I__2223\ : IoSpan4Mux
    port map (
            O => \N__9692\,
            I => \N__9689\
        );

    \I__2222\ : IoSpan4Mux
    port map (
            O => \N__9689\,
            I => \N__9686\
        );

    \I__2221\ : Span4Mux_s1_h
    port map (
            O => \N__9686\,
            I => \N__9683\
        );

    \I__2220\ : Odrv4
    port map (
            O => \N__9683\,
            I => \N_196_i\
        );

    \I__2219\ : InMux
    port map (
            O => \N__9680\,
            I => \N__9677\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__9677\,
            I => \READ_CYCLE_ACTIVE_rep16_i_ess\
        );

    \I__2217\ : IoInMux
    port map (
            O => \N__9674\,
            I => \N__9671\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__9671\,
            I => \N__9668\
        );

    \I__2215\ : IoSpan4Mux
    port map (
            O => \N__9668\,
            I => \N__9663\
        );

    \I__2214\ : IoInMux
    port map (
            O => \N__9667\,
            I => \N__9660\
        );

    \I__2213\ : IoInMux
    port map (
            O => \N__9666\,
            I => \N__9657\
        );

    \I__2212\ : IoSpan4Mux
    port map (
            O => \N__9663\,
            I => \N__9652\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__9660\,
            I => \N__9652\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__9657\,
            I => \N__9649\
        );

    \I__2209\ : IoSpan4Mux
    port map (
            O => \N__9652\,
            I => \N__9646\
        );

    \I__2208\ : Span12Mux_s0_h
    port map (
            O => \N__9649\,
            I => \N__9643\
        );

    \I__2207\ : Sp12to4
    port map (
            O => \N__9646\,
            I => \N__9639\
        );

    \I__2206\ : Span12Mux_h
    port map (
            O => \N__9643\,
            I => \N__9636\
        );

    \I__2205\ : IoInMux
    port map (
            O => \N__9642\,
            I => \N__9633\
        );

    \I__2204\ : Span12Mux_s9_v
    port map (
            O => \N__9639\,
            I => \N__9630\
        );

    \I__2203\ : Span12Mux_h
    port map (
            O => \N__9636\,
            I => \N__9625\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__9633\,
            I => \N__9625\
        );

    \I__2201\ : Odrv12
    port map (
            O => \N__9630\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__2200\ : Odrv12
    port map (
            O => \N__9625\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__2199\ : InMux
    port map (
            O => \N__9620\,
            I => \N__9617\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__9617\,
            I => \READ_CYCLE_ACTIVE_rep4_i_ess\
        );

    \I__2197\ : IoInMux
    port map (
            O => \N__9614\,
            I => \N__9611\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__9611\,
            I => \N__9608\
        );

    \I__2195\ : Span4Mux_s2_v
    port map (
            O => \N__9608\,
            I => \N__9605\
        );

    \I__2194\ : Span4Mux_v
    port map (
            O => \N__9605\,
            I => \N__9602\
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__9602\,
            I => \N_184_i\
        );

    \I__2192\ : InMux
    port map (
            O => \N__9599\,
            I => \N__9596\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__9596\,
            I => \READ_CYCLE_ACTIVE_rep2_i_ess\
        );

    \I__2190\ : IoInMux
    port map (
            O => \N__9593\,
            I => \N__9590\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__9590\,
            I => \N__9587\
        );

    \I__2188\ : Span4Mux_s2_v
    port map (
            O => \N__9587\,
            I => \N__9584\
        );

    \I__2187\ : Span4Mux_v
    port map (
            O => \N__9584\,
            I => \N__9581\
        );

    \I__2186\ : Odrv4
    port map (
            O => \N__9581\,
            I => \N_182_i\
        );

    \I__2185\ : InMux
    port map (
            O => \N__9578\,
            I => \N__9575\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__9575\,
            I => \READ_CYCLE_ACTIVE_rep0_i_ess\
        );

    \I__2183\ : IoInMux
    port map (
            O => \N__9572\,
            I => \N__9569\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__9569\,
            I => \N__9566\
        );

    \I__2181\ : IoSpan4Mux
    port map (
            O => \N__9566\,
            I => \N__9563\
        );

    \I__2180\ : Span4Mux_s2_v
    port map (
            O => \N__9563\,
            I => \N__9560\
        );

    \I__2179\ : Span4Mux_v
    port map (
            O => \N__9560\,
            I => \N__9557\
        );

    \I__2178\ : Odrv4
    port map (
            O => \N__9557\,
            I => \N_180_i\
        );

    \I__2177\ : InMux
    port map (
            O => \N__9554\,
            I => \N__9551\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__9551\,
            I => \N__9548\
        );

    \I__2175\ : Odrv4
    port map (
            O => \N__9548\,
            I => \READ_CYCLE_ACTIVE_rep7_i_ess\
        );

    \I__2174\ : IoInMux
    port map (
            O => \N__9545\,
            I => \N__9542\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__9542\,
            I => \N__9539\
        );

    \I__2172\ : Span12Mux_s6_v
    port map (
            O => \N__9539\,
            I => \N__9536\
        );

    \I__2171\ : Odrv12
    port map (
            O => \N__9536\,
            I => \N_187_i\
        );

    \I__2170\ : InMux
    port map (
            O => \N__9533\,
            I => \N__9530\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__9530\,
            I => \READ_CYCLE_ACTIVE_rep6_i_ess\
        );

    \I__2168\ : IoInMux
    port map (
            O => \N__9527\,
            I => \N__9524\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__9524\,
            I => \N__9521\
        );

    \I__2166\ : Span4Mux_s2_v
    port map (
            O => \N__9521\,
            I => \N__9518\
        );

    \I__2165\ : Span4Mux_v
    port map (
            O => \N__9518\,
            I => \N__9515\
        );

    \I__2164\ : Odrv4
    port map (
            O => \N__9515\,
            I => \N_186_i\
        );

    \I__2163\ : InMux
    port map (
            O => \N__9512\,
            I => \N__9508\
        );

    \I__2162\ : IoInMux
    port map (
            O => \N__9511\,
            I => \N__9505\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__9508\,
            I => \N__9502\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__9505\,
            I => \N__9499\
        );

    \I__2159\ : Span4Mux_h
    port map (
            O => \N__9502\,
            I => \N__9496\
        );

    \I__2158\ : Span12Mux_s9_h
    port map (
            O => \N__9499\,
            I => \N__9493\
        );

    \I__2157\ : Sp12to4
    port map (
            O => \N__9496\,
            I => \N__9490\
        );

    \I__2156\ : Span12Mux_v
    port map (
            O => \N__9493\,
            I => \N__9487\
        );

    \I__2155\ : Span12Mux_v
    port map (
            O => \N__9490\,
            I => \N__9484\
        );

    \I__2154\ : Span12Mux_h
    port map (
            O => \N__9487\,
            I => \N__9479\
        );

    \I__2153\ : Span12Mux_v
    port map (
            O => \N__9484\,
            I => \N__9479\
        );

    \I__2152\ : Odrv12
    port map (
            O => \N__9479\,
            I => \D_LM_040_in_2\
        );

    \I__2151\ : InMux
    port map (
            O => \N__9476\,
            I => \N__9473\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__9473\,
            I => \N__9470\
        );

    \I__2149\ : Span4Mux_v
    port map (
            O => \N__9470\,
            I => \N__9467\
        );

    \I__2148\ : Span4Mux_h
    port map (
            O => \N__9467\,
            I => \N__9464\
        );

    \I__2147\ : IoSpan4Mux
    port map (
            O => \N__9464\,
            I => \N__9461\
        );

    \I__2146\ : Odrv4
    port map (
            O => \N__9461\,
            I => \D_UU_040_in_2\
        );

    \I__2145\ : IoInMux
    port map (
            O => \N__9458\,
            I => \N__9455\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__9455\,
            I => \N__9452\
        );

    \I__2143\ : IoSpan4Mux
    port map (
            O => \N__9452\,
            I => \N__9449\
        );

    \I__2142\ : IoSpan4Mux
    port map (
            O => \N__9449\,
            I => \N__9446\
        );

    \I__2141\ : IoSpan4Mux
    port map (
            O => \N__9446\,
            I => \N__9443\
        );

    \I__2140\ : Span4Mux_s2_v
    port map (
            O => \N__9443\,
            I => \N__9440\
        );

    \I__2139\ : Span4Mux_v
    port map (
            O => \N__9440\,
            I => \N__9437\
        );

    \I__2138\ : Odrv4
    port map (
            O => \N__9437\,
            I => \un1_D_UU_040_2\
        );

    \I__2137\ : InMux
    port map (
            O => \N__9434\,
            I => \N__9431\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9431\,
            I => \N__9428\
        );

    \I__2135\ : Span4Mux_h
    port map (
            O => \N__9428\,
            I => \N__9425\
        );

    \I__2134\ : Span4Mux_v
    port map (
            O => \N__9425\,
            I => \N__9422\
        );

    \I__2133\ : Span4Mux_h
    port map (
            O => \N__9422\,
            I => \N__9419\
        );

    \I__2132\ : Odrv4
    port map (
            O => \N__9419\,
            I => \D_UU_040_in_0\
        );

    \I__2131\ : IoInMux
    port map (
            O => \N__9416\,
            I => \N__9413\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__9413\,
            I => \N__9409\
        );

    \I__2129\ : InMux
    port map (
            O => \N__9412\,
            I => \N__9406\
        );

    \I__2128\ : IoSpan4Mux
    port map (
            O => \N__9409\,
            I => \N__9403\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__9406\,
            I => \N__9400\
        );

    \I__2126\ : IoSpan4Mux
    port map (
            O => \N__9403\,
            I => \N__9397\
        );

    \I__2125\ : Span4Mux_v
    port map (
            O => \N__9400\,
            I => \N__9394\
        );

    \I__2124\ : Span4Mux_s2_h
    port map (
            O => \N__9397\,
            I => \N__9391\
        );

    \I__2123\ : Sp12to4
    port map (
            O => \N__9394\,
            I => \N__9388\
        );

    \I__2122\ : Sp12to4
    port map (
            O => \N__9391\,
            I => \N__9385\
        );

    \I__2121\ : Span12Mux_h
    port map (
            O => \N__9388\,
            I => \N__9382\
        );

    \I__2120\ : Span12Mux_h
    port map (
            O => \N__9385\,
            I => \N__9379\
        );

    \I__2119\ : Span12Mux_v
    port map (
            O => \N__9382\,
            I => \N__9376\
        );

    \I__2118\ : Span12Mux_h
    port map (
            O => \N__9379\,
            I => \N__9373\
        );

    \I__2117\ : Span12Mux_v
    port map (
            O => \N__9376\,
            I => \N__9370\
        );

    \I__2116\ : Odrv12
    port map (
            O => \N__9373\,
            I => \D_LM_040_in_0\
        );

    \I__2115\ : Odrv12
    port map (
            O => \N__9370\,
            I => \D_LM_040_in_0\
        );

    \I__2114\ : IoInMux
    port map (
            O => \N__9365\,
            I => \N__9362\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__9362\,
            I => \N__9359\
        );

    \I__2112\ : IoSpan4Mux
    port map (
            O => \N__9359\,
            I => \N__9356\
        );

    \I__2111\ : Sp12to4
    port map (
            O => \N__9356\,
            I => \N__9353\
        );

    \I__2110\ : Span12Mux_s6_v
    port map (
            O => \N__9353\,
            I => \N__9350\
        );

    \I__2109\ : Odrv12
    port map (
            O => \N__9350\,
            I => \un1_D_UU_040_0\
        );

    \I__2108\ : IoInMux
    port map (
            O => \N__9347\,
            I => \N__9344\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__9344\,
            I => \N__9341\
        );

    \I__2106\ : IoSpan4Mux
    port map (
            O => \N__9341\,
            I => \N__9338\
        );

    \I__2105\ : IoSpan4Mux
    port map (
            O => \N__9338\,
            I => \N__9334\
        );

    \I__2104\ : InMux
    port map (
            O => \N__9337\,
            I => \N__9331\
        );

    \I__2103\ : Span4Mux_s2_h
    port map (
            O => \N__9334\,
            I => \N__9328\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__9331\,
            I => \N__9325\
        );

    \I__2101\ : Sp12to4
    port map (
            O => \N__9328\,
            I => \N__9322\
        );

    \I__2100\ : Span4Mux_v
    port map (
            O => \N__9325\,
            I => \N__9319\
        );

    \I__2099\ : Span12Mux_h
    port map (
            O => \N__9322\,
            I => \N__9316\
        );

    \I__2098\ : Sp12to4
    port map (
            O => \N__9319\,
            I => \N__9313\
        );

    \I__2097\ : Span12Mux_h
    port map (
            O => \N__9316\,
            I => \N__9310\
        );

    \I__2096\ : Span12Mux_v
    port map (
            O => \N__9313\,
            I => \N__9307\
        );

    \I__2095\ : Odrv12
    port map (
            O => \N__9310\,
            I => \D_LM_040_in_3\
        );

    \I__2094\ : Odrv12
    port map (
            O => \N__9307\,
            I => \D_LM_040_in_3\
        );

    \I__2093\ : InMux
    port map (
            O => \N__9302\,
            I => \N__9299\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__9299\,
            I => \N__9296\
        );

    \I__2091\ : Span4Mux_v
    port map (
            O => \N__9296\,
            I => \N__9293\
        );

    \I__2090\ : Sp12to4
    port map (
            O => \N__9293\,
            I => \N__9290\
        );

    \I__2089\ : Span12Mux_h
    port map (
            O => \N__9290\,
            I => \N__9287\
        );

    \I__2088\ : Odrv12
    port map (
            O => \N__9287\,
            I => \D_UU_040_in_3\
        );

    \I__2087\ : IoInMux
    port map (
            O => \N__9284\,
            I => \N__9281\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__9281\,
            I => \N__9278\
        );

    \I__2085\ : IoSpan4Mux
    port map (
            O => \N__9278\,
            I => \N__9275\
        );

    \I__2084\ : Span4Mux_s0_v
    port map (
            O => \N__9275\,
            I => \N__9272\
        );

    \I__2083\ : Span4Mux_h
    port map (
            O => \N__9272\,
            I => \N__9269\
        );

    \I__2082\ : Sp12to4
    port map (
            O => \N__9269\,
            I => \N__9266\
        );

    \I__2081\ : Span12Mux_h
    port map (
            O => \N__9266\,
            I => \N__9263\
        );

    \I__2080\ : Odrv12
    port map (
            O => \N__9263\,
            I => \un1_D_UU_040_3\
        );

    \I__2079\ : InMux
    port map (
            O => \N__9260\,
            I => \N__9257\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__9257\,
            I => \N__9254\
        );

    \I__2077\ : Span4Mux_v
    port map (
            O => \N__9254\,
            I => \N__9251\
        );

    \I__2076\ : Span4Mux_h
    port map (
            O => \N__9251\,
            I => \N__9248\
        );

    \I__2075\ : Odrv4
    port map (
            O => \N__9248\,
            I => \D_UU_040_in_4\
        );

    \I__2074\ : IoInMux
    port map (
            O => \N__9245\,
            I => \N__9242\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__9242\,
            I => \N__9239\
        );

    \I__2072\ : Span4Mux_s1_h
    port map (
            O => \N__9239\,
            I => \N__9236\
        );

    \I__2071\ : Sp12to4
    port map (
            O => \N__9236\,
            I => \N__9232\
        );

    \I__2070\ : InMux
    port map (
            O => \N__9235\,
            I => \N__9229\
        );

    \I__2069\ : Span12Mux_v
    port map (
            O => \N__9232\,
            I => \N__9226\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__9229\,
            I => \N__9223\
        );

    \I__2067\ : Span12Mux_h
    port map (
            O => \N__9226\,
            I => \N__9220\
        );

    \I__2066\ : Span12Mux_h
    port map (
            O => \N__9223\,
            I => \N__9217\
        );

    \I__2065\ : Span12Mux_h
    port map (
            O => \N__9220\,
            I => \N__9214\
        );

    \I__2064\ : Span12Mux_v
    port map (
            O => \N__9217\,
            I => \N__9211\
        );

    \I__2063\ : Odrv12
    port map (
            O => \N__9214\,
            I => \D_LM_040_in_4\
        );

    \I__2062\ : Odrv12
    port map (
            O => \N__9211\,
            I => \D_LM_040_in_4\
        );

    \I__2061\ : IoInMux
    port map (
            O => \N__9206\,
            I => \N__9203\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__9203\,
            I => \N__9200\
        );

    \I__2059\ : IoSpan4Mux
    port map (
            O => \N__9200\,
            I => \N__9197\
        );

    \I__2058\ : Span4Mux_s2_v
    port map (
            O => \N__9197\,
            I => \N__9194\
        );

    \I__2057\ : Span4Mux_v
    port map (
            O => \N__9194\,
            I => \N__9191\
        );

    \I__2056\ : Sp12to4
    port map (
            O => \N__9191\,
            I => \N__9188\
        );

    \I__2055\ : Odrv12
    port map (
            O => \N__9188\,
            I => \un1_D_UU_040_4\
        );

    \I__2054\ : InMux
    port map (
            O => \N__9185\,
            I => \N__9182\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__9182\,
            I => \N__9179\
        );

    \I__2052\ : Span12Mux_h
    port map (
            O => \N__9179\,
            I => \N__9176\
        );

    \I__2051\ : Odrv12
    port map (
            O => \N__9176\,
            I => \D_UM_040_in_0\
        );

    \I__2050\ : IoInMux
    port map (
            O => \N__9173\,
            I => \N__9170\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__9170\,
            I => \N__9167\
        );

    \I__2048\ : IoSpan4Mux
    port map (
            O => \N__9167\,
            I => \N__9164\
        );

    \I__2047\ : Span4Mux_s2_h
    port map (
            O => \N__9164\,
            I => \N__9160\
        );

    \I__2046\ : InMux
    port map (
            O => \N__9163\,
            I => \N__9157\
        );

    \I__2045\ : Sp12to4
    port map (
            O => \N__9160\,
            I => \N__9154\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__9157\,
            I => \N__9151\
        );

    \I__2043\ : Span12Mux_h
    port map (
            O => \N__9154\,
            I => \N__9148\
        );

    \I__2042\ : Span12Mux_v
    port map (
            O => \N__9151\,
            I => \N__9145\
        );

    \I__2041\ : Span12Mux_h
    port map (
            O => \N__9148\,
            I => \N__9142\
        );

    \I__2040\ : Span12Mux_v
    port map (
            O => \N__9145\,
            I => \N__9139\
        );

    \I__2039\ : Odrv12
    port map (
            O => \N__9142\,
            I => \D_LL_040_in_0\
        );

    \I__2038\ : Odrv12
    port map (
            O => \N__9139\,
            I => \D_LL_040_in_0\
        );

    \I__2037\ : IoInMux
    port map (
            O => \N__9134\,
            I => \N__9131\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__9131\,
            I => \N__9128\
        );

    \I__2035\ : IoSpan4Mux
    port map (
            O => \N__9128\,
            I => \N__9125\
        );

    \I__2034\ : Span4Mux_s2_h
    port map (
            O => \N__9125\,
            I => \N__9122\
        );

    \I__2033\ : Span4Mux_h
    port map (
            O => \N__9122\,
            I => \N__9119\
        );

    \I__2032\ : Span4Mux_h
    port map (
            O => \N__9119\,
            I => \N__9116\
        );

    \I__2031\ : Sp12to4
    port map (
            O => \N__9116\,
            I => \N__9113\
        );

    \I__2030\ : Odrv12
    port map (
            O => \N__9113\,
            I => \un1_D_UM_040_0\
        );

    \I__2029\ : InMux
    port map (
            O => \N__9110\,
            I => \N__9107\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__9107\,
            I => \N__9104\
        );

    \I__2027\ : Span4Mux_h
    port map (
            O => \N__9104\,
            I => \N__9101\
        );

    \I__2026\ : Sp12to4
    port map (
            O => \N__9101\,
            I => \N__9098\
        );

    \I__2025\ : Span12Mux_v
    port map (
            O => \N__9098\,
            I => \N__9095\
        );

    \I__2024\ : Odrv12
    port map (
            O => \N__9095\,
            I => \D_UM_040_in_3\
        );

    \I__2023\ : IoInMux
    port map (
            O => \N__9092\,
            I => \N__9088\
        );

    \I__2022\ : InMux
    port map (
            O => \N__9091\,
            I => \N__9085\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__9088\,
            I => \N__9082\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__9085\,
            I => \N__9079\
        );

    \I__2019\ : Span4Mux_s3_h
    port map (
            O => \N__9082\,
            I => \N__9076\
        );

    \I__2018\ : Span4Mux_v
    port map (
            O => \N__9079\,
            I => \N__9073\
        );

    \I__2017\ : Sp12to4
    port map (
            O => \N__9076\,
            I => \N__9070\
        );

    \I__2016\ : Sp12to4
    port map (
            O => \N__9073\,
            I => \N__9067\
        );

    \I__2015\ : Span12Mux_v
    port map (
            O => \N__9070\,
            I => \N__9064\
        );

    \I__2014\ : Span12Mux_h
    port map (
            O => \N__9067\,
            I => \N__9061\
        );

    \I__2013\ : Span12Mux_h
    port map (
            O => \N__9064\,
            I => \N__9058\
        );

    \I__2012\ : Span12Mux_v
    port map (
            O => \N__9061\,
            I => \N__9055\
        );

    \I__2011\ : Span12Mux_h
    port map (
            O => \N__9058\,
            I => \N__9052\
        );

    \I__2010\ : Span12Mux_v
    port map (
            O => \N__9055\,
            I => \N__9049\
        );

    \I__2009\ : Odrv12
    port map (
            O => \N__9052\,
            I => \D_LL_040_in_3\
        );

    \I__2008\ : Odrv12
    port map (
            O => \N__9049\,
            I => \D_LL_040_in_3\
        );

    \I__2007\ : IoInMux
    port map (
            O => \N__9044\,
            I => \N__9041\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__9041\,
            I => \N__9038\
        );

    \I__2005\ : IoSpan4Mux
    port map (
            O => \N__9038\,
            I => \N__9035\
        );

    \I__2004\ : Span4Mux_s0_h
    port map (
            O => \N__9035\,
            I => \N__9032\
        );

    \I__2003\ : Span4Mux_h
    port map (
            O => \N__9032\,
            I => \N__9029\
        );

    \I__2002\ : Sp12to4
    port map (
            O => \N__9029\,
            I => \N__9026\
        );

    \I__2001\ : Span12Mux_h
    port map (
            O => \N__9026\,
            I => \N__9023\
        );

    \I__2000\ : Odrv12
    port map (
            O => \N__9023\,
            I => \un1_D_UM_040_3\
        );

    \I__1999\ : InMux
    port map (
            O => \N__9020\,
            I => \N__9015\
        );

    \I__1998\ : InMux
    port map (
            O => \N__9019\,
            I => \N__9012\
        );

    \I__1997\ : InMux
    port map (
            O => \N__9018\,
            I => \N__9009\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__9015\,
            I => \N__8994\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__9012\,
            I => \N__8988\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__9009\,
            I => \N__8988\
        );

    \I__1993\ : InMux
    port map (
            O => \N__9008\,
            I => \N__8985\
        );

    \I__1992\ : InMux
    port map (
            O => \N__9007\,
            I => \N__8981\
        );

    \I__1991\ : InMux
    port map (
            O => \N__9006\,
            I => \N__8976\
        );

    \I__1990\ : InMux
    port map (
            O => \N__9005\,
            I => \N__8970\
        );

    \I__1989\ : InMux
    port map (
            O => \N__9004\,
            I => \N__8966\
        );

    \I__1988\ : InMux
    port map (
            O => \N__9003\,
            I => \N__8960\
        );

    \I__1987\ : InMux
    port map (
            O => \N__9002\,
            I => \N__8953\
        );

    \I__1986\ : InMux
    port map (
            O => \N__9001\,
            I => \N__8953\
        );

    \I__1985\ : InMux
    port map (
            O => \N__9000\,
            I => \N__8948\
        );

    \I__1984\ : InMux
    port map (
            O => \N__8999\,
            I => \N__8948\
        );

    \I__1983\ : InMux
    port map (
            O => \N__8998\,
            I => \N__8945\
        );

    \I__1982\ : InMux
    port map (
            O => \N__8997\,
            I => \N__8942\
        );

    \I__1981\ : Span4Mux_v
    port map (
            O => \N__8994\,
            I => \N__8939\
        );

    \I__1980\ : InMux
    port map (
            O => \N__8993\,
            I => \N__8936\
        );

    \I__1979\ : Span4Mux_v
    port map (
            O => \N__8988\,
            I => \N__8932\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__8985\,
            I => \N__8929\
        );

    \I__1977\ : InMux
    port map (
            O => \N__8984\,
            I => \N__8926\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__8981\,
            I => \N__8923\
        );

    \I__1975\ : InMux
    port map (
            O => \N__8980\,
            I => \N__8920\
        );

    \I__1974\ : InMux
    port map (
            O => \N__8979\,
            I => \N__8916\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__8976\,
            I => \N__8912\
        );

    \I__1972\ : InMux
    port map (
            O => \N__8975\,
            I => \N__8909\
        );

    \I__1971\ : InMux
    port map (
            O => \N__8974\,
            I => \N__8906\
        );

    \I__1970\ : InMux
    port map (
            O => \N__8973\,
            I => \N__8903\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__8970\,
            I => \N__8900\
        );

    \I__1968\ : InMux
    port map (
            O => \N__8969\,
            I => \N__8897\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__8966\,
            I => \N__8894\
        );

    \I__1966\ : InMux
    port map (
            O => \N__8965\,
            I => \N__8891\
        );

    \I__1965\ : InMux
    port map (
            O => \N__8964\,
            I => \N__8887\
        );

    \I__1964\ : InMux
    port map (
            O => \N__8963\,
            I => \N__8884\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__8960\,
            I => \N__8881\
        );

    \I__1962\ : InMux
    port map (
            O => \N__8959\,
            I => \N__8878\
        );

    \I__1961\ : InMux
    port map (
            O => \N__8958\,
            I => \N__8875\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__8953\,
            I => \N__8866\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__8948\,
            I => \N__8866\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__8945\,
            I => \N__8866\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__8942\,
            I => \N__8866\
        );

    \I__1956\ : Span4Mux_h
    port map (
            O => \N__8939\,
            I => \N__8861\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__8936\,
            I => \N__8861\
        );

    \I__1954\ : InMux
    port map (
            O => \N__8935\,
            I => \N__8858\
        );

    \I__1953\ : Span4Mux_v
    port map (
            O => \N__8932\,
            I => \N__8851\
        );

    \I__1952\ : Span4Mux_h
    port map (
            O => \N__8929\,
            I => \N__8851\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__8926\,
            I => \N__8851\
        );

    \I__1950\ : Span4Mux_v
    port map (
            O => \N__8923\,
            I => \N__8846\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__8920\,
            I => \N__8846\
        );

    \I__1948\ : InMux
    port map (
            O => \N__8919\,
            I => \N__8843\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__8916\,
            I => \N__8840\
        );

    \I__1946\ : InMux
    port map (
            O => \N__8915\,
            I => \N__8837\
        );

    \I__1945\ : Span4Mux_h
    port map (
            O => \N__8912\,
            I => \N__8832\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__8909\,
            I => \N__8832\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__8906\,
            I => \N__8829\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__8903\,
            I => \N__8826\
        );

    \I__1941\ : Span4Mux_h
    port map (
            O => \N__8900\,
            I => \N__8821\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__8897\,
            I => \N__8821\
        );

    \I__1939\ : Span4Mux_v
    port map (
            O => \N__8894\,
            I => \N__8816\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__8891\,
            I => \N__8816\
        );

    \I__1937\ : InMux
    port map (
            O => \N__8890\,
            I => \N__8813\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__8887\,
            I => \N__8804\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__8884\,
            I => \N__8804\
        );

    \I__1934\ : Span12Mux_h
    port map (
            O => \N__8881\,
            I => \N__8804\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__8878\,
            I => \N__8804\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__8875\,
            I => \N__8801\
        );

    \I__1931\ : Span12Mux_h
    port map (
            O => \N__8866\,
            I => \N__8796\
        );

    \I__1930\ : Sp12to4
    port map (
            O => \N__8861\,
            I => \N__8796\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__8858\,
            I => \N__8793\
        );

    \I__1928\ : Span4Mux_v
    port map (
            O => \N__8851\,
            I => \N__8790\
        );

    \I__1927\ : Span4Mux_h
    port map (
            O => \N__8846\,
            I => \N__8785\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__8843\,
            I => \N__8785\
        );

    \I__1925\ : Span4Mux_h
    port map (
            O => \N__8840\,
            I => \N__8780\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__8837\,
            I => \N__8780\
        );

    \I__1923\ : Span4Mux_v
    port map (
            O => \N__8832\,
            I => \N__8775\
        );

    \I__1922\ : Span4Mux_h
    port map (
            O => \N__8829\,
            I => \N__8775\
        );

    \I__1921\ : Span4Mux_h
    port map (
            O => \N__8826\,
            I => \N__8770\
        );

    \I__1920\ : Span4Mux_v
    port map (
            O => \N__8821\,
            I => \N__8770\
        );

    \I__1919\ : Span4Mux_h
    port map (
            O => \N__8816\,
            I => \N__8767\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__8813\,
            I => \N__8764\
        );

    \I__1917\ : Span12Mux_v
    port map (
            O => \N__8804\,
            I => \N__8758\
        );

    \I__1916\ : Span12Mux_v
    port map (
            O => \N__8801\,
            I => \N__8758\
        );

    \I__1915\ : Span12Mux_v
    port map (
            O => \N__8796\,
            I => \N__8751\
        );

    \I__1914\ : Span12Mux_v
    port map (
            O => \N__8793\,
            I => \N__8751\
        );

    \I__1913\ : Sp12to4
    port map (
            O => \N__8790\,
            I => \N__8751\
        );

    \I__1912\ : Span4Mux_h
    port map (
            O => \N__8785\,
            I => \N__8746\
        );

    \I__1911\ : Span4Mux_v
    port map (
            O => \N__8780\,
            I => \N__8746\
        );

    \I__1910\ : Span4Mux_v
    port map (
            O => \N__8775\,
            I => \N__8737\
        );

    \I__1909\ : Span4Mux_h
    port map (
            O => \N__8770\,
            I => \N__8737\
        );

    \I__1908\ : Span4Mux_v
    port map (
            O => \N__8767\,
            I => \N__8737\
        );

    \I__1907\ : Span4Mux_h
    port map (
            O => \N__8764\,
            I => \N__8737\
        );

    \I__1906\ : InMux
    port map (
            O => \N__8763\,
            I => \N__8734\
        );

    \I__1905\ : Odrv12
    port map (
            O => \N__8758\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1904\ : Odrv12
    port map (
            O => \N__8751\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1903\ : Odrv4
    port map (
            O => \N__8746\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1902\ : Odrv4
    port map (
            O => \N__8737\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__8734\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1900\ : IoInMux
    port map (
            O => \N__8723\,
            I => \N__8720\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__8720\,
            I => \N__8717\
        );

    \I__1898\ : IoSpan4Mux
    port map (
            O => \N__8717\,
            I => \N__8713\
        );

    \I__1897\ : InMux
    port map (
            O => \N__8716\,
            I => \N__8710\
        );

    \I__1896\ : Span4Mux_s3_h
    port map (
            O => \N__8713\,
            I => \N__8707\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__8710\,
            I => \N__8704\
        );

    \I__1894\ : Sp12to4
    port map (
            O => \N__8707\,
            I => \N__8701\
        );

    \I__1893\ : Span4Mux_h
    port map (
            O => \N__8704\,
            I => \N__8698\
        );

    \I__1892\ : Span12Mux_v
    port map (
            O => \N__8701\,
            I => \N__8695\
        );

    \I__1891\ : Sp12to4
    port map (
            O => \N__8698\,
            I => \N__8692\
        );

    \I__1890\ : Span12Mux_h
    port map (
            O => \N__8695\,
            I => \N__8689\
        );

    \I__1889\ : Span12Mux_v
    port map (
            O => \N__8692\,
            I => \N__8686\
        );

    \I__1888\ : Span12Mux_h
    port map (
            O => \N__8689\,
            I => \N__8683\
        );

    \I__1887\ : Span12Mux_v
    port map (
            O => \N__8686\,
            I => \N__8680\
        );

    \I__1886\ : Odrv12
    port map (
            O => \N__8683\,
            I => \D_LL_040_in_7\
        );

    \I__1885\ : Odrv12
    port map (
            O => \N__8680\,
            I => \D_LL_040_in_7\
        );

    \I__1884\ : InMux
    port map (
            O => \N__8675\,
            I => \N__8672\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__8672\,
            I => \N__8669\
        );

    \I__1882\ : Span4Mux_v
    port map (
            O => \N__8669\,
            I => \N__8666\
        );

    \I__1881\ : Span4Mux_v
    port map (
            O => \N__8666\,
            I => \N__8663\
        );

    \I__1880\ : Sp12to4
    port map (
            O => \N__8663\,
            I => \N__8660\
        );

    \I__1879\ : Odrv12
    port map (
            O => \N__8660\,
            I => \D_UM_040_in_7\
        );

    \I__1878\ : IoInMux
    port map (
            O => \N__8657\,
            I => \N__8654\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__8654\,
            I => \N__8651\
        );

    \I__1876\ : Span4Mux_s1_h
    port map (
            O => \N__8651\,
            I => \N__8648\
        );

    \I__1875\ : Span4Mux_h
    port map (
            O => \N__8648\,
            I => \N__8645\
        );

    \I__1874\ : Span4Mux_h
    port map (
            O => \N__8645\,
            I => \N__8642\
        );

    \I__1873\ : Span4Mux_h
    port map (
            O => \N__8642\,
            I => \N__8639\
        );

    \I__1872\ : Span4Mux_h
    port map (
            O => \N__8639\,
            I => \N__8636\
        );

    \I__1871\ : Span4Mux_h
    port map (
            O => \N__8636\,
            I => \N__8633\
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__8633\,
            I => \un1_D_UM_040_7\
        );

    \I__1869\ : InMux
    port map (
            O => \N__8630\,
            I => \N__8627\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__8627\,
            I => \N__8624\
        );

    \I__1867\ : Span4Mux_v
    port map (
            O => \N__8624\,
            I => \N__8621\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__8621\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\
        );

    \I__1865\ : InMux
    port map (
            O => \N__8618\,
            I => \N__8615\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__8615\,
            I => \N__8611\
        );

    \I__1863\ : InMux
    port map (
            O => \N__8614\,
            I => \N__8608\
        );

    \I__1862\ : Span4Mux_v
    port map (
            O => \N__8611\,
            I => \N__8603\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__8608\,
            I => \N__8603\
        );

    \I__1860\ : Sp12to4
    port map (
            O => \N__8603\,
            I => \N__8599\
        );

    \I__1859\ : InMux
    port map (
            O => \N__8602\,
            I => \N__8596\
        );

    \I__1858\ : Span12Mux_v
    port map (
            O => \N__8599\,
            I => \N__8593\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__8596\,
            I => \N__8590\
        );

    \I__1856\ : Span12Mux_h
    port map (
            O => \N__8593\,
            I => \N__8587\
        );

    \I__1855\ : Span12Mux_v
    port map (
            O => \N__8590\,
            I => \N__8584\
        );

    \I__1854\ : Odrv12
    port map (
            O => \N__8587\,
            I => \D_UU_AMIGA_in_5\
        );

    \I__1853\ : Odrv12
    port map (
            O => \N__8584\,
            I => \D_UU_AMIGA_in_5\
        );

    \I__1852\ : IoInMux
    port map (
            O => \N__8579\,
            I => \N__8576\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__8576\,
            I => \N__8573\
        );

    \I__1850\ : Span4Mux_s3_v
    port map (
            O => \N__8573\,
            I => \N__8570\
        );

    \I__1849\ : Span4Mux_v
    port map (
            O => \N__8570\,
            I => \N__8567\
        );

    \I__1848\ : Sp12to4
    port map (
            O => \N__8567\,
            I => \N__8564\
        );

    \I__1847\ : Odrv12
    port map (
            O => \N__8564\,
            I => \un1_D_UU_AMIGA_5\
        );

    \I__1846\ : InMux
    port map (
            O => \N__8561\,
            I => \N__8558\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__8558\,
            I => \N__8555\
        );

    \I__1844\ : Odrv12
    port map (
            O => \N__8555\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\
        );

    \I__1843\ : InMux
    port map (
            O => \N__8552\,
            I => \N__8548\
        );

    \I__1842\ : InMux
    port map (
            O => \N__8551\,
            I => \N__8545\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__8548\,
            I => \N__8541\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__8545\,
            I => \N__8538\
        );

    \I__1839\ : InMux
    port map (
            O => \N__8544\,
            I => \N__8535\
        );

    \I__1838\ : Span4Mux_v
    port map (
            O => \N__8541\,
            I => \N__8532\
        );

    \I__1837\ : Span4Mux_v
    port map (
            O => \N__8538\,
            I => \N__8529\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__8535\,
            I => \N__8524\
        );

    \I__1835\ : Sp12to4
    port map (
            O => \N__8532\,
            I => \N__8524\
        );

    \I__1834\ : Sp12to4
    port map (
            O => \N__8529\,
            I => \N__8521\
        );

    \I__1833\ : Span12Mux_h
    port map (
            O => \N__8524\,
            I => \N__8518\
        );

    \I__1832\ : Span12Mux_h
    port map (
            O => \N__8521\,
            I => \N__8515\
        );

    \I__1831\ : Odrv12
    port map (
            O => \N__8518\,
            I => \D_UU_AMIGA_in_4\
        );

    \I__1830\ : Odrv12
    port map (
            O => \N__8515\,
            I => \D_UU_AMIGA_in_4\
        );

    \I__1829\ : IoInMux
    port map (
            O => \N__8510\,
            I => \N__8507\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__8507\,
            I => \N__8504\
        );

    \I__1827\ : Span4Mux_s2_v
    port map (
            O => \N__8504\,
            I => \N__8501\
        );

    \I__1826\ : Span4Mux_v
    port map (
            O => \N__8501\,
            I => \N__8498\
        );

    \I__1825\ : Sp12to4
    port map (
            O => \N__8498\,
            I => \N__8495\
        );

    \I__1824\ : Odrv12
    port map (
            O => \N__8495\,
            I => \un1_D_UU_AMIGA_4\
        );

    \I__1823\ : InMux
    port map (
            O => \N__8492\,
            I => \N__8488\
        );

    \I__1822\ : InMux
    port map (
            O => \N__8491\,
            I => \N__8484\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__8488\,
            I => \N__8481\
        );

    \I__1820\ : InMux
    port map (
            O => \N__8487\,
            I => \N__8478\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__8484\,
            I => \N__8475\
        );

    \I__1818\ : Span4Mux_v
    port map (
            O => \N__8481\,
            I => \N__8470\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__8478\,
            I => \N__8470\
        );

    \I__1816\ : Span4Mux_v
    port map (
            O => \N__8475\,
            I => \N__8467\
        );

    \I__1815\ : Sp12to4
    port map (
            O => \N__8470\,
            I => \N__8464\
        );

    \I__1814\ : Sp12to4
    port map (
            O => \N__8467\,
            I => \N__8461\
        );

    \I__1813\ : Span12Mux_h
    port map (
            O => \N__8464\,
            I => \N__8458\
        );

    \I__1812\ : Span12Mux_h
    port map (
            O => \N__8461\,
            I => \N__8455\
        );

    \I__1811\ : Odrv12
    port map (
            O => \N__8458\,
            I => \D_UU_AMIGA_in_6\
        );

    \I__1810\ : Odrv12
    port map (
            O => \N__8455\,
            I => \D_UU_AMIGA_in_6\
        );

    \I__1809\ : InMux
    port map (
            O => \N__8450\,
            I => \N__8447\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__8447\,
            I => \N__8434\
        );

    \I__1807\ : InMux
    port map (
            O => \N__8446\,
            I => \N__8427\
        );

    \I__1806\ : InMux
    port map (
            O => \N__8445\,
            I => \N__8427\
        );

    \I__1805\ : InMux
    port map (
            O => \N__8444\,
            I => \N__8427\
        );

    \I__1804\ : InMux
    port map (
            O => \N__8443\,
            I => \N__8422\
        );

    \I__1803\ : InMux
    port map (
            O => \N__8442\,
            I => \N__8422\
        );

    \I__1802\ : InMux
    port map (
            O => \N__8441\,
            I => \N__8417\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8440\,
            I => \N__8417\
        );

    \I__1800\ : InMux
    port map (
            O => \N__8439\,
            I => \N__8412\
        );

    \I__1799\ : InMux
    port map (
            O => \N__8438\,
            I => \N__8412\
        );

    \I__1798\ : InMux
    port map (
            O => \N__8437\,
            I => \N__8409\
        );

    \I__1797\ : Span4Mux_v
    port map (
            O => \N__8434\,
            I => \N__8404\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__8427\,
            I => \N__8393\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__8422\,
            I => \N__8393\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__8417\,
            I => \N__8393\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__8412\,
            I => \N__8393\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__8409\,
            I => \N__8393\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8408\,
            I => \N__8390\
        );

    \I__1790\ : InMux
    port map (
            O => \N__8407\,
            I => \N__8387\
        );

    \I__1789\ : Sp12to4
    port map (
            O => \N__8404\,
            I => \N__8381\
        );

    \I__1788\ : Span4Mux_v
    port map (
            O => \N__8393\,
            I => \N__8374\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__8390\,
            I => \N__8374\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__8387\,
            I => \N__8374\
        );

    \I__1785\ : InMux
    port map (
            O => \N__8386\,
            I => \N__8369\
        );

    \I__1784\ : InMux
    port map (
            O => \N__8385\,
            I => \N__8369\
        );

    \I__1783\ : CascadeMux
    port map (
            O => \N__8384\,
            I => \N__8365\
        );

    \I__1782\ : Span12Mux_h
    port map (
            O => \N__8381\,
            I => \N__8360\
        );

    \I__1781\ : Sp12to4
    port map (
            O => \N__8374\,
            I => \N__8360\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__8369\,
            I => \N__8357\
        );

    \I__1779\ : InMux
    port map (
            O => \N__8368\,
            I => \N__8354\
        );

    \I__1778\ : InMux
    port map (
            O => \N__8365\,
            I => \N__8351\
        );

    \I__1777\ : Odrv12
    port map (
            O => \N__8360\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__1776\ : Odrv4
    port map (
            O => \N__8357\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__8354\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__8351\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__1773\ : InMux
    port map (
            O => \N__8342\,
            I => \N__8339\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__8339\,
            I => \N__8336\
        );

    \I__1771\ : Odrv12
    port map (
            O => \N__8336\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\
        );

    \I__1770\ : IoInMux
    port map (
            O => \N__8333\,
            I => \N__8330\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__8330\,
            I => \N__8327\
        );

    \I__1768\ : Span12Mux_s8_v
    port map (
            O => \N__8327\,
            I => \N__8324\
        );

    \I__1767\ : Span12Mux_h
    port map (
            O => \N__8324\,
            I => \N__8321\
        );

    \I__1766\ : Odrv12
    port map (
            O => \N__8321\,
            I => \un1_D_UU_AMIGA_6\
        );

    \I__1765\ : IoInMux
    port map (
            O => \N__8318\,
            I => \N__8315\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8315\,
            I => \N__8312\
        );

    \I__1763\ : Span4Mux_s2_h
    port map (
            O => \N__8312\,
            I => \N__8309\
        );

    \I__1762\ : Span4Mux_v
    port map (
            O => \N__8309\,
            I => \N__8305\
        );

    \I__1761\ : InMux
    port map (
            O => \N__8308\,
            I => \N__8302\
        );

    \I__1760\ : Sp12to4
    port map (
            O => \N__8305\,
            I => \N__8299\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__8302\,
            I => \N__8296\
        );

    \I__1758\ : Span12Mux_h
    port map (
            O => \N__8299\,
            I => \N__8293\
        );

    \I__1757\ : Span12Mux_s11_v
    port map (
            O => \N__8296\,
            I => \N__8290\
        );

    \I__1756\ : Span12Mux_h
    port map (
            O => \N__8293\,
            I => \N__8287\
        );

    \I__1755\ : Span12Mux_h
    port map (
            O => \N__8290\,
            I => \N__8284\
        );

    \I__1754\ : Odrv12
    port map (
            O => \N__8287\,
            I => \D_LM_040_in_6\
        );

    \I__1753\ : Odrv12
    port map (
            O => \N__8284\,
            I => \D_LM_040_in_6\
        );

    \I__1752\ : InMux
    port map (
            O => \N__8279\,
            I => \N__8276\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__8276\,
            I => \N__8273\
        );

    \I__1750\ : Span4Mux_v
    port map (
            O => \N__8273\,
            I => \N__8270\
        );

    \I__1749\ : Sp12to4
    port map (
            O => \N__8270\,
            I => \N__8267\
        );

    \I__1748\ : Span12Mux_h
    port map (
            O => \N__8267\,
            I => \N__8264\
        );

    \I__1747\ : Odrv12
    port map (
            O => \N__8264\,
            I => \D_UU_040_in_6\
        );

    \I__1746\ : IoInMux
    port map (
            O => \N__8261\,
            I => \N__8258\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__8258\,
            I => \N__8255\
        );

    \I__1744\ : Span4Mux_s3_v
    port map (
            O => \N__8255\,
            I => \N__8252\
        );

    \I__1743\ : Span4Mux_h
    port map (
            O => \N__8252\,
            I => \N__8249\
        );

    \I__1742\ : Sp12to4
    port map (
            O => \N__8249\,
            I => \N__8246\
        );

    \I__1741\ : Span12Mux_h
    port map (
            O => \N__8246\,
            I => \N__8243\
        );

    \I__1740\ : Odrv12
    port map (
            O => \N__8243\,
            I => \un1_D_UU_040_6\
        );

    \I__1739\ : InMux
    port map (
            O => \N__8240\,
            I => \N__8237\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__8237\,
            I => \N__8234\
        );

    \I__1737\ : Span4Mux_v
    port map (
            O => \N__8234\,
            I => \N__8231\
        );

    \I__1736\ : Sp12to4
    port map (
            O => \N__8231\,
            I => \N__8228\
        );

    \I__1735\ : Span12Mux_h
    port map (
            O => \N__8228\,
            I => \N__8225\
        );

    \I__1734\ : Odrv12
    port map (
            O => \N__8225\,
            I => \D_UM_040_in_6\
        );

    \I__1733\ : IoInMux
    port map (
            O => \N__8222\,
            I => \N__8219\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__8219\,
            I => \N__8216\
        );

    \I__1731\ : IoSpan4Mux
    port map (
            O => \N__8216\,
            I => \N__8212\
        );

    \I__1730\ : InMux
    port map (
            O => \N__8215\,
            I => \N__8209\
        );

    \I__1729\ : IoSpan4Mux
    port map (
            O => \N__8212\,
            I => \N__8206\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__8209\,
            I => \N__8203\
        );

    \I__1727\ : Span4Mux_s2_h
    port map (
            O => \N__8206\,
            I => \N__8200\
        );

    \I__1726\ : Span4Mux_v
    port map (
            O => \N__8203\,
            I => \N__8197\
        );

    \I__1725\ : Sp12to4
    port map (
            O => \N__8200\,
            I => \N__8194\
        );

    \I__1724\ : Sp12to4
    port map (
            O => \N__8197\,
            I => \N__8191\
        );

    \I__1723\ : Span12Mux_h
    port map (
            O => \N__8194\,
            I => \N__8188\
        );

    \I__1722\ : Span12Mux_h
    port map (
            O => \N__8191\,
            I => \N__8185\
        );

    \I__1721\ : Span12Mux_h
    port map (
            O => \N__8188\,
            I => \N__8182\
        );

    \I__1720\ : Span12Mux_v
    port map (
            O => \N__8185\,
            I => \N__8179\
        );

    \I__1719\ : Odrv12
    port map (
            O => \N__8182\,
            I => \D_LL_040_in_6\
        );

    \I__1718\ : Odrv12
    port map (
            O => \N__8179\,
            I => \D_LL_040_in_6\
        );

    \I__1717\ : IoInMux
    port map (
            O => \N__8174\,
            I => \N__8171\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__8171\,
            I => \N__8168\
        );

    \I__1715\ : Span12Mux_s2_h
    port map (
            O => \N__8168\,
            I => \N__8165\
        );

    \I__1714\ : Span12Mux_v
    port map (
            O => \N__8165\,
            I => \N__8162\
        );

    \I__1713\ : Span12Mux_h
    port map (
            O => \N__8162\,
            I => \N__8159\
        );

    \I__1712\ : Odrv12
    port map (
            O => \N__8159\,
            I => \un1_D_UM_040_6\
        );

    \I__1711\ : InMux
    port map (
            O => \N__8156\,
            I => \N__8152\
        );

    \I__1710\ : IoInMux
    port map (
            O => \N__8155\,
            I => \N__8149\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__8152\,
            I => \N__8146\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__8149\,
            I => \N__8143\
        );

    \I__1707\ : Span4Mux_v
    port map (
            O => \N__8146\,
            I => \N__8140\
        );

    \I__1706\ : Span4Mux_s2_h
    port map (
            O => \N__8143\,
            I => \N__8137\
        );

    \I__1705\ : Sp12to4
    port map (
            O => \N__8140\,
            I => \N__8134\
        );

    \I__1704\ : Span4Mux_v
    port map (
            O => \N__8137\,
            I => \N__8131\
        );

    \I__1703\ : Span12Mux_h
    port map (
            O => \N__8134\,
            I => \N__8128\
        );

    \I__1702\ : Sp12to4
    port map (
            O => \N__8131\,
            I => \N__8125\
        );

    \I__1701\ : Span12Mux_v
    port map (
            O => \N__8128\,
            I => \N__8122\
        );

    \I__1700\ : Span12Mux_h
    port map (
            O => \N__8125\,
            I => \N__8119\
        );

    \I__1699\ : Span12Mux_v
    port map (
            O => \N__8122\,
            I => \N__8114\
        );

    \I__1698\ : Span12Mux_h
    port map (
            O => \N__8119\,
            I => \N__8114\
        );

    \I__1697\ : Odrv12
    port map (
            O => \N__8114\,
            I => \D_LL_040_in_4\
        );

    \I__1696\ : InMux
    port map (
            O => \N__8111\,
            I => \N__8108\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__8108\,
            I => \N__8105\
        );

    \I__1694\ : Span12Mux_v
    port map (
            O => \N__8105\,
            I => \N__8102\
        );

    \I__1693\ : Span12Mux_h
    port map (
            O => \N__8102\,
            I => \N__8099\
        );

    \I__1692\ : Odrv12
    port map (
            O => \N__8099\,
            I => \D_UM_040_in_4\
        );

    \I__1691\ : IoInMux
    port map (
            O => \N__8096\,
            I => \N__8093\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__8093\,
            I => \N__8090\
        );

    \I__1689\ : Span4Mux_s3_h
    port map (
            O => \N__8090\,
            I => \N__8087\
        );

    \I__1688\ : Span4Mux_h
    port map (
            O => \N__8087\,
            I => \N__8084\
        );

    \I__1687\ : Sp12to4
    port map (
            O => \N__8084\,
            I => \N__8081\
        );

    \I__1686\ : Span12Mux_s7_v
    port map (
            O => \N__8081\,
            I => \N__8078\
        );

    \I__1685\ : Odrv12
    port map (
            O => \N__8078\,
            I => \un1_D_UM_040_4\
        );

    \I__1684\ : InMux
    port map (
            O => \N__8075\,
            I => \N__8072\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__8072\,
            I => \N__8069\
        );

    \I__1682\ : Span4Mux_v
    port map (
            O => \N__8069\,
            I => \N__8066\
        );

    \I__1681\ : Sp12to4
    port map (
            O => \N__8066\,
            I => \N__8063\
        );

    \I__1680\ : Span12Mux_h
    port map (
            O => \N__8063\,
            I => \N__8060\
        );

    \I__1679\ : Odrv12
    port map (
            O => \N__8060\,
            I => \D_UM_040_in_5\
        );

    \I__1678\ : IoInMux
    port map (
            O => \N__8057\,
            I => \N__8054\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__8054\,
            I => \N__8051\
        );

    \I__1676\ : IoSpan4Mux
    port map (
            O => \N__8051\,
            I => \N__8048\
        );

    \I__1675\ : Span4Mux_s2_h
    port map (
            O => \N__8048\,
            I => \N__8044\
        );

    \I__1674\ : InMux
    port map (
            O => \N__8047\,
            I => \N__8041\
        );

    \I__1673\ : Span4Mux_h
    port map (
            O => \N__8044\,
            I => \N__8038\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__8041\,
            I => \N__8035\
        );

    \I__1671\ : Span4Mux_v
    port map (
            O => \N__8038\,
            I => \N__8032\
        );

    \I__1670\ : Sp12to4
    port map (
            O => \N__8035\,
            I => \N__8029\
        );

    \I__1669\ : Sp12to4
    port map (
            O => \N__8032\,
            I => \N__8026\
        );

    \I__1668\ : Span12Mux_v
    port map (
            O => \N__8029\,
            I => \N__8023\
        );

    \I__1667\ : Span12Mux_h
    port map (
            O => \N__8026\,
            I => \N__8018\
        );

    \I__1666\ : Span12Mux_v
    port map (
            O => \N__8023\,
            I => \N__8018\
        );

    \I__1665\ : Span12Mux_h
    port map (
            O => \N__8018\,
            I => \N__8015\
        );

    \I__1664\ : Odrv12
    port map (
            O => \N__8015\,
            I => \D_LL_040_in_5\
        );

    \I__1663\ : IoInMux
    port map (
            O => \N__8012\,
            I => \N__8009\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__8009\,
            I => \N__8006\
        );

    \I__1661\ : IoSpan4Mux
    port map (
            O => \N__8006\,
            I => \N__8003\
        );

    \I__1660\ : IoSpan4Mux
    port map (
            O => \N__8003\,
            I => \N__8000\
        );

    \I__1659\ : IoSpan4Mux
    port map (
            O => \N__8000\,
            I => \N__7997\
        );

    \I__1658\ : IoSpan4Mux
    port map (
            O => \N__7997\,
            I => \N__7994\
        );

    \I__1657\ : Span4Mux_s3_v
    port map (
            O => \N__7994\,
            I => \N__7991\
        );

    \I__1656\ : Odrv4
    port map (
            O => \N__7991\,
            I => \un1_D_UM_040_5\
        );

    \I__1655\ : IoInMux
    port map (
            O => \N__7988\,
            I => \N__7985\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__7985\,
            I => \N__7982\
        );

    \I__1653\ : Span4Mux_s3_h
    port map (
            O => \N__7982\,
            I => \N__7978\
        );

    \I__1652\ : InMux
    port map (
            O => \N__7981\,
            I => \N__7975\
        );

    \I__1651\ : Sp12to4
    port map (
            O => \N__7978\,
            I => \N__7972\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__7975\,
            I => \N__7969\
        );

    \I__1649\ : Span12Mux_v
    port map (
            O => \N__7972\,
            I => \N__7966\
        );

    \I__1648\ : Span12Mux_v
    port map (
            O => \N__7969\,
            I => \N__7963\
        );

    \I__1647\ : Span12Mux_h
    port map (
            O => \N__7966\,
            I => \N__7960\
        );

    \I__1646\ : Span12Mux_v
    port map (
            O => \N__7963\,
            I => \N__7957\
        );

    \I__1645\ : Span12Mux_h
    port map (
            O => \N__7960\,
            I => \N__7954\
        );

    \I__1644\ : Span12Mux_h
    port map (
            O => \N__7957\,
            I => \N__7951\
        );

    \I__1643\ : Odrv12
    port map (
            O => \N__7954\,
            I => \D_LL_040_in_1\
        );

    \I__1642\ : Odrv12
    port map (
            O => \N__7951\,
            I => \D_LL_040_in_1\
        );

    \I__1641\ : InMux
    port map (
            O => \N__7946\,
            I => \N__7943\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__7943\,
            I => \N__7940\
        );

    \I__1639\ : Span4Mux_h
    port map (
            O => \N__7940\,
            I => \N__7937\
        );

    \I__1638\ : Sp12to4
    port map (
            O => \N__7937\,
            I => \N__7934\
        );

    \I__1637\ : Span12Mux_v
    port map (
            O => \N__7934\,
            I => \N__7931\
        );

    \I__1636\ : Odrv12
    port map (
            O => \N__7931\,
            I => \D_UM_040_in_1\
        );

    \I__1635\ : IoInMux
    port map (
            O => \N__7928\,
            I => \N__7925\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__7925\,
            I => \N__7922\
        );

    \I__1633\ : IoSpan4Mux
    port map (
            O => \N__7922\,
            I => \N__7919\
        );

    \I__1632\ : Span4Mux_s0_h
    port map (
            O => \N__7919\,
            I => \N__7916\
        );

    \I__1631\ : Sp12to4
    port map (
            O => \N__7916\,
            I => \N__7913\
        );

    \I__1630\ : Span12Mux_s8_h
    port map (
            O => \N__7913\,
            I => \N__7910\
        );

    \I__1629\ : Odrv12
    port map (
            O => \N__7910\,
            I => \un1_D_UM_040_1\
        );

    \I__1628\ : CEMux
    port map (
            O => \N__7907\,
            I => \N__7900\
        );

    \I__1627\ : CEMux
    port map (
            O => \N__7906\,
            I => \N__7897\
        );

    \I__1626\ : CEMux
    port map (
            O => \N__7905\,
            I => \N__7894\
        );

    \I__1625\ : CEMux
    port map (
            O => \N__7904\,
            I => \N__7891\
        );

    \I__1624\ : CEMux
    port map (
            O => \N__7903\,
            I => \N__7888\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__7900\,
            I => \U111_CYCLE_SM.N_159_0\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__7897\,
            I => \U111_CYCLE_SM.N_159_0\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__7894\,
            I => \U111_CYCLE_SM.N_159_0\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__7891\,
            I => \U111_CYCLE_SM.N_159_0\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__7888\,
            I => \U111_CYCLE_SM.N_159_0\
        );

    \I__1618\ : SRMux
    port map (
            O => \N__7877\,
            I => \N__7873\
        );

    \I__1617\ : SRMux
    port map (
            O => \N__7876\,
            I => \N__7868\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__7873\,
            I => \N__7865\
        );

    \I__1615\ : SRMux
    port map (
            O => \N__7872\,
            I => \N__7862\
        );

    \I__1614\ : SRMux
    port map (
            O => \N__7871\,
            I => \N__7858\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__7868\,
            I => \N__7851\
        );

    \I__1612\ : Span4Mux_h
    port map (
            O => \N__7865\,
            I => \N__7851\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__7862\,
            I => \N__7851\
        );

    \I__1610\ : SRMux
    port map (
            O => \N__7861\,
            I => \N__7848\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__7858\,
            I => \N__7845\
        );

    \I__1608\ : Span4Mux_v
    port map (
            O => \N__7851\,
            I => \N__7840\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__7848\,
            I => \N__7840\
        );

    \I__1606\ : Span4Mux_h
    port map (
            O => \N__7845\,
            I => \N__7837\
        );

    \I__1605\ : Span4Mux_h
    port map (
            O => \N__7840\,
            I => \N__7834\
        );

    \I__1604\ : Odrv4
    port map (
            O => \N__7837\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1\
        );

    \I__1603\ : Odrv4
    port map (
            O => \N__7834\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1\
        );

    \I__1602\ : InMux
    port map (
            O => \N__7829\,
            I => \N__7826\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__7826\,
            I => \N__7823\
        );

    \I__1600\ : Span4Mux_v
    port map (
            O => \N__7823\,
            I => \N__7819\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7822\,
            I => \N__7816\
        );

    \I__1598\ : Odrv4
    port map (
            O => \N__7819\,
            I => \U111_CYCLE_SM.TA_DISZ0\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__7816\,
            I => \U111_CYCLE_SM.TA_DISZ0\
        );

    \I__1596\ : IoInMux
    port map (
            O => \N__7811\,
            I => \N__7808\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__7808\,
            I => \N__7805\
        );

    \I__1594\ : Span4Mux_s2_v
    port map (
            O => \N__7805\,
            I => \N__7802\
        );

    \I__1593\ : Span4Mux_v
    port map (
            O => \N__7802\,
            I => \N__7799\
        );

    \I__1592\ : Span4Mux_v
    port map (
            O => \N__7799\,
            I => \N__7796\
        );

    \I__1591\ : Odrv4
    port map (
            O => \N__7796\,
            I => \TAn_1_i\
        );

    \I__1590\ : InMux
    port map (
            O => \N__7793\,
            I => \N__7790\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__7790\,
            I => \N__7787\
        );

    \I__1588\ : Odrv4
    port map (
            O => \N__7787\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\
        );

    \I__1587\ : InMux
    port map (
            O => \N__7784\,
            I => \N__7780\
        );

    \I__1586\ : InMux
    port map (
            O => \N__7783\,
            I => \N__7777\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__7780\,
            I => \N__7774\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__7777\,
            I => \N__7770\
        );

    \I__1583\ : Span4Mux_v
    port map (
            O => \N__7774\,
            I => \N__7767\
        );

    \I__1582\ : InMux
    port map (
            O => \N__7773\,
            I => \N__7764\
        );

    \I__1581\ : Span4Mux_v
    port map (
            O => \N__7770\,
            I => \N__7761\
        );

    \I__1580\ : Span4Mux_h
    port map (
            O => \N__7767\,
            I => \N__7758\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__7764\,
            I => \N__7755\
        );

    \I__1578\ : Sp12to4
    port map (
            O => \N__7761\,
            I => \N__7752\
        );

    \I__1577\ : Sp12to4
    port map (
            O => \N__7758\,
            I => \N__7747\
        );

    \I__1576\ : Span12Mux_h
    port map (
            O => \N__7755\,
            I => \N__7747\
        );

    \I__1575\ : Span12Mux_h
    port map (
            O => \N__7752\,
            I => \N__7744\
        );

    \I__1574\ : Span12Mux_h
    port map (
            O => \N__7747\,
            I => \N__7741\
        );

    \I__1573\ : Span12Mux_v
    port map (
            O => \N__7744\,
            I => \N__7738\
        );

    \I__1572\ : Odrv12
    port map (
            O => \N__7741\,
            I => \D_UU_AMIGA_in_3\
        );

    \I__1571\ : Odrv12
    port map (
            O => \N__7738\,
            I => \D_UU_AMIGA_in_3\
        );

    \I__1570\ : IoInMux
    port map (
            O => \N__7733\,
            I => \N__7730\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__7730\,
            I => \N__7727\
        );

    \I__1568\ : Span4Mux_s0_v
    port map (
            O => \N__7727\,
            I => \N__7724\
        );

    \I__1567\ : Span4Mux_v
    port map (
            O => \N__7724\,
            I => \N__7721\
        );

    \I__1566\ : Sp12to4
    port map (
            O => \N__7721\,
            I => \N__7718\
        );

    \I__1565\ : Span12Mux_h
    port map (
            O => \N__7718\,
            I => \N__7715\
        );

    \I__1564\ : Odrv12
    port map (
            O => \N__7715\,
            I => \un1_D_UU_AMIGA_3\
        );

    \I__1563\ : InMux
    port map (
            O => \N__7712\,
            I => \N__7709\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__7709\,
            I => \N__7706\
        );

    \I__1561\ : Odrv4
    port map (
            O => \N__7706\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\
        );

    \I__1560\ : InMux
    port map (
            O => \N__7703\,
            I => \N__7699\
        );

    \I__1559\ : InMux
    port map (
            O => \N__7702\,
            I => \N__7695\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__7699\,
            I => \N__7692\
        );

    \I__1557\ : InMux
    port map (
            O => \N__7698\,
            I => \N__7689\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__7695\,
            I => \N__7686\
        );

    \I__1555\ : Span4Mux_v
    port map (
            O => \N__7692\,
            I => \N__7681\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__7689\,
            I => \N__7681\
        );

    \I__1553\ : Span12Mux_v
    port map (
            O => \N__7686\,
            I => \N__7678\
        );

    \I__1552\ : Span4Mux_v
    port map (
            O => \N__7681\,
            I => \N__7675\
        );

    \I__1551\ : Span12Mux_v
    port map (
            O => \N__7678\,
            I => \N__7672\
        );

    \I__1550\ : Sp12to4
    port map (
            O => \N__7675\,
            I => \N__7669\
        );

    \I__1549\ : Span12Mux_h
    port map (
            O => \N__7672\,
            I => \N__7666\
        );

    \I__1548\ : Span12Mux_h
    port map (
            O => \N__7669\,
            I => \N__7663\
        );

    \I__1547\ : Odrv12
    port map (
            O => \N__7666\,
            I => \D_UM_AMIGA_in_3\
        );

    \I__1546\ : Odrv12
    port map (
            O => \N__7663\,
            I => \D_UM_AMIGA_in_3\
        );

    \I__1545\ : IoInMux
    port map (
            O => \N__7658\,
            I => \N__7655\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__7655\,
            I => \N__7652\
        );

    \I__1543\ : IoSpan4Mux
    port map (
            O => \N__7652\,
            I => \N__7649\
        );

    \I__1542\ : Span4Mux_s1_h
    port map (
            O => \N__7649\,
            I => \N__7646\
        );

    \I__1541\ : Sp12to4
    port map (
            O => \N__7646\,
            I => \N__7643\
        );

    \I__1540\ : Span12Mux_h
    port map (
            O => \N__7643\,
            I => \N__7640\
        );

    \I__1539\ : Odrv12
    port map (
            O => \N__7640\,
            I => \un1_D_UM_AMIGA_3\
        );

    \I__1538\ : InMux
    port map (
            O => \N__7637\,
            I => \N__7633\
        );

    \I__1537\ : InMux
    port map (
            O => \N__7636\,
            I => \N__7629\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__7633\,
            I => \N__7626\
        );

    \I__1535\ : InMux
    port map (
            O => \N__7632\,
            I => \N__7623\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__7629\,
            I => \N__7620\
        );

    \I__1533\ : Span4Mux_v
    port map (
            O => \N__7626\,
            I => \N__7615\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__7623\,
            I => \N__7615\
        );

    \I__1531\ : Span12Mux_v
    port map (
            O => \N__7620\,
            I => \N__7612\
        );

    \I__1530\ : Span4Mux_v
    port map (
            O => \N__7615\,
            I => \N__7609\
        );

    \I__1529\ : Span12Mux_h
    port map (
            O => \N__7612\,
            I => \N__7606\
        );

    \I__1528\ : Sp12to4
    port map (
            O => \N__7609\,
            I => \N__7603\
        );

    \I__1527\ : Span12Mux_v
    port map (
            O => \N__7606\,
            I => \N__7600\
        );

    \I__1526\ : Span12Mux_h
    port map (
            O => \N__7603\,
            I => \N__7597\
        );

    \I__1525\ : Odrv12
    port map (
            O => \N__7600\,
            I => \D_UM_AMIGA_in_4\
        );

    \I__1524\ : Odrv12
    port map (
            O => \N__7597\,
            I => \D_UM_AMIGA_in_4\
        );

    \I__1523\ : InMux
    port map (
            O => \N__7592\,
            I => \N__7589\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__7589\,
            I => \N__7586\
        );

    \I__1521\ : Odrv12
    port map (
            O => \N__7586\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\
        );

    \I__1520\ : IoInMux
    port map (
            O => \N__7583\,
            I => \N__7580\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__7580\,
            I => \N__7577\
        );

    \I__1518\ : IoSpan4Mux
    port map (
            O => \N__7577\,
            I => \N__7574\
        );

    \I__1517\ : IoSpan4Mux
    port map (
            O => \N__7574\,
            I => \N__7571\
        );

    \I__1516\ : Span4Mux_s3_v
    port map (
            O => \N__7571\,
            I => \N__7568\
        );

    \I__1515\ : Span4Mux_h
    port map (
            O => \N__7568\,
            I => \N__7565\
        );

    \I__1514\ : Span4Mux_v
    port map (
            O => \N__7565\,
            I => \N__7562\
        );

    \I__1513\ : Odrv4
    port map (
            O => \N__7562\,
            I => \un1_D_UM_AMIGA_4\
        );

    \I__1512\ : IoInMux
    port map (
            O => \N__7559\,
            I => \N__7556\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__7556\,
            I => \N__7553\
        );

    \I__1510\ : IoSpan4Mux
    port map (
            O => \N__7553\,
            I => \N__7550\
        );

    \I__1509\ : Span4Mux_s1_h
    port map (
            O => \N__7550\,
            I => \N__7547\
        );

    \I__1508\ : Sp12to4
    port map (
            O => \N__7547\,
            I => \N__7544\
        );

    \I__1507\ : Span12Mux_h
    port map (
            O => \N__7544\,
            I => \N__7541\
        );

    \I__1506\ : Odrv12
    port map (
            O => \N__7541\,
            I => \un1_D_UM_AMIGA_0\
        );

    \I__1505\ : CascadeMux
    port map (
            O => \N__7538\,
            I => \N__7534\
        );

    \I__1504\ : InMux
    port map (
            O => \N__7537\,
            I => \N__7530\
        );

    \I__1503\ : InMux
    port map (
            O => \N__7534\,
            I => \N__7525\
        );

    \I__1502\ : InMux
    port map (
            O => \N__7533\,
            I => \N__7525\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__7530\,
            I => \U111_CYCLE_SM.LW_TRANSZ0\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__7525\,
            I => \U111_CYCLE_SM.LW_TRANSZ0\
        );

    \I__1499\ : CascadeMux
    port map (
            O => \N__7520\,
            I => \N__7517\
        );

    \I__1498\ : InMux
    port map (
            O => \N__7517\,
            I => \N__7513\
        );

    \I__1497\ : InMux
    port map (
            O => \N__7516\,
            I => \N__7510\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__7513\,
            I => \N__7505\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__7510\,
            I => \N__7505\
        );

    \I__1494\ : Span4Mux_v
    port map (
            O => \N__7505\,
            I => \N__7501\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7504\,
            I => \N__7498\
        );

    \I__1492\ : Sp12to4
    port map (
            O => \N__7501\,
            I => \N__7493\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__7498\,
            I => \N__7493\
        );

    \I__1490\ : Span12Mux_h
    port map (
            O => \N__7493\,
            I => \N__7490\
        );

    \I__1489\ : Span12Mux_v
    port map (
            O => \N__7490\,
            I => \N__7487\
        );

    \I__1488\ : Odrv12
    port map (
            O => \N__7487\,
            I => \PORTSIZE_c\
        );

    \I__1487\ : InMux
    port map (
            O => \N__7484\,
            I => \N__7481\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__7481\,
            I => \N__7477\
        );

    \I__1485\ : InMux
    port map (
            O => \N__7480\,
            I => \N__7474\
        );

    \I__1484\ : Span4Mux_v
    port map (
            O => \N__7477\,
            I => \N__7466\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__7474\,
            I => \N__7466\
        );

    \I__1482\ : InMux
    port map (
            O => \N__7473\,
            I => \N__7463\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7472\,
            I => \N__7460\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7471\,
            I => \N__7457\
        );

    \I__1479\ : Odrv4
    port map (
            O => \N__7466\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__7463\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__7460\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__7457\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7448\,
            I => \N__7444\
        );

    \I__1474\ : InMux
    port map (
            O => \N__7447\,
            I => \N__7440\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__7444\,
            I => \N__7436\
        );

    \I__1472\ : InMux
    port map (
            O => \N__7443\,
            I => \N__7433\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__7440\,
            I => \N__7430\
        );

    \I__1470\ : InMux
    port map (
            O => \N__7439\,
            I => \N__7427\
        );

    \I__1469\ : Odrv4
    port map (
            O => \N__7436\,
            I => \U111_CYCLE_SM.PORT_MISMATCHZ0\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__7433\,
            I => \U111_CYCLE_SM.PORT_MISMATCHZ0\
        );

    \I__1467\ : Odrv4
    port map (
            O => \N__7430\,
            I => \U111_CYCLE_SM.PORT_MISMATCHZ0\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7427\,
            I => \U111_CYCLE_SM.PORT_MISMATCHZ0\
        );

    \I__1465\ : IoInMux
    port map (
            O => \N__7418\,
            I => \N__7415\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__7415\,
            I => \N__7412\
        );

    \I__1463\ : Span12Mux_s3_h
    port map (
            O => \N__7412\,
            I => \N__7409\
        );

    \I__1462\ : Span12Mux_h
    port map (
            O => \N__7409\,
            I => \N__7406\
        );

    \I__1461\ : Odrv12
    port map (
            O => \N__7406\,
            I => \un1_D_UM_AMIGA_2\
        );

    \I__1460\ : InMux
    port map (
            O => \N__7403\,
            I => \N__7400\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__7400\,
            I => \N__7397\
        );

    \I__1458\ : Span4Mux_v
    port map (
            O => \N__7397\,
            I => \N__7394\
        );

    \I__1457\ : Span4Mux_v
    port map (
            O => \N__7394\,
            I => \N__7389\
        );

    \I__1456\ : InMux
    port map (
            O => \N__7393\,
            I => \N__7386\
        );

    \I__1455\ : InMux
    port map (
            O => \N__7392\,
            I => \N__7383\
        );

    \I__1454\ : Sp12to4
    port map (
            O => \N__7389\,
            I => \N__7378\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__7386\,
            I => \N__7378\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__7383\,
            I => \N__7375\
        );

    \I__1451\ : Span12Mux_h
    port map (
            O => \N__7378\,
            I => \N__7372\
        );

    \I__1450\ : Span12Mux_v
    port map (
            O => \N__7375\,
            I => \N__7369\
        );

    \I__1449\ : Span12Mux_v
    port map (
            O => \N__7372\,
            I => \N__7366\
        );

    \I__1448\ : Span12Mux_h
    port map (
            O => \N__7369\,
            I => \N__7363\
        );

    \I__1447\ : Odrv12
    port map (
            O => \N__7366\,
            I => \D_UM_AMIGA_in_6\
        );

    \I__1446\ : Odrv12
    port map (
            O => \N__7363\,
            I => \D_UM_AMIGA_in_6\
        );

    \I__1445\ : InMux
    port map (
            O => \N__7358\,
            I => \N__7355\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__7355\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\
        );

    \I__1443\ : IoInMux
    port map (
            O => \N__7352\,
            I => \N__7349\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__7349\,
            I => \N__7346\
        );

    \I__1441\ : IoSpan4Mux
    port map (
            O => \N__7346\,
            I => \N__7343\
        );

    \I__1440\ : Span4Mux_s2_h
    port map (
            O => \N__7343\,
            I => \N__7340\
        );

    \I__1439\ : Span4Mux_h
    port map (
            O => \N__7340\,
            I => \N__7337\
        );

    \I__1438\ : Sp12to4
    port map (
            O => \N__7337\,
            I => \N__7334\
        );

    \I__1437\ : Odrv12
    port map (
            O => \N__7334\,
            I => \un1_D_UM_AMIGA_6\
        );

    \I__1436\ : InMux
    port map (
            O => \N__7331\,
            I => \N__7328\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__7328\,
            I => \N__7325\
        );

    \I__1434\ : Span4Mux_v
    port map (
            O => \N__7325\,
            I => \N__7320\
        );

    \I__1433\ : InMux
    port map (
            O => \N__7324\,
            I => \N__7317\
        );

    \I__1432\ : InMux
    port map (
            O => \N__7323\,
            I => \N__7314\
        );

    \I__1431\ : Span4Mux_v
    port map (
            O => \N__7320\,
            I => \N__7307\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__7317\,
            I => \N__7307\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__7314\,
            I => \N__7307\
        );

    \I__1428\ : Span4Mux_v
    port map (
            O => \N__7307\,
            I => \N__7304\
        );

    \I__1427\ : Sp12to4
    port map (
            O => \N__7304\,
            I => \N__7301\
        );

    \I__1426\ : Span12Mux_h
    port map (
            O => \N__7301\,
            I => \N__7298\
        );

    \I__1425\ : Odrv12
    port map (
            O => \N__7298\,
            I => \D_UM_AMIGA_in_2\
        );

    \I__1424\ : InMux
    port map (
            O => \N__7295\,
            I => \N__7292\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__7292\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\
        );

    \I__1422\ : InMux
    port map (
            O => \N__7289\,
            I => \N__7286\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__7286\,
            I => \N__7283\
        );

    \I__1420\ : Span4Mux_v
    port map (
            O => \N__7283\,
            I => \N__7278\
        );

    \I__1419\ : InMux
    port map (
            O => \N__7282\,
            I => \N__7275\
        );

    \I__1418\ : InMux
    port map (
            O => \N__7281\,
            I => \N__7272\
        );

    \I__1417\ : Span4Mux_v
    port map (
            O => \N__7278\,
            I => \N__7269\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__7275\,
            I => \N__7266\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__7272\,
            I => \N__7263\
        );

    \I__1414\ : Span4Mux_v
    port map (
            O => \N__7269\,
            I => \N__7256\
        );

    \I__1413\ : Span4Mux_v
    port map (
            O => \N__7266\,
            I => \N__7256\
        );

    \I__1412\ : Span4Mux_v
    port map (
            O => \N__7263\,
            I => \N__7256\
        );

    \I__1411\ : Sp12to4
    port map (
            O => \N__7256\,
            I => \N__7253\
        );

    \I__1410\ : Span12Mux_h
    port map (
            O => \N__7253\,
            I => \N__7250\
        );

    \I__1409\ : Odrv12
    port map (
            O => \N__7250\,
            I => \D_UM_AMIGA_in_0\
        );

    \I__1408\ : InMux
    port map (
            O => \N__7247\,
            I => \N__7244\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__7244\,
            I => \N__7241\
        );

    \I__1406\ : Odrv4
    port map (
            O => \N__7241\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\
        );

    \I__1405\ : InMux
    port map (
            O => \N__7238\,
            I => \N__7235\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__7235\,
            I => \N__7231\
        );

    \I__1403\ : InMux
    port map (
            O => \N__7234\,
            I => \N__7228\
        );

    \I__1402\ : Odrv12
    port map (
            O => \N__7231\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__7228\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__1400\ : InMux
    port map (
            O => \N__7223\,
            I => \N__7220\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__7220\,
            I => \N__7217\
        );

    \I__1398\ : Odrv12
    port map (
            O => \N__7217\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\
        );

    \I__1397\ : InMux
    port map (
            O => \N__7214\,
            I => \N__7211\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__7211\,
            I => \N__7207\
        );

    \I__1395\ : InMux
    port map (
            O => \N__7210\,
            I => \N__7204\
        );

    \I__1394\ : Span4Mux_v
    port map (
            O => \N__7207\,
            I => \N__7201\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__7204\,
            I => \N__7197\
        );

    \I__1392\ : Span4Mux_h
    port map (
            O => \N__7201\,
            I => \N__7194\
        );

    \I__1391\ : InMux
    port map (
            O => \N__7200\,
            I => \N__7191\
        );

    \I__1390\ : Sp12to4
    port map (
            O => \N__7197\,
            I => \N__7188\
        );

    \I__1389\ : Sp12to4
    port map (
            O => \N__7194\,
            I => \N__7185\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__7191\,
            I => \N__7180\
        );

    \I__1387\ : Span12Mux_s11_v
    port map (
            O => \N__7188\,
            I => \N__7180\
        );

    \I__1386\ : Span12Mux_v
    port map (
            O => \N__7185\,
            I => \N__7177\
        );

    \I__1385\ : Span12Mux_h
    port map (
            O => \N__7180\,
            I => \N__7174\
        );

    \I__1384\ : Odrv12
    port map (
            O => \N__7177\,
            I => \D_UM_AMIGA_in_5\
        );

    \I__1383\ : Odrv12
    port map (
            O => \N__7174\,
            I => \D_UM_AMIGA_in_5\
        );

    \I__1382\ : IoInMux
    port map (
            O => \N__7169\,
            I => \N__7166\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__7166\,
            I => \N__7163\
        );

    \I__1380\ : IoSpan4Mux
    port map (
            O => \N__7163\,
            I => \N__7160\
        );

    \I__1379\ : Span4Mux_s3_v
    port map (
            O => \N__7160\,
            I => \N__7157\
        );

    \I__1378\ : Span4Mux_h
    port map (
            O => \N__7157\,
            I => \N__7154\
        );

    \I__1377\ : Span4Mux_h
    port map (
            O => \N__7154\,
            I => \N__7151\
        );

    \I__1376\ : Span4Mux_v
    port map (
            O => \N__7151\,
            I => \N__7148\
        );

    \I__1375\ : Odrv4
    port map (
            O => \N__7148\,
            I => \un1_D_UM_AMIGA_5\
        );

    \I__1374\ : InMux
    port map (
            O => \N__7145\,
            I => \N__7142\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__7142\,
            I => \N__7137\
        );

    \I__1372\ : InMux
    port map (
            O => \N__7141\,
            I => \N__7134\
        );

    \I__1371\ : InMux
    port map (
            O => \N__7140\,
            I => \N__7131\
        );

    \I__1370\ : Span4Mux_v
    port map (
            O => \N__7137\,
            I => \N__7128\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__7134\,
            I => \N__7123\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__7131\,
            I => \N__7123\
        );

    \I__1367\ : Sp12to4
    port map (
            O => \N__7128\,
            I => \N__7120\
        );

    \I__1366\ : Span12Mux_v
    port map (
            O => \N__7123\,
            I => \N__7117\
        );

    \I__1365\ : Span12Mux_v
    port map (
            O => \N__7120\,
            I => \N__7114\
        );

    \I__1364\ : Span12Mux_h
    port map (
            O => \N__7117\,
            I => \N__7111\
        );

    \I__1363\ : Odrv12
    port map (
            O => \N__7114\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__1362\ : Odrv12
    port map (
            O => \N__7111\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__1361\ : InMux
    port map (
            O => \N__7106\,
            I => \N__7103\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__7103\,
            I => \N__7100\
        );

    \I__1359\ : Odrv12
    port map (
            O => \N__7100\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\
        );

    \I__1358\ : IoInMux
    port map (
            O => \N__7097\,
            I => \N__7094\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__7094\,
            I => \N__7091\
        );

    \I__1356\ : IoSpan4Mux
    port map (
            O => \N__7091\,
            I => \N__7088\
        );

    \I__1355\ : Span4Mux_s2_h
    port map (
            O => \N__7088\,
            I => \N__7085\
        );

    \I__1354\ : Span4Mux_h
    port map (
            O => \N__7085\,
            I => \N__7082\
        );

    \I__1353\ : Sp12to4
    port map (
            O => \N__7082\,
            I => \N__7079\
        );

    \I__1352\ : Span12Mux_s7_v
    port map (
            O => \N__7079\,
            I => \N__7076\
        );

    \I__1351\ : Odrv12
    port map (
            O => \N__7076\,
            I => \un1_D_UM_AMIGA_7\
        );

    \I__1350\ : InMux
    port map (
            O => \N__7073\,
            I => \N__7070\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__7070\,
            I => \N__7067\
        );

    \I__1348\ : Span4Mux_v
    port map (
            O => \N__7067\,
            I => \N__7062\
        );

    \I__1347\ : InMux
    port map (
            O => \N__7066\,
            I => \N__7059\
        );

    \I__1346\ : InMux
    port map (
            O => \N__7065\,
            I => \N__7056\
        );

    \I__1345\ : Span4Mux_v
    port map (
            O => \N__7062\,
            I => \N__7053\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__7059\,
            I => \N__7050\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__7056\,
            I => \N__7047\
        );

    \I__1342\ : Span4Mux_v
    port map (
            O => \N__7053\,
            I => \N__7040\
        );

    \I__1341\ : Span4Mux_v
    port map (
            O => \N__7050\,
            I => \N__7040\
        );

    \I__1340\ : Span4Mux_v
    port map (
            O => \N__7047\,
            I => \N__7040\
        );

    \I__1339\ : Sp12to4
    port map (
            O => \N__7040\,
            I => \N__7037\
        );

    \I__1338\ : Span12Mux_h
    port map (
            O => \N__7037\,
            I => \N__7034\
        );

    \I__1337\ : Odrv12
    port map (
            O => \N__7034\,
            I => \D_UU_AMIGA_in_0\
        );

    \I__1336\ : InMux
    port map (
            O => \N__7031\,
            I => \N__7028\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__7028\,
            I => \N__7025\
        );

    \I__1334\ : Odrv12
    port map (
            O => \N__7025\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\
        );

    \I__1333\ : IoInMux
    port map (
            O => \N__7022\,
            I => \N__7019\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__7019\,
            I => \N__7016\
        );

    \I__1331\ : Span12Mux_s9_v
    port map (
            O => \N__7016\,
            I => \N__7013\
        );

    \I__1330\ : Span12Mux_h
    port map (
            O => \N__7013\,
            I => \N__7010\
        );

    \I__1329\ : Odrv12
    port map (
            O => \N__7010\,
            I => \un1_D_UU_AMIGA_0\
        );

    \I__1328\ : InMux
    port map (
            O => \N__7007\,
            I => \N__7004\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__7004\,
            I => \N__7001\
        );

    \I__1326\ : Span4Mux_v
    port map (
            O => \N__7001\,
            I => \N__6998\
        );

    \I__1325\ : Odrv4
    port map (
            O => \N__6998\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\
        );

    \I__1324\ : InMux
    port map (
            O => \N__6995\,
            I => \N__6990\
        );

    \I__1323\ : InMux
    port map (
            O => \N__6994\,
            I => \N__6987\
        );

    \I__1322\ : InMux
    port map (
            O => \N__6993\,
            I => \N__6984\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__6990\,
            I => \N__6981\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__6987\,
            I => \N__6978\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__6984\,
            I => \N__6975\
        );

    \I__1318\ : Span12Mux_v
    port map (
            O => \N__6981\,
            I => \N__6972\
        );

    \I__1317\ : Span12Mux_s7_v
    port map (
            O => \N__6978\,
            I => \N__6969\
        );

    \I__1316\ : Span4Mux_h
    port map (
            O => \N__6975\,
            I => \N__6966\
        );

    \I__1315\ : Span12Mux_h
    port map (
            O => \N__6972\,
            I => \N__6963\
        );

    \I__1314\ : Span12Mux_h
    port map (
            O => \N__6969\,
            I => \N__6958\
        );

    \I__1313\ : Sp12to4
    port map (
            O => \N__6966\,
            I => \N__6958\
        );

    \I__1312\ : Odrv12
    port map (
            O => \N__6963\,
            I => \D_UU_AMIGA_in_7\
        );

    \I__1311\ : Odrv12
    port map (
            O => \N__6958\,
            I => \D_UU_AMIGA_in_7\
        );

    \I__1310\ : IoInMux
    port map (
            O => \N__6953\,
            I => \N__6950\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__6950\,
            I => \N__6947\
        );

    \I__1308\ : Span4Mux_s2_v
    port map (
            O => \N__6947\,
            I => \N__6944\
        );

    \I__1307\ : Span4Mux_v
    port map (
            O => \N__6944\,
            I => \N__6941\
        );

    \I__1306\ : Sp12to4
    port map (
            O => \N__6941\,
            I => \N__6938\
        );

    \I__1305\ : Odrv12
    port map (
            O => \N__6938\,
            I => \un1_D_UU_AMIGA_7\
        );

    \I__1304\ : InMux
    port map (
            O => \N__6935\,
            I => \N__6932\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__6932\,
            I => \N__6929\
        );

    \I__1302\ : Odrv12
    port map (
            O => \N__6929\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\
        );

    \I__1301\ : InMux
    port map (
            O => \N__6926\,
            I => \N__6922\
        );

    \I__1300\ : InMux
    port map (
            O => \N__6925\,
            I => \N__6919\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__6922\,
            I => \N__6915\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__6919\,
            I => \N__6912\
        );

    \I__1297\ : InMux
    port map (
            O => \N__6918\,
            I => \N__6909\
        );

    \I__1296\ : Span4Mux_v
    port map (
            O => \N__6915\,
            I => \N__6906\
        );

    \I__1295\ : Span4Mux_v
    port map (
            O => \N__6912\,
            I => \N__6903\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__6909\,
            I => \N__6898\
        );

    \I__1293\ : Sp12to4
    port map (
            O => \N__6906\,
            I => \N__6898\
        );

    \I__1292\ : Sp12to4
    port map (
            O => \N__6903\,
            I => \N__6895\
        );

    \I__1291\ : Span12Mux_h
    port map (
            O => \N__6898\,
            I => \N__6892\
        );

    \I__1290\ : Span12Mux_h
    port map (
            O => \N__6895\,
            I => \N__6889\
        );

    \I__1289\ : Odrv12
    port map (
            O => \N__6892\,
            I => \D_UU_AMIGA_in_2\
        );

    \I__1288\ : Odrv12
    port map (
            O => \N__6889\,
            I => \D_UU_AMIGA_in_2\
        );

    \I__1287\ : IoInMux
    port map (
            O => \N__6884\,
            I => \N__6881\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__6881\,
            I => \N__6878\
        );

    \I__1285\ : Span4Mux_s0_v
    port map (
            O => \N__6878\,
            I => \N__6875\
        );

    \I__1284\ : Sp12to4
    port map (
            O => \N__6875\,
            I => \N__6872\
        );

    \I__1283\ : Span12Mux_h
    port map (
            O => \N__6872\,
            I => \N__6869\
        );

    \I__1282\ : Odrv12
    port map (
            O => \N__6869\,
            I => \un1_D_UU_AMIGA_2\
        );

    \I__1281\ : CascadeMux
    port map (
            O => \N__6866\,
            I => \N__6863\
        );

    \I__1280\ : InMux
    port map (
            O => \N__6863\,
            I => \N__6860\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__6860\,
            I => \N__6857\
        );

    \I__1278\ : Span4Mux_v
    port map (
            O => \N__6857\,
            I => \N__6854\
        );

    \I__1277\ : Odrv4
    port map (
            O => \N__6854\,
            I => \U111_CYCLE_SM.FLIP_WORD_2\
        );

    \I__1276\ : InMux
    port map (
            O => \N__6851\,
            I => \N__6843\
        );

    \I__1275\ : InMux
    port map (
            O => \N__6850\,
            I => \N__6840\
        );

    \I__1274\ : InMux
    port map (
            O => \N__6849\,
            I => \N__6837\
        );

    \I__1273\ : InMux
    port map (
            O => \N__6848\,
            I => \N__6834\
        );

    \I__1272\ : InMux
    port map (
            O => \N__6847\,
            I => \N__6829\
        );

    \I__1271\ : InMux
    port map (
            O => \N__6846\,
            I => \N__6829\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__6843\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__6840\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__6837\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__6834\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__6829\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1265\ : InMux
    port map (
            O => \N__6818\,
            I => \N__6815\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__6815\,
            I => \U111_CYCLE_SM.N_160\
        );

    \I__1263\ : InMux
    port map (
            O => \N__6812\,
            I => \N__6806\
        );

    \I__1262\ : InMux
    port map (
            O => \N__6811\,
            I => \N__6806\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__6806\,
            I => \N__6803\
        );

    \I__1260\ : Span12Mux_v
    port map (
            O => \N__6803\,
            I => \N__6799\
        );

    \I__1259\ : InMux
    port map (
            O => \N__6802\,
            I => \N__6796\
        );

    \I__1258\ : Odrv12
    port map (
            O => \N__6799\,
            I => \U111_CYCLE_SM.A2_ENZ0\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__6796\,
            I => \U111_CYCLE_SM.A2_ENZ0\
        );

    \I__1256\ : InMux
    port map (
            O => \N__6791\,
            I => \N__6787\
        );

    \I__1255\ : InMux
    port map (
            O => \N__6790\,
            I => \N__6784\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__6787\,
            I => \U111_CYCLE_SM.un1_CYCLE_STATE_1_0\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__6784\,
            I => \U111_CYCLE_SM.un1_CYCLE_STATE_1_0\
        );

    \I__1252\ : InMux
    port map (
            O => \N__6779\,
            I => \N__6775\
        );

    \I__1251\ : InMux
    port map (
            O => \N__6778\,
            I => \N__6772\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__6775\,
            I => \N__6768\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__6772\,
            I => \N__6765\
        );

    \I__1248\ : InMux
    port map (
            O => \N__6771\,
            I => \N__6762\
        );

    \I__1247\ : Span4Mux_h
    port map (
            O => \N__6768\,
            I => \N__6759\
        );

    \I__1246\ : Span4Mux_h
    port map (
            O => \N__6765\,
            I => \N__6754\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__6762\,
            I => \N__6751\
        );

    \I__1244\ : Span4Mux_h
    port map (
            O => \N__6759\,
            I => \N__6748\
        );

    \I__1243\ : InMux
    port map (
            O => \N__6758\,
            I => \N__6743\
        );

    \I__1242\ : InMux
    port map (
            O => \N__6757\,
            I => \N__6743\
        );

    \I__1241\ : Odrv4
    port map (
            O => \N__6754\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1240\ : Odrv4
    port map (
            O => \N__6751\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1239\ : Odrv4
    port map (
            O => \N__6748\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6743\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1237\ : InMux
    port map (
            O => \N__6734\,
            I => \N__6727\
        );

    \I__1236\ : InMux
    port map (
            O => \N__6733\,
            I => \N__6727\
        );

    \I__1235\ : InMux
    port map (
            O => \N__6732\,
            I => \N__6724\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__6727\,
            I => \N__6720\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__6724\,
            I => \N__6714\
        );

    \I__1232\ : InMux
    port map (
            O => \N__6723\,
            I => \N__6711\
        );

    \I__1231\ : Span4Mux_v
    port map (
            O => \N__6720\,
            I => \N__6706\
        );

    \I__1230\ : InMux
    port map (
            O => \N__6719\,
            I => \N__6703\
        );

    \I__1229\ : InMux
    port map (
            O => \N__6718\,
            I => \N__6700\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6717\,
            I => \N__6697\
        );

    \I__1227\ : Span4Mux_v
    port map (
            O => \N__6714\,
            I => \N__6692\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__6711\,
            I => \N__6692\
        );

    \I__1225\ : InMux
    port map (
            O => \N__6710\,
            I => \N__6689\
        );

    \I__1224\ : InMux
    port map (
            O => \N__6709\,
            I => \N__6686\
        );

    \I__1223\ : Sp12to4
    port map (
            O => \N__6706\,
            I => \N__6675\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__6703\,
            I => \N__6675\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__6700\,
            I => \N__6675\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__6697\,
            I => \N__6675\
        );

    \I__1219\ : Sp12to4
    port map (
            O => \N__6692\,
            I => \N__6675\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__6689\,
            I => \N__6672\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__6686\,
            I => \N__6669\
        );

    \I__1216\ : Span12Mux_v
    port map (
            O => \N__6675\,
            I => \N__6666\
        );

    \I__1215\ : Span12Mux_h
    port map (
            O => \N__6672\,
            I => \N__6661\
        );

    \I__1214\ : Span12Mux_s7_h
    port map (
            O => \N__6669\,
            I => \N__6661\
        );

    \I__1213\ : Span12Mux_h
    port map (
            O => \N__6666\,
            I => \N__6658\
        );

    \I__1212\ : Span12Mux_v
    port map (
            O => \N__6661\,
            I => \N__6655\
        );

    \I__1211\ : Odrv12
    port map (
            O => \N__6658\,
            I => \RESETn_c\
        );

    \I__1210\ : Odrv12
    port map (
            O => \N__6655\,
            I => \RESETn_c\
        );

    \I__1209\ : CascadeMux
    port map (
            O => \N__6650\,
            I => \U111_CYCLE_SM.CYCLE_STATE_srsts_i_1_2_cascade_\
        );

    \I__1208\ : InMux
    port map (
            O => \N__6647\,
            I => \N__6640\
        );

    \I__1207\ : InMux
    port map (
            O => \N__6646\,
            I => \N__6640\
        );

    \I__1206\ : InMux
    port map (
            O => \N__6645\,
            I => \N__6637\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__6640\,
            I => \N__6632\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__6637\,
            I => \N__6629\
        );

    \I__1203\ : InMux
    port map (
            O => \N__6636\,
            I => \N__6624\
        );

    \I__1202\ : InMux
    port map (
            O => \N__6635\,
            I => \N__6624\
        );

    \I__1201\ : Odrv4
    port map (
            O => \N__6632\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\
        );

    \I__1200\ : Odrv12
    port map (
            O => \N__6629\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__6624\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\
        );

    \I__1198\ : InMux
    port map (
            O => \N__6617\,
            I => \N__6614\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__6614\,
            I => \N__6610\
        );

    \I__1196\ : InMux
    port map (
            O => \N__6613\,
            I => \N__6607\
        );

    \I__1195\ : Span4Mux_v
    port map (
            O => \N__6610\,
            I => \N__6604\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__6607\,
            I => \N__6601\
        );

    \I__1193\ : Sp12to4
    port map (
            O => \N__6604\,
            I => \N__6597\
        );

    \I__1192\ : Span4Mux_v
    port map (
            O => \N__6601\,
            I => \N__6594\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6600\,
            I => \N__6591\
        );

    \I__1190\ : Span12Mux_h
    port map (
            O => \N__6597\,
            I => \N__6588\
        );

    \I__1189\ : Sp12to4
    port map (
            O => \N__6594\,
            I => \N__6583\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__6591\,
            I => \N__6583\
        );

    \I__1187\ : Span12Mux_v
    port map (
            O => \N__6588\,
            I => \N__6578\
        );

    \I__1186\ : Span12Mux_h
    port map (
            O => \N__6583\,
            I => \N__6578\
        );

    \I__1185\ : Odrv12
    port map (
            O => \N__6578\,
            I => \D_UM_AMIGA_in_1\
        );

    \I__1184\ : InMux
    port map (
            O => \N__6575\,
            I => \N__6572\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__6572\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\
        );

    \I__1182\ : IoInMux
    port map (
            O => \N__6569\,
            I => \N__6566\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__6566\,
            I => \N__6563\
        );

    \I__1180\ : IoSpan4Mux
    port map (
            O => \N__6563\,
            I => \N__6560\
        );

    \I__1179\ : Span4Mux_s2_h
    port map (
            O => \N__6560\,
            I => \N__6557\
        );

    \I__1178\ : Sp12to4
    port map (
            O => \N__6557\,
            I => \N__6554\
        );

    \I__1177\ : Span12Mux_h
    port map (
            O => \N__6554\,
            I => \N__6551\
        );

    \I__1176\ : Odrv12
    port map (
            O => \N__6551\,
            I => \un1_D_UM_AMIGA_1\
        );

    \I__1175\ : InMux
    port map (
            O => \N__6548\,
            I => \N__6545\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__6545\,
            I => \N__6542\
        );

    \I__1173\ : Glb2LocalMux
    port map (
            O => \N__6542\,
            I => \N__6539\
        );

    \I__1172\ : GlobalMux
    port map (
            O => \N__6539\,
            I => \CLK80\
        );

    \I__1171\ : IoInMux
    port map (
            O => \N__6536\,
            I => \N__6533\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__6533\,
            I => \N__6530\
        );

    \I__1169\ : IoSpan4Mux
    port map (
            O => \N__6530\,
            I => \N__6526\
        );

    \I__1168\ : IoInMux
    port map (
            O => \N__6529\,
            I => \N__6523\
        );

    \I__1167\ : Span4Mux_s3_v
    port map (
            O => \N__6526\,
            I => \N__6520\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__6523\,
            I => \N__6517\
        );

    \I__1165\ : Span4Mux_v
    port map (
            O => \N__6520\,
            I => \N__6514\
        );

    \I__1164\ : IoSpan4Mux
    port map (
            O => \N__6517\,
            I => \N__6511\
        );

    \I__1163\ : Span4Mux_v
    port map (
            O => \N__6514\,
            I => \N__6508\
        );

    \I__1162\ : IoSpan4Mux
    port map (
            O => \N__6511\,
            I => \N__6505\
        );

    \I__1161\ : Sp12to4
    port map (
            O => \N__6508\,
            I => \N__6502\
        );

    \I__1160\ : Span4Mux_s3_h
    port map (
            O => \N__6505\,
            I => \N__6499\
        );

    \I__1159\ : Span12Mux_v
    port map (
            O => \N__6502\,
            I => \N__6494\
        );

    \I__1158\ : Sp12to4
    port map (
            O => \N__6499\,
            I => \N__6494\
        );

    \I__1157\ : Odrv12
    port map (
            O => \N__6494\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__1156\ : InMux
    port map (
            O => \N__6491\,
            I => \N__6488\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__6488\,
            I => \N__6485\
        );

    \I__1154\ : Span4Mux_v
    port map (
            O => \N__6485\,
            I => \N__6482\
        );

    \I__1153\ : Sp12to4
    port map (
            O => \N__6482\,
            I => \N__6479\
        );

    \I__1152\ : Span12Mux_h
    port map (
            O => \N__6479\,
            I => \N__6476\
        );

    \I__1151\ : Odrv12
    port map (
            O => \N__6476\,
            I => \D_LM_AMIGA_in_6\
        );

    \I__1150\ : IoInMux
    port map (
            O => \N__6473\,
            I => \N__6470\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__6470\,
            I => \N__6467\
        );

    \I__1148\ : IoSpan4Mux
    port map (
            O => \N__6467\,
            I => \N__6464\
        );

    \I__1147\ : Span4Mux_s3_h
    port map (
            O => \N__6464\,
            I => \N__6461\
        );

    \I__1146\ : Span4Mux_h
    port map (
            O => \N__6461\,
            I => \N__6458\
        );

    \I__1145\ : Sp12to4
    port map (
            O => \N__6458\,
            I => \N__6455\
        );

    \I__1144\ : Odrv12
    port map (
            O => \N__6455\,
            I => \un2_D_LM_AMIGA_6\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__6452\,
            I => \U111_CYCLE_SM.un7_CYCLE_STATE_0_cascade_\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6449\,
            I => \N__6446\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__6446\,
            I => \U111_CYCLE_SM.N_149\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6443\,
            I => \N__6436\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6442\,
            I => \N__6433\
        );

    \I__1138\ : InMux
    port map (
            O => \N__6441\,
            I => \N__6430\
        );

    \I__1137\ : InMux
    port map (
            O => \N__6440\,
            I => \N__6425\
        );

    \I__1136\ : InMux
    port map (
            O => \N__6439\,
            I => \N__6422\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__6436\,
            I => \N__6417\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__6433\,
            I => \N__6417\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__6430\,
            I => \N__6414\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6429\,
            I => \N__6411\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6428\,
            I => \N__6408\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__6425\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6422\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__1128\ : Odrv4
    port map (
            O => \N__6417\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__1127\ : Odrv4
    port map (
            O => \N__6414\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__6411\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__6408\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__1124\ : InMux
    port map (
            O => \N__6395\,
            I => \N__6387\
        );

    \I__1123\ : InMux
    port map (
            O => \N__6394\,
            I => \N__6384\
        );

    \I__1122\ : InMux
    port map (
            O => \N__6393\,
            I => \N__6379\
        );

    \I__1121\ : InMux
    port map (
            O => \N__6392\,
            I => \N__6379\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6391\,
            I => \N__6374\
        );

    \I__1119\ : InMux
    port map (
            O => \N__6390\,
            I => \N__6374\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__6387\,
            I => \N__6369\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__6384\,
            I => \N__6369\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__6379\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__6374\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\
        );

    \I__1114\ : Odrv4
    port map (
            O => \N__6369\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\
        );

    \I__1113\ : CascadeMux
    port map (
            O => \N__6362\,
            I => \N__6359\
        );

    \I__1112\ : InMux
    port map (
            O => \N__6359\,
            I => \N__6354\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6358\,
            I => \N__6351\
        );

    \I__1110\ : InMux
    port map (
            O => \N__6357\,
            I => \N__6348\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__6354\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_0\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__6351\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_0\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__6348\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_0\
        );

    \I__1106\ : CascadeMux
    port map (
            O => \N__6341\,
            I => \U111_CYCLE_SM.N_132_0_cascade_\
        );

    \I__1105\ : InMux
    port map (
            O => \N__6338\,
            I => \N__6334\
        );

    \I__1104\ : InMux
    port map (
            O => \N__6337\,
            I => \N__6331\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__6334\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_1\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__6331\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_1\
        );

    \I__1101\ : CascadeMux
    port map (
            O => \N__6326\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNIGD6KZ0Z_2_cascade_\
        );

    \I__1100\ : CascadeMux
    port map (
            O => \N__6323\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1_cascade_\
        );

    \I__1099\ : InMux
    port map (
            O => \N__6320\,
            I => \N__6317\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__6317\,
            I => \N__6310\
        );

    \I__1097\ : InMux
    port map (
            O => \N__6316\,
            I => \N__6307\
        );

    \I__1096\ : InMux
    port map (
            O => \N__6315\,
            I => \N__6302\
        );

    \I__1095\ : InMux
    port map (
            O => \N__6314\,
            I => \N__6302\
        );

    \I__1094\ : InMux
    port map (
            O => \N__6313\,
            I => \N__6299\
        );

    \I__1093\ : Span4Mux_v
    port map (
            O => \N__6310\,
            I => \N__6292\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__6307\,
            I => \N__6292\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__6302\,
            I => \N__6292\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__6299\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNIGD6KZ0Z_2\
        );

    \I__1089\ : Odrv4
    port map (
            O => \N__6292\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNIGD6KZ0Z_2\
        );

    \I__1088\ : IoInMux
    port map (
            O => \N__6287\,
            I => \N__6282\
        );

    \I__1087\ : InMux
    port map (
            O => \N__6286\,
            I => \N__6277\
        );

    \I__1086\ : InMux
    port map (
            O => \N__6285\,
            I => \N__6277\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__6282\,
            I => \N__6273\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__6277\,
            I => \N__6270\
        );

    \I__1083\ : InMux
    port map (
            O => \N__6276\,
            I => \N__6267\
        );

    \I__1082\ : Span4Mux_s1_v
    port map (
            O => \N__6273\,
            I => \N__6262\
        );

    \I__1081\ : Span4Mux_v
    port map (
            O => \N__6270\,
            I => \N__6257\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__6267\,
            I => \N__6257\
        );

    \I__1079\ : InMux
    port map (
            O => \N__6266\,
            I => \N__6254\
        );

    \I__1078\ : InMux
    port map (
            O => \N__6265\,
            I => \N__6251\
        );

    \I__1077\ : Span4Mux_v
    port map (
            O => \N__6262\,
            I => \N__6248\
        );

    \I__1076\ : Span4Mux_v
    port map (
            O => \N__6257\,
            I => \N__6240\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__6254\,
            I => \N__6240\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__6251\,
            I => \N__6240\
        );

    \I__1073\ : Sp12to4
    port map (
            O => \N__6248\,
            I => \N__6237\
        );

    \I__1072\ : InMux
    port map (
            O => \N__6247\,
            I => \N__6234\
        );

    \I__1071\ : Span4Mux_v
    port map (
            O => \N__6240\,
            I => \N__6231\
        );

    \I__1070\ : Span12Mux_h
    port map (
            O => \N__6237\,
            I => \N__6225\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__6234\,
            I => \N__6225\
        );

    \I__1068\ : Sp12to4
    port map (
            O => \N__6231\,
            I => \N__6222\
        );

    \I__1067\ : InMux
    port map (
            O => \N__6230\,
            I => \N__6219\
        );

    \I__1066\ : Span12Mux_v
    port map (
            O => \N__6225\,
            I => \N__6212\
        );

    \I__1065\ : Span12Mux_h
    port map (
            O => \N__6222\,
            I => \N__6212\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__6219\,
            I => \N__6212\
        );

    \I__1063\ : Span12Mux_v
    port map (
            O => \N__6212\,
            I => \N__6209\
        );

    \I__1062\ : Odrv12
    port map (
            O => \N__6209\,
            I => \TACKn_in\
        );

    \I__1061\ : CascadeMux
    port map (
            O => \N__6206\,
            I => \N__6202\
        );

    \I__1060\ : IoInMux
    port map (
            O => \N__6205\,
            I => \N__6198\
        );

    \I__1059\ : InMux
    port map (
            O => \N__6202\,
            I => \N__6193\
        );

    \I__1058\ : InMux
    port map (
            O => \N__6201\,
            I => \N__6193\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__6198\,
            I => \N__6189\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__6193\,
            I => \N__6186\
        );

    \I__1055\ : InMux
    port map (
            O => \N__6192\,
            I => \N__6183\
        );

    \I__1054\ : Span4Mux_s1_v
    port map (
            O => \N__6189\,
            I => \N__6179\
        );

    \I__1053\ : Span4Mux_v
    port map (
            O => \N__6186\,
            I => \N__6174\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__6183\,
            I => \N__6174\
        );

    \I__1051\ : InMux
    port map (
            O => \N__6182\,
            I => \N__6171\
        );

    \I__1050\ : Span4Mux_v
    port map (
            O => \N__6179\,
            I => \N__6168\
        );

    \I__1049\ : Span4Mux_v
    port map (
            O => \N__6174\,
            I => \N__6162\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__6171\,
            I => \N__6162\
        );

    \I__1047\ : Sp12to4
    port map (
            O => \N__6168\,
            I => \N__6158\
        );

    \I__1046\ : InMux
    port map (
            O => \N__6167\,
            I => \N__6155\
        );

    \I__1045\ : Span4Mux_v
    port map (
            O => \N__6162\,
            I => \N__6152\
        );

    \I__1044\ : InMux
    port map (
            O => \N__6161\,
            I => \N__6149\
        );

    \I__1043\ : Span12Mux_h
    port map (
            O => \N__6158\,
            I => \N__6146\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__6155\,
            I => \N__6139\
        );

    \I__1041\ : Sp12to4
    port map (
            O => \N__6152\,
            I => \N__6139\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__6149\,
            I => \N__6139\
        );

    \I__1039\ : Span12Mux_v
    port map (
            O => \N__6146\,
            I => \N__6134\
        );

    \I__1038\ : Span12Mux_h
    port map (
            O => \N__6139\,
            I => \N__6134\
        );

    \I__1037\ : Span12Mux_v
    port map (
            O => \N__6134\,
            I => \N__6131\
        );

    \I__1036\ : Odrv12
    port map (
            O => \N__6131\,
            I => \TEAn_c\
        );

    \I__1035\ : InMux
    port map (
            O => \N__6128\,
            I => \N__6125\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__6125\,
            I => \N__6122\
        );

    \I__1033\ : Odrv4
    port map (
            O => \N__6122\,
            I => \U111_CYCLE_SM.un7_CYCLE_STATE_0\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__6119\,
            I => \U111_CYCLE_SM.N_160_cascade_\
        );

    \I__1031\ : InMux
    port map (
            O => \N__6116\,
            I => \N__6110\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6115\,
            I => \N__6110\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__6110\,
            I => \N__6107\
        );

    \I__1028\ : Span4Mux_v
    port map (
            O => \N__6107\,
            I => \N__6104\
        );

    \I__1027\ : Sp12to4
    port map (
            O => \N__6104\,
            I => \N__6101\
        );

    \I__1026\ : Span12Mux_h
    port map (
            O => \N__6101\,
            I => \N__6098\
        );

    \I__1025\ : Span12Mux_v
    port map (
            O => \N__6098\,
            I => \N__6095\
        );

    \I__1024\ : Odrv12
    port map (
            O => \N__6095\,
            I => \SIZ_c_1\
        );

    \I__1023\ : CascadeMux
    port map (
            O => \N__6092\,
            I => \N__6088\
        );

    \I__1022\ : InMux
    port map (
            O => \N__6091\,
            I => \N__6083\
        );

    \I__1021\ : InMux
    port map (
            O => \N__6088\,
            I => \N__6083\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__6083\,
            I => \N__6080\
        );

    \I__1019\ : Span4Mux_v
    port map (
            O => \N__6080\,
            I => \N__6077\
        );

    \I__1018\ : Sp12to4
    port map (
            O => \N__6077\,
            I => \N__6074\
        );

    \I__1017\ : Span12Mux_h
    port map (
            O => \N__6074\,
            I => \N__6071\
        );

    \I__1016\ : Span12Mux_v
    port map (
            O => \N__6071\,
            I => \N__6068\
        );

    \I__1015\ : Odrv12
    port map (
            O => \N__6068\,
            I => \SIZ_c_0\
        );

    \I__1014\ : CascadeMux
    port map (
            O => \N__6065\,
            I => \U111_CYCLE_SM.PORT_MISMATCH_2_cascade_\
        );

    \I__1013\ : InMux
    port map (
            O => \N__6062\,
            I => \N__6057\
        );

    \I__1012\ : InMux
    port map (
            O => \N__6061\,
            I => \N__6052\
        );

    \I__1011\ : InMux
    port map (
            O => \N__6060\,
            I => \N__6049\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__6057\,
            I => \N__6046\
        );

    \I__1009\ : InMux
    port map (
            O => \N__6056\,
            I => \N__6043\
        );

    \I__1008\ : InMux
    port map (
            O => \N__6055\,
            I => \N__6040\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__6052\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__6049\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__1005\ : Odrv4
    port map (
            O => \N__6046\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__6043\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__6040\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__1002\ : InMux
    port map (
            O => \N__6029\,
            I => \N__6026\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__6026\,
            I => \U111_CYCLE_SM.N_142_0\
        );

    \I__1000\ : CascadeMux
    port map (
            O => \N__6023\,
            I => \N__6020\
        );

    \I__999\ : InMux
    port map (
            O => \N__6020\,
            I => \N__6017\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__6017\,
            I => \N__6014\
        );

    \I__997\ : Span4Mux_h
    port map (
            O => \N__6014\,
            I => \N__6011\
        );

    \I__996\ : Span4Mux_h
    port map (
            O => \N__6011\,
            I => \N__6007\
        );

    \I__995\ : IoInMux
    port map (
            O => \N__6010\,
            I => \N__6004\
        );

    \I__994\ : Sp12to4
    port map (
            O => \N__6007\,
            I => \N__6001\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__6004\,
            I => \N__5998\
        );

    \I__992\ : Span12Mux_v
    port map (
            O => \N__6001\,
            I => \N__5995\
        );

    \I__991\ : IoSpan4Mux
    port map (
            O => \N__5998\,
            I => \N__5992\
        );

    \I__990\ : Odrv12
    port map (
            O => \N__5995\,
            I => \TBIn_c\
        );

    \I__989\ : Odrv4
    port map (
            O => \N__5992\,
            I => \TBIn_c\
        );

    \I__988\ : InMux
    port map (
            O => \N__5987\,
            I => \N__5983\
        );

    \I__987\ : InMux
    port map (
            O => \N__5986\,
            I => \N__5980\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__5983\,
            I => \N__5976\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__5980\,
            I => \N__5973\
        );

    \I__984\ : InMux
    port map (
            O => \N__5979\,
            I => \N__5970\
        );

    \I__983\ : Span4Mux_v
    port map (
            O => \N__5976\,
            I => \N__5967\
        );

    \I__982\ : Span4Mux_v
    port map (
            O => \N__5973\,
            I => \N__5962\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__5970\,
            I => \N__5962\
        );

    \I__980\ : Span4Mux_v
    port map (
            O => \N__5967\,
            I => \N__5959\
        );

    \I__979\ : Span4Mux_v
    port map (
            O => \N__5962\,
            I => \N__5956\
        );

    \I__978\ : Span4Mux_v
    port map (
            O => \N__5959\,
            I => \N__5953\
        );

    \I__977\ : Span4Mux_h
    port map (
            O => \N__5956\,
            I => \N__5950\
        );

    \I__976\ : Sp12to4
    port map (
            O => \N__5953\,
            I => \N__5945\
        );

    \I__975\ : Sp12to4
    port map (
            O => \N__5950\,
            I => \N__5945\
        );

    \I__974\ : Odrv12
    port map (
            O => \N__5945\,
            I => \D_UU_AMIGA_in_1\
        );

    \I__973\ : InMux
    port map (
            O => \N__5942\,
            I => \N__5939\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__5939\,
            I => \N__5936\
        );

    \I__971\ : Odrv4
    port map (
            O => \N__5936\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\
        );

    \I__970\ : IoInMux
    port map (
            O => \N__5933\,
            I => \N__5930\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__5930\,
            I => \N__5927\
        );

    \I__968\ : Span4Mux_s2_h
    port map (
            O => \N__5927\,
            I => \N__5924\
        );

    \I__967\ : Span4Mux_h
    port map (
            O => \N__5924\,
            I => \N__5921\
        );

    \I__966\ : Sp12to4
    port map (
            O => \N__5921\,
            I => \N__5918\
        );

    \I__965\ : Span12Mux_s8_v
    port map (
            O => \N__5918\,
            I => \N__5915\
        );

    \I__964\ : Odrv12
    port map (
            O => \N__5915\,
            I => \un1_D_UU_AMIGA_1\
        );

    \I__963\ : InMux
    port map (
            O => \N__5912\,
            I => \N__5909\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__5909\,
            I => \N__5906\
        );

    \I__961\ : Span4Mux_v
    port map (
            O => \N__5906\,
            I => \N__5903\
        );

    \I__960\ : Sp12to4
    port map (
            O => \N__5903\,
            I => \N__5900\
        );

    \I__959\ : Span12Mux_h
    port map (
            O => \N__5900\,
            I => \N__5897\
        );

    \I__958\ : Odrv12
    port map (
            O => \N__5897\,
            I => \D_LL_AMIGA_in_2\
        );

    \I__957\ : IoInMux
    port map (
            O => \N__5894\,
            I => \N__5891\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__5891\,
            I => \N__5888\
        );

    \I__955\ : IoSpan4Mux
    port map (
            O => \N__5888\,
            I => \N__5885\
        );

    \I__954\ : IoSpan4Mux
    port map (
            O => \N__5885\,
            I => \N__5882\
        );

    \I__953\ : Span4Mux_s3_h
    port map (
            O => \N__5882\,
            I => \N__5879\
        );

    \I__952\ : Sp12to4
    port map (
            O => \N__5879\,
            I => \N__5876\
        );

    \I__951\ : Odrv12
    port map (
            O => \N__5876\,
            I => \un2_D_LL_AMIGA_2\
        );

    \I__950\ : InMux
    port map (
            O => \N__5873\,
            I => \N__5870\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__5870\,
            I => \N__5866\
        );

    \I__948\ : InMux
    port map (
            O => \N__5869\,
            I => \N__5863\
        );

    \I__947\ : Odrv4
    port map (
            O => \N__5866\,
            I => \U111_CYCLE_SM.TS_ENZ0Z6\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__5863\,
            I => \U111_CYCLE_SM.TS_ENZ0Z6\
        );

    \I__945\ : CascadeMux
    port map (
            O => \N__5858\,
            I => \U111_CYCLE_SM.N_158_cascade_\
        );

    \I__944\ : InMux
    port map (
            O => \N__5855\,
            I => \N__5852\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__5852\,
            I => \U111_CYCLE_SM.N_130_0\
        );

    \I__942\ : CascadeMux
    port map (
            O => \N__5849\,
            I => \N__5845\
        );

    \I__941\ : InMux
    port map (
            O => \N__5848\,
            I => \N__5842\
        );

    \I__940\ : InMux
    port map (
            O => \N__5845\,
            I => \N__5839\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__5842\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__5839\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\
        );

    \I__937\ : CascadeMux
    port map (
            O => \N__5834\,
            I => \N__5831\
        );

    \I__936\ : InMux
    port map (
            O => \N__5831\,
            I => \N__5828\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__5828\,
            I => \U111_CYCLE_SM.TS_EN_6\
        );

    \I__934\ : InMux
    port map (
            O => \N__5825\,
            I => \N__5822\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__5822\,
            I => \N__5819\
        );

    \I__932\ : Sp12to4
    port map (
            O => \N__5819\,
            I => \N__5815\
        );

    \I__931\ : InMux
    port map (
            O => \N__5818\,
            I => \N__5812\
        );

    \I__930\ : Span12Mux_v
    port map (
            O => \N__5815\,
            I => \N__5807\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__5812\,
            I => \N__5807\
        );

    \I__928\ : Span12Mux_h
    port map (
            O => \N__5807\,
            I => \N__5804\
        );

    \I__927\ : Odrv12
    port map (
            O => \N__5804\,
            I => \A_040_c_1\
        );

    \I__926\ : IoInMux
    port map (
            O => \N__5801\,
            I => \N__5798\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__5798\,
            I => \N__5795\
        );

    \I__924\ : Sp12to4
    port map (
            O => \N__5795\,
            I => \N__5792\
        );

    \I__923\ : Span12Mux_v
    port map (
            O => \N__5792\,
            I => \N__5789\
        );

    \I__922\ : Odrv12
    port map (
            O => \N__5789\,
            I => \TSn_c\
        );

    \I__921\ : InMux
    port map (
            O => \N__5786\,
            I => \N__5782\
        );

    \I__920\ : InMux
    port map (
            O => \N__5785\,
            I => \N__5779\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__5782\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__5779\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__917\ : CascadeMux
    port map (
            O => \N__5774\,
            I => \U111_CYCLE_SM.CYCLE_STATE_srsts_i_o2_0_5_cascade_\
        );

    \I__916\ : CascadeMux
    port map (
            O => \N__5771\,
            I => \U111_CYCLE_SM.N_148_cascade_\
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__5768\,
            I => \U111_CYCLE_SM.CYCLE_STATE_srsts_0_1_0_cascade_\
        );

    \I__914\ : InMux
    port map (
            O => \N__5765\,
            I => \N__5762\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__5762\,
            I => \N__5759\
        );

    \I__912\ : Span4Mux_v
    port map (
            O => \N__5759\,
            I => \N__5756\
        );

    \I__911\ : Span4Mux_h
    port map (
            O => \N__5756\,
            I => \N__5753\
        );

    \I__910\ : Sp12to4
    port map (
            O => \N__5753\,
            I => \N__5750\
        );

    \I__909\ : Span12Mux_h
    port map (
            O => \N__5750\,
            I => \N__5747\
        );

    \I__908\ : Odrv12
    port map (
            O => \N__5747\,
            I => \D_UU_040_in_5\
        );

    \I__907\ : IoInMux
    port map (
            O => \N__5744\,
            I => \N__5741\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__5741\,
            I => \N__5738\
        );

    \I__905\ : IoSpan4Mux
    port map (
            O => \N__5738\,
            I => \N__5734\
        );

    \I__904\ : InMux
    port map (
            O => \N__5737\,
            I => \N__5731\
        );

    \I__903\ : IoSpan4Mux
    port map (
            O => \N__5734\,
            I => \N__5728\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__5731\,
            I => \N__5725\
        );

    \I__901\ : Span4Mux_s2_h
    port map (
            O => \N__5728\,
            I => \N__5722\
        );

    \I__900\ : Span4Mux_v
    port map (
            O => \N__5725\,
            I => \N__5719\
        );

    \I__899\ : Sp12to4
    port map (
            O => \N__5722\,
            I => \N__5716\
        );

    \I__898\ : Sp12to4
    port map (
            O => \N__5719\,
            I => \N__5713\
        );

    \I__897\ : Span12Mux_h
    port map (
            O => \N__5716\,
            I => \N__5710\
        );

    \I__896\ : Span12Mux_h
    port map (
            O => \N__5713\,
            I => \N__5707\
        );

    \I__895\ : Span12Mux_h
    port map (
            O => \N__5710\,
            I => \N__5702\
        );

    \I__894\ : Span12Mux_v
    port map (
            O => \N__5707\,
            I => \N__5702\
        );

    \I__893\ : Odrv12
    port map (
            O => \N__5702\,
            I => \D_LM_040_in_5\
        );

    \I__892\ : IoInMux
    port map (
            O => \N__5699\,
            I => \N__5696\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__5696\,
            I => \N__5693\
        );

    \I__890\ : Span4Mux_s2_h
    port map (
            O => \N__5693\,
            I => \N__5690\
        );

    \I__889\ : Span4Mux_v
    port map (
            O => \N__5690\,
            I => \N__5687\
        );

    \I__888\ : Sp12to4
    port map (
            O => \N__5687\,
            I => \N__5684\
        );

    \I__887\ : Odrv12
    port map (
            O => \N__5684\,
            I => \un1_D_UU_040_5\
        );

    \I__886\ : InMux
    port map (
            O => \N__5681\,
            I => \N__5678\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5678\,
            I => \N__5675\
        );

    \I__884\ : Span4Mux_v
    port map (
            O => \N__5675\,
            I => \N__5672\
        );

    \I__883\ : Sp12to4
    port map (
            O => \N__5672\,
            I => \N__5669\
        );

    \I__882\ : Odrv12
    port map (
            O => \N__5669\,
            I => \D_LL_AMIGA_in_6\
        );

    \I__881\ : IoInMux
    port map (
            O => \N__5666\,
            I => \N__5663\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__5663\,
            I => \N__5660\
        );

    \I__879\ : Span4Mux_s2_h
    port map (
            O => \N__5660\,
            I => \N__5657\
        );

    \I__878\ : Span4Mux_v
    port map (
            O => \N__5657\,
            I => \N__5654\
        );

    \I__877\ : Span4Mux_v
    port map (
            O => \N__5654\,
            I => \N__5651\
        );

    \I__876\ : Sp12to4
    port map (
            O => \N__5651\,
            I => \N__5648\
        );

    \I__875\ : Span12Mux_s11_h
    port map (
            O => \N__5648\,
            I => \N__5645\
        );

    \I__874\ : Odrv12
    port map (
            O => \N__5645\,
            I => \un2_D_LL_AMIGA_6\
        );

    \I__873\ : InMux
    port map (
            O => \N__5642\,
            I => \N__5639\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__5639\,
            I => \N__5636\
        );

    \I__871\ : Span4Mux_v
    port map (
            O => \N__5636\,
            I => \N__5633\
        );

    \I__870\ : Sp12to4
    port map (
            O => \N__5633\,
            I => \N__5630\
        );

    \I__869\ : Span12Mux_h
    port map (
            O => \N__5630\,
            I => \N__5627\
        );

    \I__868\ : Odrv12
    port map (
            O => \N__5627\,
            I => \D_LM_AMIGA_in_0\
        );

    \I__867\ : IoInMux
    port map (
            O => \N__5624\,
            I => \N__5621\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__5621\,
            I => \N__5618\
        );

    \I__865\ : IoSpan4Mux
    port map (
            O => \N__5618\,
            I => \N__5615\
        );

    \I__864\ : Sp12to4
    port map (
            O => \N__5615\,
            I => \N__5612\
        );

    \I__863\ : Span12Mux_s7_h
    port map (
            O => \N__5612\,
            I => \N__5609\
        );

    \I__862\ : Span12Mux_h
    port map (
            O => \N__5609\,
            I => \N__5606\
        );

    \I__861\ : Odrv12
    port map (
            O => \N__5606\,
            I => \un2_D_LM_AMIGA_0\
        );

    \I__860\ : InMux
    port map (
            O => \N__5603\,
            I => \N__5600\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__5600\,
            I => \N__5597\
        );

    \I__858\ : Span4Mux_v
    port map (
            O => \N__5597\,
            I => \N__5594\
        );

    \I__857\ : Sp12to4
    port map (
            O => \N__5594\,
            I => \N__5591\
        );

    \I__856\ : Span12Mux_h
    port map (
            O => \N__5591\,
            I => \N__5588\
        );

    \I__855\ : Odrv12
    port map (
            O => \N__5588\,
            I => \D_LL_AMIGA_in_3\
        );

    \I__854\ : IoInMux
    port map (
            O => \N__5585\,
            I => \N__5582\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__5582\,
            I => \N__5579\
        );

    \I__852\ : Span4Mux_s2_h
    port map (
            O => \N__5579\,
            I => \N__5576\
        );

    \I__851\ : Span4Mux_v
    port map (
            O => \N__5576\,
            I => \N__5573\
        );

    \I__850\ : Span4Mux_h
    port map (
            O => \N__5573\,
            I => \N__5570\
        );

    \I__849\ : Sp12to4
    port map (
            O => \N__5570\,
            I => \N__5567\
        );

    \I__848\ : Span12Mux_h
    port map (
            O => \N__5567\,
            I => \N__5564\
        );

    \I__847\ : Odrv12
    port map (
            O => \N__5564\,
            I => \un2_D_LL_AMIGA_3\
        );

    \I__846\ : InMux
    port map (
            O => \N__5561\,
            I => \N__5558\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__5558\,
            I => \N__5555\
        );

    \I__844\ : Span4Mux_v
    port map (
            O => \N__5555\,
            I => \N__5552\
        );

    \I__843\ : Sp12to4
    port map (
            O => \N__5552\,
            I => \N__5549\
        );

    \I__842\ : Span12Mux_h
    port map (
            O => \N__5549\,
            I => \N__5546\
        );

    \I__841\ : Odrv12
    port map (
            O => \N__5546\,
            I => \D_LL_AMIGA_in_4\
        );

    \I__840\ : IoInMux
    port map (
            O => \N__5543\,
            I => \N__5540\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__5540\,
            I => \N__5537\
        );

    \I__838\ : Span12Mux_s6_h
    port map (
            O => \N__5537\,
            I => \N__5534\
        );

    \I__837\ : Span12Mux_h
    port map (
            O => \N__5534\,
            I => \N__5531\
        );

    \I__836\ : Odrv12
    port map (
            O => \N__5531\,
            I => \un2_D_LL_AMIGA_4\
        );

    \I__835\ : InMux
    port map (
            O => \N__5528\,
            I => \N__5525\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__5525\,
            I => \N__5522\
        );

    \I__833\ : Span4Mux_v
    port map (
            O => \N__5522\,
            I => \N__5519\
        );

    \I__832\ : Sp12to4
    port map (
            O => \N__5519\,
            I => \N__5516\
        );

    \I__831\ : Span12Mux_h
    port map (
            O => \N__5516\,
            I => \N__5513\
        );

    \I__830\ : Odrv12
    port map (
            O => \N__5513\,
            I => \D_LM_AMIGA_in_4\
        );

    \I__829\ : IoInMux
    port map (
            O => \N__5510\,
            I => \N__5507\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__5507\,
            I => \N__5504\
        );

    \I__827\ : IoSpan4Mux
    port map (
            O => \N__5504\,
            I => \N__5501\
        );

    \I__826\ : Span4Mux_s2_h
    port map (
            O => \N__5501\,
            I => \N__5498\
        );

    \I__825\ : Span4Mux_h
    port map (
            O => \N__5498\,
            I => \N__5495\
        );

    \I__824\ : Sp12to4
    port map (
            O => \N__5495\,
            I => \N__5492\
        );

    \I__823\ : Span12Mux_h
    port map (
            O => \N__5492\,
            I => \N__5489\
        );

    \I__822\ : Odrv12
    port map (
            O => \N__5489\,
            I => \un2_D_LM_AMIGA_4\
        );

    \I__821\ : IoInMux
    port map (
            O => \N__5486\,
            I => \N__5482\
        );

    \I__820\ : IoInMux
    port map (
            O => \N__5485\,
            I => \N__5479\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__5482\,
            I => \N__5476\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__5479\,
            I => \N__5473\
        );

    \I__817\ : Span4Mux_s2_v
    port map (
            O => \N__5476\,
            I => \N__5470\
        );

    \I__816\ : IoSpan4Mux
    port map (
            O => \N__5473\,
            I => \N__5467\
        );

    \I__815\ : Span4Mux_h
    port map (
            O => \N__5470\,
            I => \N__5464\
        );

    \I__814\ : Span4Mux_s2_v
    port map (
            O => \N__5467\,
            I => \N__5461\
        );

    \I__813\ : Span4Mux_v
    port map (
            O => \N__5464\,
            I => \N__5458\
        );

    \I__812\ : Span4Mux_v
    port map (
            O => \N__5461\,
            I => \N__5455\
        );

    \I__811\ : Odrv4
    port map (
            O => \N__5458\,
            I => \CONSTANT_ONE_NET\
        );

    \I__810\ : Odrv4
    port map (
            O => \N__5455\,
            I => \CONSTANT_ONE_NET\
        );

    \I__809\ : IoInMux
    port map (
            O => \N__5450\,
            I => \N__5447\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__5447\,
            I => \N__5444\
        );

    \I__807\ : Odrv12
    port map (
            O => \N__5444\,
            I => \LBENn_c_i_0\
        );

    \I__806\ : InMux
    port map (
            O => \N__5441\,
            I => \N__5438\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__5438\,
            I => \N__5435\
        );

    \I__804\ : Span4Mux_v
    port map (
            O => \N__5435\,
            I => \N__5432\
        );

    \I__803\ : Sp12to4
    port map (
            O => \N__5432\,
            I => \N__5429\
        );

    \I__802\ : Span12Mux_h
    port map (
            O => \N__5429\,
            I => \N__5426\
        );

    \I__801\ : Odrv12
    port map (
            O => \N__5426\,
            I => \D_LL_AMIGA_in_1\
        );

    \I__800\ : IoInMux
    port map (
            O => \N__5423\,
            I => \N__5420\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__5420\,
            I => \N__5417\
        );

    \I__798\ : IoSpan4Mux
    port map (
            O => \N__5417\,
            I => \N__5414\
        );

    \I__797\ : IoSpan4Mux
    port map (
            O => \N__5414\,
            I => \N__5411\
        );

    \I__796\ : Span4Mux_s2_h
    port map (
            O => \N__5411\,
            I => \N__5408\
        );

    \I__795\ : Sp12to4
    port map (
            O => \N__5408\,
            I => \N__5405\
        );

    \I__794\ : Span12Mux_s9_h
    port map (
            O => \N__5405\,
            I => \N__5402\
        );

    \I__793\ : Odrv12
    port map (
            O => \N__5402\,
            I => \un2_D_LL_AMIGA_1\
        );

    \I__792\ : IoInMux
    port map (
            O => \N__5399\,
            I => \N__5396\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__5396\,
            I => \N__5393\
        );

    \I__790\ : Span4Mux_s1_h
    port map (
            O => \N__5393\,
            I => \N__5390\
        );

    \I__789\ : Span4Mux_h
    port map (
            O => \N__5390\,
            I => \N__5387\
        );

    \I__788\ : Span4Mux_h
    port map (
            O => \N__5387\,
            I => \N__5384\
        );

    \I__787\ : Odrv4
    port map (
            O => \N__5384\,
            I => \un1_D_UU_040_1\
        );

    \I__786\ : InMux
    port map (
            O => \N__5381\,
            I => \N__5378\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__5378\,
            I => \WRITE_CYCLE_ACTIVE_rep0_i_ess\
        );

    \I__784\ : IoInMux
    port map (
            O => \N__5375\,
            I => \N__5372\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__5372\,
            I => \N__5369\
        );

    \I__782\ : IoSpan4Mux
    port map (
            O => \N__5369\,
            I => \N__5366\
        );

    \I__781\ : Span4Mux_s3_v
    port map (
            O => \N__5366\,
            I => \N__5363\
        );

    \I__780\ : Span4Mux_v
    port map (
            O => \N__5363\,
            I => \N__5360\
        );

    \I__779\ : Odrv4
    port map (
            O => \N__5360\,
            I => \N_212_i\
        );

    \I__778\ : InMux
    port map (
            O => \N__5357\,
            I => \N__5354\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__5354\,
            I => \WRITE_CYCLE_ACTIVE_rep4_i_ess\
        );

    \I__776\ : IoInMux
    port map (
            O => \N__5351\,
            I => \N__5348\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__5348\,
            I => \N__5345\
        );

    \I__774\ : IoSpan4Mux
    port map (
            O => \N__5345\,
            I => \N__5342\
        );

    \I__773\ : Span4Mux_s3_v
    port map (
            O => \N__5342\,
            I => \N__5339\
        );

    \I__772\ : Odrv4
    port map (
            O => \N__5339\,
            I => \N_216_i\
        );

    \I__771\ : InMux
    port map (
            O => \N__5336\,
            I => \N__5333\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__5333\,
            I => \WRITE_CYCLE_ACTIVE_rep2_i_ess\
        );

    \I__769\ : IoInMux
    port map (
            O => \N__5330\,
            I => \N__5327\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__5327\,
            I => \N__5324\
        );

    \I__767\ : Span12Mux_s7_v
    port map (
            O => \N__5324\,
            I => \N__5321\
        );

    \I__766\ : Odrv12
    port map (
            O => \N__5321\,
            I => \N_225_i\
        );

    \I__765\ : IoInMux
    port map (
            O => \N__5318\,
            I => \N__5315\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__5315\,
            I => \N__5312\
        );

    \I__763\ : IoSpan4Mux
    port map (
            O => \N__5312\,
            I => \N__5309\
        );

    \I__762\ : Span4Mux_s2_v
    port map (
            O => \N__5309\,
            I => \N__5306\
        );

    \I__761\ : Span4Mux_v
    port map (
            O => \N__5306\,
            I => \N__5303\
        );

    \I__760\ : Odrv4
    port map (
            O => \N__5303\,
            I => \LBENn_c_i\
        );

    \I__759\ : InMux
    port map (
            O => \N__5300\,
            I => \N__5297\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__5297\,
            I => \N__5294\
        );

    \I__757\ : Span4Mux_v
    port map (
            O => \N__5294\,
            I => \N__5291\
        );

    \I__756\ : Span4Mux_h
    port map (
            O => \N__5291\,
            I => \N__5288\
        );

    \I__755\ : Span4Mux_h
    port map (
            O => \N__5288\,
            I => \N__5285\
        );

    \I__754\ : Odrv4
    port map (
            O => \N__5285\,
            I => \D_LL_AMIGA_in_0\
        );

    \I__753\ : IoInMux
    port map (
            O => \N__5282\,
            I => \N__5279\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__5279\,
            I => \N__5276\
        );

    \I__751\ : Span4Mux_s0_h
    port map (
            O => \N__5276\,
            I => \N__5273\
        );

    \I__750\ : Sp12to4
    port map (
            O => \N__5273\,
            I => \N__5270\
        );

    \I__749\ : Span12Mux_s6_v
    port map (
            O => \N__5270\,
            I => \N__5267\
        );

    \I__748\ : Span12Mux_h
    port map (
            O => \N__5267\,
            I => \N__5264\
        );

    \I__747\ : Odrv12
    port map (
            O => \N__5264\,
            I => \un2_D_LL_AMIGA_0\
        );

    \I__746\ : InMux
    port map (
            O => \N__5261\,
            I => \N__5258\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__5258\,
            I => \N__5255\
        );

    \I__744\ : Span12Mux_h
    port map (
            O => \N__5255\,
            I => \N__5252\
        );

    \I__743\ : Odrv12
    port map (
            O => \N__5252\,
            I => \D_LM_AMIGA_in_2\
        );

    \I__742\ : IoInMux
    port map (
            O => \N__5249\,
            I => \N__5246\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__5246\,
            I => \N__5243\
        );

    \I__740\ : Span12Mux_s8_h
    port map (
            O => \N__5243\,
            I => \N__5240\
        );

    \I__739\ : Span12Mux_v
    port map (
            O => \N__5240\,
            I => \N__5237\
        );

    \I__738\ : Odrv12
    port map (
            O => \N__5237\,
            I => \un2_D_LM_AMIGA_2\
        );

    \I__737\ : InMux
    port map (
            O => \N__5234\,
            I => \N__5231\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__5231\,
            I => \WRITE_CYCLE_ACTIVE_rep13_i_ess\
        );

    \I__735\ : IoInMux
    port map (
            O => \N__5228\,
            I => \N__5225\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__5225\,
            I => \N__5222\
        );

    \I__733\ : IoSpan4Mux
    port map (
            O => \N__5222\,
            I => \N__5219\
        );

    \I__732\ : Span4Mux_s2_h
    port map (
            O => \N__5219\,
            I => \N__5216\
        );

    \I__731\ : Sp12to4
    port map (
            O => \N__5216\,
            I => \N__5213\
        );

    \I__730\ : Span12Mux_s11_h
    port map (
            O => \N__5213\,
            I => \N__5210\
        );

    \I__729\ : Span12Mux_h
    port map (
            O => \N__5210\,
            I => \N__5207\
        );

    \I__728\ : Odrv12
    port map (
            O => \N__5207\,
            I => \un2_D_LM_AMIGA_1\
        );

    \I__727\ : InMux
    port map (
            O => \N__5204\,
            I => \N__5201\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__5201\,
            I => \N__5198\
        );

    \I__725\ : Odrv12
    port map (
            O => \N__5198\,
            I => \WRITE_CYCLE_ACTIVE_rep15_i_ess\
        );

    \I__724\ : InMux
    port map (
            O => \N__5195\,
            I => \N__5192\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__5192\,
            I => \N__5189\
        );

    \I__722\ : Odrv12
    port map (
            O => \N__5189\,
            I => \WRITE_CYCLE_ACTIVE_rep3_i_ess\
        );

    \I__721\ : InMux
    port map (
            O => \N__5186\,
            I => \N__5183\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__5183\,
            I => \N__5180\
        );

    \I__719\ : Odrv4
    port map (
            O => \N__5180\,
            I => \WRITE_CYCLE_ACTIVE_rep7_i_ess\
        );

    \I__718\ : InMux
    port map (
            O => \N__5177\,
            I => \N__5174\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__5174\,
            I => \N__5171\
        );

    \I__716\ : Span12Mux_h
    port map (
            O => \N__5171\,
            I => \N__5168\
        );

    \I__715\ : Odrv12
    port map (
            O => \N__5168\,
            I => \D_LM_AMIGA_in_3\
        );

    \I__714\ : IoInMux
    port map (
            O => \N__5165\,
            I => \N__5162\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__5162\,
            I => \N__5159\
        );

    \I__712\ : Span4Mux_s1_h
    port map (
            O => \N__5159\,
            I => \N__5156\
        );

    \I__711\ : Span4Mux_h
    port map (
            O => \N__5156\,
            I => \N__5153\
        );

    \I__710\ : Sp12to4
    port map (
            O => \N__5153\,
            I => \N__5150\
        );

    \I__709\ : Span12Mux_v
    port map (
            O => \N__5150\,
            I => \N__5147\
        );

    \I__708\ : Span12Mux_h
    port map (
            O => \N__5147\,
            I => \N__5144\
        );

    \I__707\ : Odrv12
    port map (
            O => \N__5144\,
            I => \un2_D_LM_AMIGA_3\
        );

    \I__706\ : InMux
    port map (
            O => \N__5141\,
            I => \N__5138\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__5138\,
            I => \N__5135\
        );

    \I__704\ : Span4Mux_v
    port map (
            O => \N__5135\,
            I => \N__5132\
        );

    \I__703\ : Sp12to4
    port map (
            O => \N__5132\,
            I => \N__5129\
        );

    \I__702\ : Odrv12
    port map (
            O => \N__5129\,
            I => \D_LM_AMIGA_in_5\
        );

    \I__701\ : IoInMux
    port map (
            O => \N__5126\,
            I => \N__5123\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__5123\,
            I => \N__5120\
        );

    \I__699\ : IoSpan4Mux
    port map (
            O => \N__5120\,
            I => \N__5117\
        );

    \I__698\ : Span4Mux_s3_h
    port map (
            O => \N__5117\,
            I => \N__5114\
        );

    \I__697\ : Span4Mux_v
    port map (
            O => \N__5114\,
            I => \N__5111\
        );

    \I__696\ : Sp12to4
    port map (
            O => \N__5111\,
            I => \N__5108\
        );

    \I__695\ : Span12Mux_h
    port map (
            O => \N__5108\,
            I => \N__5105\
        );

    \I__694\ : Odrv12
    port map (
            O => \N__5105\,
            I => \un2_D_LM_AMIGA_5\
        );

    \I__693\ : IoInMux
    port map (
            O => \N__5102\,
            I => \N__5099\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__5099\,
            I => \N__5096\
        );

    \I__691\ : Span4Mux_s1_v
    port map (
            O => \N__5096\,
            I => \N__5093\
        );

    \I__690\ : Span4Mux_h
    port map (
            O => \N__5093\,
            I => \N__5090\
        );

    \I__689\ : Span4Mux_v
    port map (
            O => \N__5090\,
            I => \N__5087\
        );

    \I__688\ : Odrv4
    port map (
            O => \N__5087\,
            I => \N_214_i\
        );

    \I__687\ : InMux
    port map (
            O => \N__5084\,
            I => \N__5081\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__5081\,
            I => \N__5078\
        );

    \I__685\ : Span4Mux_v
    port map (
            O => \N__5078\,
            I => \N__5075\
        );

    \I__684\ : Span4Mux_v
    port map (
            O => \N__5075\,
            I => \N__5072\
        );

    \I__683\ : Sp12to4
    port map (
            O => \N__5072\,
            I => \N__5069\
        );

    \I__682\ : Span12Mux_h
    port map (
            O => \N__5069\,
            I => \N__5066\
        );

    \I__681\ : Odrv12
    port map (
            O => \N__5066\,
            I => \D_UU_040_in_1\
        );

    \I__680\ : InMux
    port map (
            O => \N__5063\,
            I => \N__5059\
        );

    \I__679\ : IoInMux
    port map (
            O => \N__5062\,
            I => \N__5056\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__5059\,
            I => \N__5053\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__5056\,
            I => \N__5050\
        );

    \I__676\ : Span4Mux_v
    port map (
            O => \N__5053\,
            I => \N__5047\
        );

    \I__675\ : Span4Mux_s3_h
    port map (
            O => \N__5050\,
            I => \N__5044\
        );

    \I__674\ : Span4Mux_h
    port map (
            O => \N__5047\,
            I => \N__5041\
        );

    \I__673\ : Sp12to4
    port map (
            O => \N__5044\,
            I => \N__5038\
        );

    \I__672\ : Span4Mux_v
    port map (
            O => \N__5041\,
            I => \N__5035\
        );

    \I__671\ : Span12Mux_v
    port map (
            O => \N__5038\,
            I => \N__5032\
        );

    \I__670\ : Sp12to4
    port map (
            O => \N__5035\,
            I => \N__5029\
        );

    \I__669\ : Span12Mux_h
    port map (
            O => \N__5032\,
            I => \N__5026\
        );

    \I__668\ : Span12Mux_h
    port map (
            O => \N__5029\,
            I => \N__5023\
        );

    \I__667\ : Span12Mux_h
    port map (
            O => \N__5026\,
            I => \N__5018\
        );

    \I__666\ : Span12Mux_v
    port map (
            O => \N__5023\,
            I => \N__5018\
        );

    \I__665\ : Odrv12
    port map (
            O => \N__5018\,
            I => \D_LM_040_in_1\
        );

    \I__664\ : InMux
    port map (
            O => \N__5015\,
            I => \N__5012\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__5012\,
            I => \N__5009\
        );

    \I__662\ : Span4Mux_v
    port map (
            O => \N__5009\,
            I => \N__5006\
        );

    \I__661\ : Span4Mux_h
    port map (
            O => \N__5006\,
            I => \N__5003\
        );

    \I__660\ : Odrv4
    port map (
            O => \N__5003\,
            I => \D_LM_AMIGA_in_7\
        );

    \I__659\ : IoInMux
    port map (
            O => \N__5000\,
            I => \N__4997\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__4997\,
            I => \N__4994\
        );

    \I__657\ : Span12Mux_s9_h
    port map (
            O => \N__4994\,
            I => \N__4991\
        );

    \I__656\ : Span12Mux_h
    port map (
            O => \N__4991\,
            I => \N__4988\
        );

    \I__655\ : Odrv12
    port map (
            O => \N__4988\,
            I => \un2_D_LM_AMIGA_7\
        );

    \I__654\ : InMux
    port map (
            O => \N__4985\,
            I => \N__4982\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__4982\,
            I => \N__4979\
        );

    \I__652\ : Span4Mux_v
    port map (
            O => \N__4979\,
            I => \N__4976\
        );

    \I__651\ : Odrv4
    port map (
            O => \N__4976\,
            I => \WRITE_CYCLE_ACTIVE_rep12_i_ess\
        );

    \I__650\ : InMux
    port map (
            O => \N__4973\,
            I => \N__4970\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__4970\,
            I => \N__4967\
        );

    \I__648\ : Odrv4
    port map (
            O => \N__4967\,
            I => \WRITE_CYCLE_ACTIVE_rep14_i_ess\
        );

    \I__647\ : InMux
    port map (
            O => \N__4964\,
            I => \N__4961\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__4961\,
            I => \WRITE_CYCLE_ACTIVE_rep6_i_ess\
        );

    \I__645\ : IoInMux
    port map (
            O => \N__4958\,
            I => \N__4955\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__4955\,
            I => \N__4952\
        );

    \I__643\ : IoSpan4Mux
    port map (
            O => \N__4952\,
            I => \N__4949\
        );

    \I__642\ : Span4Mux_s2_v
    port map (
            O => \N__4949\,
            I => \N__4946\
        );

    \I__641\ : Span4Mux_v
    port map (
            O => \N__4946\,
            I => \N__4943\
        );

    \I__640\ : Odrv4
    port map (
            O => \N__4943\,
            I => \N_218_i\
        );

    \I__639\ : InMux
    port map (
            O => \N__4940\,
            I => \N__4937\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__4937\,
            I => \N__4934\
        );

    \I__637\ : Span4Mux_v
    port map (
            O => \N__4934\,
            I => \N__4931\
        );

    \I__636\ : Sp12to4
    port map (
            O => \N__4931\,
            I => \N__4928\
        );

    \I__635\ : Span12Mux_h
    port map (
            O => \N__4928\,
            I => \N__4925\
        );

    \I__634\ : Span12Mux_h
    port map (
            O => \N__4925\,
            I => \N__4922\
        );

    \I__633\ : Odrv12
    port map (
            O => \N__4922\,
            I => \D_UU_040_in_7\
        );

    \I__632\ : IoInMux
    port map (
            O => \N__4919\,
            I => \N__4916\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__4916\,
            I => \N__4913\
        );

    \I__630\ : IoSpan4Mux
    port map (
            O => \N__4913\,
            I => \N__4909\
        );

    \I__629\ : InMux
    port map (
            O => \N__4912\,
            I => \N__4906\
        );

    \I__628\ : Span4Mux_s2_h
    port map (
            O => \N__4909\,
            I => \N__4903\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__4906\,
            I => \N__4900\
        );

    \I__626\ : Span4Mux_h
    port map (
            O => \N__4903\,
            I => \N__4895\
        );

    \I__625\ : Span4Mux_v
    port map (
            O => \N__4900\,
            I => \N__4895\
        );

    \I__624\ : Span4Mux_h
    port map (
            O => \N__4895\,
            I => \N__4892\
        );

    \I__623\ : Sp12to4
    port map (
            O => \N__4892\,
            I => \N__4889\
        );

    \I__622\ : Span12Mux_h
    port map (
            O => \N__4889\,
            I => \N__4886\
        );

    \I__621\ : Odrv12
    port map (
            O => \N__4886\,
            I => \D_LM_040_in_7\
        );

    \I__620\ : IoInMux
    port map (
            O => \N__4883\,
            I => \N__4880\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__4880\,
            I => \N__4877\
        );

    \I__618\ : IoSpan4Mux
    port map (
            O => \N__4877\,
            I => \N__4874\
        );

    \I__617\ : Span4Mux_s2_v
    port map (
            O => \N__4874\,
            I => \N__4871\
        );

    \I__616\ : Span4Mux_v
    port map (
            O => \N__4871\,
            I => \N__4868\
        );

    \I__615\ : Odrv4
    port map (
            O => \N__4868\,
            I => \un1_D_UU_040_7\
        );

    \I__614\ : IoInMux
    port map (
            O => \N__4865\,
            I => \N__4862\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__4862\,
            I => \N__4859\
        );

    \I__612\ : Span4Mux_s3_v
    port map (
            O => \N__4859\,
            I => \N__4856\
        );

    \I__611\ : Span4Mux_h
    port map (
            O => \N__4856\,
            I => \N__4853\
        );

    \I__610\ : Odrv4
    port map (
            O => \N__4853\,
            I => \N_219_i\
        );

    \I__609\ : InMux
    port map (
            O => \N__4850\,
            I => \N__4847\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__4847\,
            I => \N__4844\
        );

    \I__607\ : Span4Mux_v
    port map (
            O => \N__4844\,
            I => \N__4841\
        );

    \I__606\ : Sp12to4
    port map (
            O => \N__4841\,
            I => \N__4838\
        );

    \I__605\ : Odrv12
    port map (
            O => \N__4838\,
            I => \D_LL_AMIGA_in_5\
        );

    \I__604\ : IoInMux
    port map (
            O => \N__4835\,
            I => \N__4832\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__4832\,
            I => \N__4829\
        );

    \I__602\ : Span4Mux_s1_h
    port map (
            O => \N__4829\,
            I => \N__4826\
        );

    \I__601\ : Span4Mux_h
    port map (
            O => \N__4826\,
            I => \N__4823\
        );

    \I__600\ : Sp12to4
    port map (
            O => \N__4823\,
            I => \N__4820\
        );

    \I__599\ : Span12Mux_s11_v
    port map (
            O => \N__4820\,
            I => \N__4817\
        );

    \I__598\ : Span12Mux_h
    port map (
            O => \N__4817\,
            I => \N__4814\
        );

    \I__597\ : Odrv12
    port map (
            O => \N__4814\,
            I => \un2_D_LL_AMIGA_5\
        );

    \I__596\ : InMux
    port map (
            O => \N__4811\,
            I => \N__4808\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__4808\,
            I => \N__4805\
        );

    \I__594\ : Odrv12
    port map (
            O => \N__4805\,
            I => \D_LM_AMIGA_in_1\
        );

    \I__593\ : InMux
    port map (
            O => \N__4802\,
            I => \N__4799\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__4799\,
            I => \WRITE_CYCLE_ACTIVE_rep1_i_ess\
        );

    \I__591\ : InMux
    port map (
            O => \N__4796\,
            I => \N__4793\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__4793\,
            I => \WRITE_CYCLE_ACTIVE_rep5_i_ess\
        );

    \I__589\ : IoInMux
    port map (
            O => \N__4790\,
            I => \N__4787\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__4787\,
            I => \N__4784\
        );

    \I__587\ : Span4Mux_s3_v
    port map (
            O => \N__4784\,
            I => \N__4781\
        );

    \I__586\ : Span4Mux_h
    port map (
            O => \N__4781\,
            I => \N__4778\
        );

    \I__585\ : Odrv4
    port map (
            O => \N__4778\,
            I => \N_215_i\
        );

    \I__584\ : IoInMux
    port map (
            O => \N__4775\,
            I => \N__4772\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__4772\,
            I => \N__4769\
        );

    \I__582\ : Odrv12
    port map (
            O => \N__4769\,
            I => \U111_CYCLE_SM_A_AMIGA_0_i_1\
        );

    \I__581\ : InMux
    port map (
            O => \N__4766\,
            I => \N__4763\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__4763\,
            I => \N__4760\
        );

    \I__579\ : Span4Mux_h
    port map (
            O => \N__4760\,
            I => \N__4757\
        );

    \I__578\ : Span4Mux_v
    port map (
            O => \N__4757\,
            I => \N__4754\
        );

    \I__577\ : Odrv4
    port map (
            O => \N__4754\,
            I => \A_040_c_0\
        );

    \I__576\ : IoInMux
    port map (
            O => \N__4751\,
            I => \N__4748\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__4748\,
            I => \N__4745\
        );

    \I__574\ : IoSpan4Mux
    port map (
            O => \N__4745\,
            I => \N__4742\
        );

    \I__573\ : Span4Mux_s2_v
    port map (
            O => \N__4742\,
            I => \N__4739\
        );

    \I__572\ : Span4Mux_v
    port map (
            O => \N__4739\,
            I => \N__4736\
        );

    \I__571\ : Odrv4
    port map (
            O => \N__4736\,
            I => \A_AMIGA_c_0\
        );

    \I__570\ : InMux
    port map (
            O => \N__4733\,
            I => \N__4730\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__4730\,
            I => \N__4727\
        );

    \I__568\ : Span4Mux_v
    port map (
            O => \N__4727\,
            I => \N__4724\
        );

    \I__567\ : Span4Mux_h
    port map (
            O => \N__4724\,
            I => \N__4721\
        );

    \I__566\ : Odrv4
    port map (
            O => \N__4721\,
            I => \D_LL_AMIGA_in_7\
        );

    \I__565\ : IoInMux
    port map (
            O => \N__4718\,
            I => \N__4715\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__4715\,
            I => \N__4712\
        );

    \I__563\ : Span4Mux_s2_h
    port map (
            O => \N__4712\,
            I => \N__4709\
        );

    \I__562\ : Span4Mux_v
    port map (
            O => \N__4709\,
            I => \N__4706\
        );

    \I__561\ : Sp12to4
    port map (
            O => \N__4706\,
            I => \N__4703\
        );

    \I__560\ : Span12Mux_h
    port map (
            O => \N__4703\,
            I => \N__4700\
        );

    \I__559\ : Span12Mux_h
    port map (
            O => \N__4700\,
            I => \N__4697\
        );

    \I__558\ : Odrv12
    port map (
            O => \N__4697\,
            I => \un2_D_LL_AMIGA_7\
        );

    \I__557\ : InMux
    port map (
            O => \N__4694\,
            I => \N__4690\
        );

    \I__556\ : IoInMux
    port map (
            O => \N__4693\,
            I => \N__4687\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__4690\,
            I => \N__4684\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__4687\,
            I => \N__4681\
        );

    \I__553\ : Span4Mux_v
    port map (
            O => \N__4684\,
            I => \N__4678\
        );

    \I__552\ : IoSpan4Mux
    port map (
            O => \N__4681\,
            I => \N__4675\
        );

    \I__551\ : Sp12to4
    port map (
            O => \N__4678\,
            I => \N__4672\
        );

    \I__550\ : Span4Mux_s2_h
    port map (
            O => \N__4675\,
            I => \N__4669\
        );

    \I__549\ : Span12Mux_h
    port map (
            O => \N__4672\,
            I => \N__4666\
        );

    \I__548\ : Sp12to4
    port map (
            O => \N__4669\,
            I => \N__4663\
        );

    \I__547\ : Span12Mux_v
    port map (
            O => \N__4666\,
            I => \N__4660\
        );

    \I__546\ : Span12Mux_h
    port map (
            O => \N__4663\,
            I => \N__4657\
        );

    \I__545\ : Span12Mux_h
    port map (
            O => \N__4660\,
            I => \N__4654\
        );

    \I__544\ : Span12Mux_h
    port map (
            O => \N__4657\,
            I => \N__4651\
        );

    \I__543\ : Odrv12
    port map (
            O => \N__4654\,
            I => \D_LL_040_in_2\
        );

    \I__542\ : Odrv12
    port map (
            O => \N__4651\,
            I => \D_LL_040_in_2\
        );

    \I__541\ : InMux
    port map (
            O => \N__4646\,
            I => \N__4643\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__4643\,
            I => \N__4640\
        );

    \I__539\ : Span12Mux_h
    port map (
            O => \N__4640\,
            I => \N__4637\
        );

    \I__538\ : Span12Mux_h
    port map (
            O => \N__4637\,
            I => \N__4634\
        );

    \I__537\ : Odrv12
    port map (
            O => \N__4634\,
            I => \D_UM_040_in_2\
        );

    \I__536\ : IoInMux
    port map (
            O => \N__4631\,
            I => \N__4628\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__4628\,
            I => \N__4625\
        );

    \I__534\ : Span4Mux_s1_h
    port map (
            O => \N__4625\,
            I => \N__4622\
        );

    \I__533\ : Span4Mux_h
    port map (
            O => \N__4622\,
            I => \N__4619\
        );

    \I__532\ : Span4Mux_v
    port map (
            O => \N__4619\,
            I => \N__4616\
        );

    \I__531\ : Odrv4
    port map (
            O => \N__4616\,
            I => \un1_D_UM_040_2\
        );

    \I__530\ : InMux
    port map (
            O => \N__4613\,
            I => \N__4610\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__4610\,
            I => \N__4607\
        );

    \I__528\ : Odrv4
    port map (
            O => \N__4607\,
            I => \WRITE_CYCLE_ACTIVE_rep8_i_ess\
        );

    \I__527\ : InMux
    port map (
            O => \N__4604\,
            I => \N__4601\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__4601\,
            I => \N__4598\
        );

    \I__525\ : Odrv4
    port map (
            O => \N__4598\,
            I => \WRITE_CYCLE_ACTIVE_rep10_i_ess\
        );

    \I__524\ : InMux
    port map (
            O => \N__4595\,
            I => \N__4592\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__4592\,
            I => \WRITE_CYCLE_ACTIVE_rep17_i_ess\
        );

    \I__522\ : InMux
    port map (
            O => \N__4589\,
            I => \N__4586\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__4586\,
            I => \WRITE_CYCLE_ACTIVE_rep19_i_ess\
        );

    \I__520\ : InMux
    port map (
            O => \N__4583\,
            I => \N__4580\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__4580\,
            I => \WRITE_CYCLE_ACTIVE_rep18_i_ess\
        );

    \I__518\ : InMux
    port map (
            O => \N__4577\,
            I => \N__4574\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__4574\,
            I => \WRITE_CYCLE_ACTIVE_rep20_i_ess\
        );

    \I__516\ : InMux
    port map (
            O => \N__4571\,
            I => \N__4568\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__4568\,
            I => \WRITE_CYCLE_ACTIVE_rep21_i_ess\
        );

    \I__514\ : InMux
    port map (
            O => \N__4565\,
            I => \N__4562\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__4562\,
            I => \WRITE_CYCLE_ACTIVE_rep22_i_ess\
        );

    \I__512\ : InMux
    port map (
            O => \N__4559\,
            I => \N__4556\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__4556\,
            I => \WRITE_CYCLE_ACTIVE_rep9_i_ess\
        );

    \I__510\ : InMux
    port map (
            O => \N__4553\,
            I => \N__4550\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__4550\,
            I => \WRITE_CYCLE_ACTIVE_rep23_i_ess\
        );

    \I__508\ : InMux
    port map (
            O => \N__4547\,
            I => \N__4544\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__4544\,
            I => \WRITE_CYCLE_ACTIVE_rep11_i_ess\
        );

    \I__506\ : InMux
    port map (
            O => \N__4541\,
            I => \N__4538\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4538\,
            I => \N__4535\
        );

    \I__504\ : Odrv4
    port map (
            O => \N__4535\,
            I => \WRITE_CYCLE_ACTIVE_rep24_i_ess\
        );

    \I__503\ : InMux
    port map (
            O => \N__4532\,
            I => \N__4529\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__4529\,
            I => \WRITE_CYCLE_ACTIVE_rep25_i_ess\
        );

    \I__501\ : InMux
    port map (
            O => \N__4526\,
            I => \N__4523\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4523\,
            I => \WRITE_CYCLE_ACTIVE_rep28_i_ess\
        );

    \I__499\ : InMux
    port map (
            O => \N__4520\,
            I => \N__4517\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__4517\,
            I => \N__4514\
        );

    \I__497\ : Odrv4
    port map (
            O => \N__4514\,
            I => \WRITE_CYCLE_ACTIVE_rep27_i_ess\
        );

    \I__496\ : InMux
    port map (
            O => \N__4511\,
            I => \N__4508\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__4508\,
            I => \N__4505\
        );

    \I__494\ : Odrv12
    port map (
            O => \N__4505\,
            I => \WRITE_CYCLE_ACTIVE_rep26_i_ess\
        );

    \I__493\ : InMux
    port map (
            O => \N__4502\,
            I => \N__4499\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__4499\,
            I => \WRITE_CYCLE_ACTIVE_rep30_i_ess\
        );

    \I__491\ : InMux
    port map (
            O => \N__4496\,
            I => \N__4493\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__4493\,
            I => \WRITE_CYCLE_ACTIVE_rep16_i_ess\
        );

    \I__489\ : InMux
    port map (
            O => \N__4490\,
            I => \N__4487\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__4487\,
            I => \WRITE_CYCLE_ACTIVE_rep29_i_ess\
        );

    \I__487\ : InMux
    port map (
            O => \N__4484\,
            I => \N__4481\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__4481\,
            I => \WRITE_CYCLE_ACTIVE_i_ess\
        );

    \I__485\ : IoInMux
    port map (
            O => \N__4478\,
            I => \N__4475\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__4475\,
            I => \N__4472\
        );

    \I__483\ : IoSpan4Mux
    port map (
            O => \N__4472\,
            I => \N__4469\
        );

    \I__482\ : Span4Mux_s3_h
    port map (
            O => \N__4469\,
            I => \N__4466\
        );

    \I__481\ : Odrv4
    port map (
            O => \N__4466\,
            I => \N_235_i\
        );

    \I__480\ : IoInMux
    port map (
            O => \N__4463\,
            I => \N__4460\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4460\,
            I => \N__4457\
        );

    \I__478\ : IoSpan4Mux
    port map (
            O => \N__4457\,
            I => \N__4454\
        );

    \I__477\ : Span4Mux_s3_h
    port map (
            O => \N__4454\,
            I => \N__4451\
        );

    \I__476\ : Odrv4
    port map (
            O => \N__4451\,
            I => \N_213_i\
        );

    \I__475\ : IoInMux
    port map (
            O => \N__4448\,
            I => \N__4445\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__4445\,
            I => \N__4442\
        );

    \I__473\ : Span4Mux_s0_h
    port map (
            O => \N__4442\,
            I => \N__4439\
        );

    \I__472\ : Span4Mux_h
    port map (
            O => \N__4439\,
            I => \N__4436\
        );

    \I__471\ : Odrv4
    port map (
            O => \N__4436\,
            I => \N_223_i\
        );

    \I__470\ : IoInMux
    port map (
            O => \N__4433\,
            I => \N__4430\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__4430\,
            I => \N__4427\
        );

    \I__468\ : IoSpan4Mux
    port map (
            O => \N__4427\,
            I => \N__4424\
        );

    \I__467\ : Span4Mux_s3_h
    port map (
            O => \N__4424\,
            I => \N__4421\
        );

    \I__466\ : Odrv4
    port map (
            O => \N__4421\,
            I => \N_224_i\
        );

    \I__465\ : IoInMux
    port map (
            O => \N__4418\,
            I => \N__4415\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__4415\,
            I => \N__4412\
        );

    \I__463\ : IoSpan4Mux
    port map (
            O => \N__4412\,
            I => \N__4409\
        );

    \I__462\ : Span4Mux_s3_v
    port map (
            O => \N__4409\,
            I => \N__4406\
        );

    \I__461\ : Span4Mux_v
    port map (
            O => \N__4406\,
            I => \N__4403\
        );

    \I__460\ : Odrv4
    port map (
            O => \N__4403\,
            I => \N_217_i\
        );

    \I__459\ : IoInMux
    port map (
            O => \N__4400\,
            I => \N__4397\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__4397\,
            I => \N__4394\
        );

    \I__457\ : Span4Mux_s0_h
    port map (
            O => \N__4394\,
            I => \N__4391\
        );

    \I__456\ : Span4Mux_h
    port map (
            O => \N__4391\,
            I => \N__4388\
        );

    \I__455\ : Odrv4
    port map (
            O => \N__4388\,
            I => \N_227_i\
        );

    \I__454\ : IoInMux
    port map (
            O => \N__4385\,
            I => \N__4382\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__4382\,
            I => \N__4379\
        );

    \I__452\ : IoSpan4Mux
    port map (
            O => \N__4379\,
            I => \N__4376\
        );

    \I__451\ : Span4Mux_s0_h
    port map (
            O => \N__4376\,
            I => \N__4373\
        );

    \I__450\ : Span4Mux_h
    port map (
            O => \N__4373\,
            I => \N__4370\
        );

    \I__449\ : Odrv4
    port map (
            O => \N__4370\,
            I => \N_226_i\
        );

    \I__448\ : IoInMux
    port map (
            O => \N__4367\,
            I => \N__4364\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__4364\,
            I => \N__4361\
        );

    \I__446\ : IoSpan4Mux
    port map (
            O => \N__4361\,
            I => \N__4358\
        );

    \I__445\ : Span4Mux_s3_h
    port map (
            O => \N__4358\,
            I => \N__4355\
        );

    \I__444\ : Odrv4
    port map (
            O => \N__4355\,
            I => \N_236_i\
        );

    \I__443\ : IoInMux
    port map (
            O => \N__4352\,
            I => \N__4349\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__4349\,
            I => \N__4346\
        );

    \I__441\ : IoSpan4Mux
    port map (
            O => \N__4346\,
            I => \N__4343\
        );

    \I__440\ : Span4Mux_s1_h
    port map (
            O => \N__4343\,
            I => \N__4340\
        );

    \I__439\ : Span4Mux_h
    port map (
            O => \N__4340\,
            I => \N__4337\
        );

    \I__438\ : Odrv4
    port map (
            O => \N__4337\,
            I => \N_239_i\
        );

    \I__437\ : IoInMux
    port map (
            O => \N__4334\,
            I => \N__4331\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__4331\,
            I => \N__4328\
        );

    \I__435\ : IoSpan4Mux
    port map (
            O => \N__4328\,
            I => \N__4325\
        );

    \I__434\ : Span4Mux_s1_h
    port map (
            O => \N__4325\,
            I => \N__4322\
        );

    \I__433\ : Span4Mux_h
    port map (
            O => \N__4322\,
            I => \N__4319\
        );

    \I__432\ : Odrv4
    port map (
            O => \N__4319\,
            I => \N_238_i\
        );

    \I__431\ : IoInMux
    port map (
            O => \N__4316\,
            I => \N__4313\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__4313\,
            I => \N__4310\
        );

    \I__429\ : Odrv12
    port map (
            O => \N__4310\,
            I => \RESETn_c_i\
        );

    \I__428\ : IoInMux
    port map (
            O => \N__4307\,
            I => \N__4304\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__4304\,
            I => \N__4301\
        );

    \I__426\ : Odrv12
    port map (
            O => \N__4301\,
            I => \N_231_i\
        );

    \I__425\ : IoInMux
    port map (
            O => \N__4298\,
            I => \N__4295\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__4295\,
            I => \N__4292\
        );

    \I__423\ : Odrv12
    port map (
            O => \N__4292\,
            I => \N_220_i\
        );

    \I__422\ : IoInMux
    port map (
            O => \N__4289\,
            I => \N__4286\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__4286\,
            I => \N__4283\
        );

    \I__420\ : Odrv12
    port map (
            O => \N__4283\,
            I => \N_230_i\
        );

    \I__419\ : IoInMux
    port map (
            O => \N__4280\,
            I => \N__4277\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__4277\,
            I => \N__4274\
        );

    \I__417\ : Span12Mux_s4_h
    port map (
            O => \N__4274\,
            I => \N__4271\
        );

    \I__416\ : Odrv12
    port map (
            O => \N__4271\,
            I => \N_232_i\
        );

    \I__415\ : IoInMux
    port map (
            O => \N__4268\,
            I => \N__4265\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__4265\,
            I => \N__4262\
        );

    \I__413\ : IoSpan4Mux
    port map (
            O => \N__4262\,
            I => \N__4259\
        );

    \I__412\ : Span4Mux_s3_h
    port map (
            O => \N__4259\,
            I => \N__4256\
        );

    \I__411\ : Odrv4
    port map (
            O => \N__4256\,
            I => \N_222_i\
        );

    \I__410\ : IoInMux
    port map (
            O => \N__4253\,
            I => \N__4250\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__4250\,
            I => \N__4247\
        );

    \I__408\ : IoSpan4Mux
    port map (
            O => \N__4247\,
            I => \N__4244\
        );

    \I__407\ : Span4Mux_s3_h
    port map (
            O => \N__4244\,
            I => \N__4241\
        );

    \I__406\ : Odrv4
    port map (
            O => \N__4241\,
            I => \N_221_i\
        );

    \I__405\ : IoInMux
    port map (
            O => \N__4238\,
            I => \N__4235\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__4235\,
            I => \N__4232\
        );

    \I__403\ : IoSpan4Mux
    port map (
            O => \N__4232\,
            I => \N__4229\
        );

    \I__402\ : Span4Mux_s2_h
    port map (
            O => \N__4229\,
            I => \N__4226\
        );

    \I__401\ : Odrv4
    port map (
            O => \N__4226\,
            I => \N_233_i\
        );

    \I__400\ : IoInMux
    port map (
            O => \N__4223\,
            I => \N__4220\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__4220\,
            I => \N__4217\
        );

    \I__398\ : IoSpan4Mux
    port map (
            O => \N__4217\,
            I => \N__4214\
        );

    \I__397\ : Span4Mux_s3_h
    port map (
            O => \N__4214\,
            I => \N__4211\
        );

    \I__396\ : Odrv4
    port map (
            O => \N__4211\,
            I => \N_234_i\
        );

    \I__395\ : IoInMux
    port map (
            O => \N__4208\,
            I => \N__4205\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__4205\,
            I => \N__4202\
        );

    \I__393\ : Span4Mux_s0_v
    port map (
            O => \N__4202\,
            I => \N__4199\
        );

    \I__392\ : Sp12to4
    port map (
            O => \N__4199\,
            I => \N__4196\
        );

    \I__391\ : Span12Mux_h
    port map (
            O => \N__4196\,
            I => \N__4193\
        );

    \I__390\ : Span12Mux_v
    port map (
            O => \N__4193\,
            I => \N__4190\
        );

    \I__389\ : Span12Mux_v
    port map (
            O => \N__4190\,
            I => \N__4187\
        );

    \I__388\ : Odrv12
    port map (
            O => \N__4187\,
            I => \TAn_in\
        );

    \I__387\ : IoInMux
    port map (
            O => \N__4184\,
            I => \N__4181\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__4181\,
            I => \N__4178\
        );

    \I__385\ : Span12Mux_s4_h
    port map (
            O => \N__4178\,
            I => \N__4175\
        );

    \I__384\ : Odrv12
    port map (
            O => \N__4175\,
            I => \N_237_i\
        );

    \I__383\ : IoInMux
    port map (
            O => \N__4172\,
            I => \N__4169\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__4169\,
            I => \N__4166\
        );

    \I__381\ : IoSpan4Mux
    port map (
            O => \N__4166\,
            I => \N__4163\
        );

    \I__380\ : Span4Mux_s1_h
    port map (
            O => \N__4163\,
            I => \N__4160\
        );

    \I__379\ : Odrv4
    port map (
            O => \N__4160\,
            I => \N_240_i\
        );

    \I__378\ : IoInMux
    port map (
            O => \N__4157\,
            I => \N__4154\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__4154\,
            I => \N__4151\
        );

    \I__376\ : Span4Mux_s0_h
    port map (
            O => \N__4151\,
            I => \N__4148\
        );

    \I__375\ : Span4Mux_h
    port map (
            O => \N__4148\,
            I => \N__4145\
        );

    \I__374\ : Odrv4
    port map (
            O => \N__4145\,
            I => \N_242_i\
        );

    \I__373\ : IoInMux
    port map (
            O => \N__4142\,
            I => \N__4139\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__4139\,
            I => \N__4136\
        );

    \I__371\ : Span4Mux_s0_h
    port map (
            O => \N__4136\,
            I => \N__4133\
        );

    \I__370\ : Span4Mux_h
    port map (
            O => \N__4133\,
            I => \N__4130\
        );

    \I__369\ : Odrv4
    port map (
            O => \N__4130\,
            I => \N_228_i\
        );

    \I__368\ : IoInMux
    port map (
            O => \N__4127\,
            I => \N__4124\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__4124\,
            I => \N__4121\
        );

    \I__366\ : IoSpan4Mux
    port map (
            O => \N__4121\,
            I => \N__4118\
        );

    \I__365\ : Span4Mux_s3_h
    port map (
            O => \N__4118\,
            I => \N__4115\
        );

    \I__364\ : Odrv4
    port map (
            O => \N__4115\,
            I => \N_241_i\
        );

    \I__363\ : IoInMux
    port map (
            O => \N__4112\,
            I => \N__4109\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__4109\,
            I => \N__4106\
        );

    \I__361\ : Span12Mux_s4_h
    port map (
            O => \N__4106\,
            I => \N__4103\
        );

    \I__360\ : Odrv12
    port map (
            O => \N__4103\,
            I => \N_243_i\
        );

    \I__359\ : IoInMux
    port map (
            O => \N__4100\,
            I => \N__4097\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__4097\,
            I => \N__4094\
        );

    \I__357\ : Span4Mux_s0_h
    port map (
            O => \N__4094\,
            I => \N__4091\
        );

    \I__356\ : Span4Mux_h
    port map (
            O => \N__4091\,
            I => \N__4088\
        );

    \I__355\ : Odrv4
    port map (
            O => \N__4088\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_0\
        );

    \I__354\ : IoInMux
    port map (
            O => \N__4085\,
            I => \N__4082\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__4082\,
            I => \N__4079\
        );

    \I__352\ : Odrv12
    port map (
            O => \N__4079\,
            I => \N_229_i\
        );

    \I__351\ : IoInMux
    port map (
            O => \N__4076\,
            I => \N__4073\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__4073\,
            I => \N__4070\
        );

    \I__349\ : IoSpan4Mux
    port map (
            O => \N__4070\,
            I => \N__4067\
        );

    \I__348\ : Span4Mux_s3_h
    port map (
            O => \N__4067\,
            I => \N__4064\
        );

    \I__347\ : Sp12to4
    port map (
            O => \N__4064\,
            I => \N__4061\
        );

    \I__346\ : Span12Mux_s8_h
    port map (
            O => \N__4061\,
            I => \N__4058\
        );

    \I__345\ : Span12Mux_v
    port map (
            O => \N__4058\,
            I => \N__4055\
        );

    \I__344\ : Span12Mux_v
    port map (
            O => \N__4055\,
            I => \N__4052\
        );

    \I__343\ : Span12Mux_h
    port map (
            O => \N__4052\,
            I => \N__4049\
        );

    \I__342\ : Odrv12
    port map (
            O => \N__4049\,
            I => \TCIn_c\
        );

    \INVU111_CYCLE_SM.TSnC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.TSnC_net\,
            I => \N__10601\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4316\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIICIM_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4100\,
            GLOBALBUFFEROUTPUT => \U111_CYCLE_SM.CYCLE_STATE_0_g_0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \D_LL_AMIGA_iobuf_RNO_1_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4532\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_237_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_AMIGA_iobuf_RNO_4_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4526\,
            lcout => \N_240_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_AMIGA_iobuf_RNO_6_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4502\,
            lcout => \N_242_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_AMIGA_iobuf_RNO_0_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4496\,
            lcout => \N_228_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_AMIGA_iobuf_RNO_5_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4490\,
            lcout => \N_241_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_AMIGA_iobuf_RNO_7_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4484\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_243_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIICIM_0_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10319\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6779\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_AMIGA_iobuf_RNO_1_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4595\,
            lcout => \N_229_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6709\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_AMIGA_iobuf_RNO_3_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4589\,
            lcout => \N_231_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_0_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4613\,
            lcout => \N_220_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_AMIGA_iobuf_RNO_2_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4583\,
            lcout => \N_230_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_AMIGA_iobuf_RNO_4_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4577\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_232_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_2_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4604\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_222_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_1_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4559\,
            lcout => \N_221_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_AMIGA_iobuf_RNO_5_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4571\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_233_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_AMIGA_iobuf_RNO_6_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4565\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_234_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_AMIGA_iobuf_RNO_7_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4553\,
            lcout => \N_235_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_AMIGA_iobuf_RNO_1_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4802\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_213_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_3_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4547\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_223_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_4_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4985\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_224_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_AMIGA_iobuf_RNO_5_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4796\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_217_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_7_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5204\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_227_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_AMIGA_iobuf_RNO_6_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4973\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_226_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_AMIGA_iobuf_RNO_0_LC_2_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4541\,
            lcout => \N_236_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_AMIGA_iobuf_RNO_3_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4520\,
            lcout => \N_239_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_AMIGA_iobuf_RNO_2_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4511\,
            lcout => \N_238_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep24_i_ess_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__12545\,
            in1 => \N__11117\,
            in2 => \N__12184\,
            in3 => \N__11231\,
            lcout => \WRITE_CYCLE_ACTIVE_rep24_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10625\,
            ce => \N__10422\,
            sr => \N__10283\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep25_i_ess_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__11232\,
            in1 => \N__11079\,
            in2 => \N__12185\,
            in3 => \N__12546\,
            lcout => \WRITE_CYCLE_ACTIVE_rep25_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10625\,
            ce => \N__10422\,
            sr => \N__10283\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep28_i_ess_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__12547\,
            in1 => \N__12183\,
            in2 => \N__11113\,
            in3 => \N__11233\,
            lcout => \WRITE_CYCLE_ACTIVE_rep28_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10625\,
            ce => \N__10422\,
            sr => \N__10283\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep27_i_ess_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__12168\,
            in1 => \N__11116\,
            in2 => \N__12722\,
            in3 => \N__11430\,
            lcout => \WRITE_CYCLE_ACTIVE_rep27_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10622\,
            ce => \N__10419\,
            sr => \N__10281\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep26_i_ess_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__11115\,
            in1 => \N__12167\,
            in2 => \N__11509\,
            in3 => \N__12713\,
            lcout => \WRITE_CYCLE_ACTIVE_rep26_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10621\,
            ce => \N__10417\,
            sr => \N__10279\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep30_i_ess_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__12166\,
            in1 => \N__11114\,
            in2 => \N__12721\,
            in3 => \N__11434\,
            lcout => \WRITE_CYCLE_ACTIVE_rep30_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10619\,
            ce => \N__10416\,
            sr => \N__10277\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep16_i_ess_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__11093\,
            in1 => \N__12165\,
            in2 => \N__11510\,
            in3 => \N__12717\,
            lcout => \WRITE_CYCLE_ACTIVE_rep16_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10617\,
            ce => \N__10414\,
            sr => \N__10274\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep29_i_ess_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__11092\,
            in1 => \N__12144\,
            in2 => \N__11564\,
            in3 => \N__12689\,
            lcout => \WRITE_CYCLE_ACTIVE_rep29_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10616\,
            ce => \N__10412\,
            sr => \N__10272\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_i_ess_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__11091\,
            in1 => \N__11514\,
            in2 => \N__12164\,
            in3 => \N__12679\,
            lcout => \WRITE_CYCLE_ACTIVE_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10614\,
            ce => \N__10409\,
            sr => \N__10270\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep17_i_ess_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__11090\,
            in1 => \N__12678\,
            in2 => \N__12163\,
            in3 => \N__11515\,
            lcout => \WRITE_CYCLE_ACTIVE_rep17_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10610\,
            ce => \N__10407\,
            sr => \N__10269\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep19_i_ess_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__11033\,
            in1 => \N__12137\,
            in2 => \N__12720\,
            in3 => \N__11516\,
            lcout => \WRITE_CYCLE_ACTIVE_rep19_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10609\,
            ce => \N__10406\,
            sr => \N__10271\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep18_i_ess_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__11032\,
            in1 => \N__12620\,
            in2 => \N__11606\,
            in3 => \N__12106\,
            lcout => \WRITE_CYCLE_ACTIVE_rep18_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10607\,
            ce => \N__10408\,
            sr => \N__10273\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep20_i_ess_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__12099\,
            in1 => \N__11030\,
            in2 => \N__12677\,
            in3 => \N__11570\,
            lcout => \WRITE_CYCLE_ACTIVE_rep20_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10605\,
            ce => \N__10410\,
            sr => \N__10275\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep21_i_ess_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__11057\,
            in1 => \N__12096\,
            in2 => \N__12544\,
            in3 => \N__11571\,
            lcout => \WRITE_CYCLE_ACTIVE_rep21_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10603\,
            ce => \N__10415\,
            sr => \N__10280\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep22_i_ess_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__12467\,
            in1 => \N__12097\,
            in2 => \N__11106\,
            in3 => \N__11572\,
            lcout => \WRITE_CYCLE_ACTIVE_rep22_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10603\,
            ce => \N__10415\,
            sr => \N__10280\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep9_i_ess_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__12468\,
            in1 => \N__12098\,
            in2 => \N__11107\,
            in3 => \N__11573\,
            lcout => \WRITE_CYCLE_ACTIVE_rep9_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10603\,
            ce => \N__10415\,
            sr => \N__10280\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep23_i_ess_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__12640\,
            in1 => \N__11065\,
            in2 => \N__12095\,
            in3 => \N__11608\,
            lcout => \WRITE_CYCLE_ACTIVE_rep23_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10600\,
            ce => \N__10418\,
            sr => \N__10282\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep11_i_ess_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__11108\,
            in1 => \N__12641\,
            in2 => \N__11629\,
            in3 => \N__12034\,
            lcout => \WRITE_CYCLE_ACTIVE_rep11_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10595\,
            ce => \N__10420\,
            sr => \N__10284\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep1_i_ess_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__11109\,
            in1 => \N__12642\,
            in2 => \N__11630\,
            in3 => \N__12035\,
            lcout => \WRITE_CYCLE_ACTIVE_rep1_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10595\,
            ce => \N__10420\,
            sr => \N__10284\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep5_i_ess_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__11112\,
            in1 => \N__12033\,
            in2 => \N__12695\,
            in3 => \N__11617\,
            lcout => \WRITE_CYCLE_ACTIVE_rep5_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10588\,
            ce => \N__10421\,
            sr => \N__10285\
        );

    \D_UU_AMIGA_iobuf_RNO_3_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5195\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_215_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5818\,
            in2 => \_gnd_net_\,
            in3 => \N__6812\,
            lcout => \U111_CYCLE_SM_A_AMIGA_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__4766\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6811\,
            lcout => \A_AMIGA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_3_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8958\,
            in1 => \N__7145\,
            in2 => \_gnd_net_\,
            in3 => \N__4733\,
            lcout => \un2_D_LL_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8959\,
            in1 => \N__4694\,
            in2 => \_gnd_net_\,
            in3 => \N__4646\,
            lcout => \un1_D_UM_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep8_i_ess_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__11565\,
            in1 => \N__11031\,
            in2 => \N__12136\,
            in3 => \N__12670\,
            lcout => \WRITE_CYCLE_ACTIVE_rep8_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10606\,
            ce => \N__10411\,
            sr => \N__10276\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep10_i_ess_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__11566\,
            in1 => \N__11029\,
            in2 => \N__12019\,
            in3 => \N__12669\,
            lcout => \WRITE_CYCLE_ACTIVE_rep10_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10604\,
            ce => \N__10413\,
            sr => \N__10278\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5015\,
            in1 => \N__6993\,
            in2 => \_gnd_net_\,
            in3 => \N__8963\,
            lcout => \un2_D_LM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep12_i_ess_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__11064\,
            in1 => \N__11607\,
            in2 => \N__12709\,
            in3 => \N__12032\,
            lcout => \WRITE_CYCLE_ACTIVE_rep12_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10589\,
            ce => \N__10423\,
            sr => \N__10286\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep6_i_ess_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__11958\,
            in1 => \N__11111\,
            in2 => \N__12694\,
            in3 => \N__11616\,
            lcout => \WRITE_CYCLE_ACTIVE_rep6_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10584\,
            ce => \N__10424\,
            sr => \N__10288\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep14_i_ess_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__11957\,
            in1 => \N__11110\,
            in2 => \N__12693\,
            in3 => \N__11615\,
            lcout => \WRITE_CYCLE_ACTIVE_rep14_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10584\,
            ce => \N__10424\,
            sr => \N__10288\
        );

    \D_UU_AMIGA_iobuf_RNO_6_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4964\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_218_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8964\,
            in1 => \N__4940\,
            in2 => \_gnd_net_\,
            in3 => \N__4912\,
            lcout => \un1_D_UU_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_AMIGA_iobuf_RNO_7_LC_3_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5186\,
            lcout => \N_219_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4850\,
            in1 => \N__7214\,
            in2 => \_gnd_net_\,
            in3 => \N__8980\,
            lcout => \un2_D_LL_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9007\,
            in1 => \N__5987\,
            in2 => \_gnd_net_\,
            in3 => \N__4811\,
            lcout => \un2_D_LM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep0_i_ess_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__11619\,
            in1 => \N__11085\,
            in2 => \N__11990\,
            in3 => \N__12603\,
            lcout => \WRITE_CYCLE_ACTIVE_rep0_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10579\,
            ce => \N__10425\,
            sr => \N__10294\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep15_i_ess_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__11620\,
            in1 => \N__11086\,
            in2 => \N__11991\,
            in3 => \N__12604\,
            lcout => \WRITE_CYCLE_ACTIVE_rep15_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10579\,
            ce => \N__10425\,
            sr => \N__10294\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep3_i_ess_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__12699\,
            in1 => \N__11087\,
            in2 => \N__11988\,
            in3 => \N__11631\,
            lcout => \WRITE_CYCLE_ACTIVE_rep3_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10575\,
            ce => \N__10427\,
            sr => \N__10297\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep7_i_ess_LC_5_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__11089\,
            in1 => \N__11633\,
            in2 => \N__12719\,
            in3 => \N__11905\,
            lcout => \WRITE_CYCLE_ACTIVE_rep7_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10575\,
            ce => \N__10427\,
            sr => \N__10297\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep4_i_ess_LC_5_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__12700\,
            in1 => \N__11088\,
            in2 => \N__11989\,
            in3 => \N__11632\,
            lcout => \WRITE_CYCLE_ACTIVE_rep4_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10575\,
            ce => \N__10427\,
            sr => \N__10297\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5177\,
            in1 => \N__7783\,
            in2 => \_gnd_net_\,
            in3 => \N__8973\,
            lcout => \un2_D_LM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5141\,
            in1 => \N__8602\,
            in2 => \_gnd_net_\,
            in3 => \N__9005\,
            lcout => \un2_D_LM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_AMIGA_iobuf_RNO_2_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5336\,
            lcout => \N_214_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_6_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9020\,
            in1 => \N__5084\,
            in2 => \_gnd_net_\,
            in3 => \N__5063\,
            lcout => \un1_D_UU_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_AMIGA_iobuf_RNO_0_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5381\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_212_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_AMIGA_iobuf_RNO_4_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5357\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_216_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep2_i_ess_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__11505\,
            in1 => \N__11016\,
            in2 => \N__12031\,
            in3 => \N__12528\,
            lcout => \WRITE_CYCLE_ACTIVE_rep2_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10573\,
            ce => \N__10426\,
            sr => \N__10295\
        );

    \D_UM_AMIGA_iobuf_RNO_5_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5234\,
            lcout => \N_225_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \BUFENn_obuf_RNO_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11563\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \LBENn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9004\,
            in1 => \N__5300\,
            in2 => \_gnd_net_\,
            in3 => \N__7289\,
            lcout => \un2_D_LL_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8969\,
            in1 => \N__6926\,
            in2 => \_gnd_net_\,
            in3 => \N__5261\,
            lcout => \un2_D_LM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep13_i_ess_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__11015\,
            in1 => \N__11875\,
            in2 => \N__11618\,
            in3 => \N__12452\,
            lcout => \WRITE_CYCLE_ACTIVE_rep13_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10568\,
            ce => \N__10428\,
            sr => \N__10298\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5765\,
            in1 => \N__5737\,
            in2 => \_gnd_net_\,
            in3 => \N__9003\,
            lcout => \un1_D_UU_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7403\,
            in1 => \N__5681\,
            in2 => \_gnd_net_\,
            in3 => \N__8919\,
            lcout => \un2_D_LL_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8890\,
            in1 => \N__7073\,
            in2 => \_gnd_net_\,
            in3 => \N__5642\,
            lcout => \un2_D_LM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_10_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5603\,
            in1 => \N__7702\,
            in2 => \_gnd_net_\,
            in3 => \N__8979\,
            lcout => \un2_D_LL_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_10_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7636\,
            in1 => \N__5561\,
            in2 => \_gnd_net_\,
            in3 => \N__8965\,
            lcout => \un2_D_LL_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5528\,
            in1 => \N__8552\,
            in2 => \_gnd_net_\,
            in3 => \N__8993\,
            lcout => \un2_D_LM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LBENn_c_sbtinv_LC_11_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11216\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \LBENn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8935\,
            in1 => \N__5441\,
            in2 => \_gnd_net_\,
            in3 => \N__6617\,
            lcout => \un2_D_LL_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7504\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5825\,
            lcout => \U111_CYCLE_SM.FLIP_WORD_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TSn_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__6723\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5785\,
            lcout => \TSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TSnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001110111011"
        )
    port map (
            in0 => \N__5786\,
            in1 => \N__6791\,
            in2 => \N__5834\,
            in3 => \N__5855\,
            lcout => \U111_CYCLE_SM.TS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10596\,
            ce => 'H',
            sr => \N__10289\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__6230\,
            in1 => \N__6161\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_srsts_i_o2_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_5_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__6732\,
            in1 => \N__5848\,
            in2 => \N__5774\,
            in3 => \N__6061\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10591\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_3_0_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__6247\,
            in1 => \N__6428\,
            in2 => \_gnd_net_\,
            in3 => \N__6056\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.N_148_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100000000"
        )
    port map (
            in0 => \N__6758\,
            in1 => \N__5869\,
            in2 => \N__5771\,
            in3 => \N__6710\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_srsts_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_0_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100011111"
        )
    port map (
            in0 => \N__6029\,
            in1 => \N__6192\,
            in2 => \N__5768\,
            in3 => \N__6449\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10586\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIDUAQ_0_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__11083\,
            in1 => \N__12134\,
            in2 => \N__11408\,
            in3 => \N__6757\,
            lcout => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN6_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__12135\,
            in1 => \N__11084\,
            in2 => \_gnd_net_\,
            in3 => \N__11308\,
            lcout => \U111_CYCLE_SM.TS_ENZ0Z6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.BURST_COUNT_0_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011000"
        )
    port map (
            in0 => \N__6316\,
            in1 => \N__6443\,
            in2 => \N__6362\,
            in3 => \N__6395\,
            lcout => \U111_CYCLE_SM.BURST_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10580\,
            ce => 'H',
            sr => \N__10290\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_1_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5986\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10570\,
            ce => \N__7905\,
            sr => \N__7871\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNIUR6Q_1_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5979\,
            in1 => \N__5942\,
            in2 => \_gnd_net_\,
            in3 => \N__8450\,
            lcout => \un1_D_UU_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8915\,
            in1 => \N__7331\,
            in2 => \_gnd_net_\,
            in3 => \N__5912\,
            lcout => \un2_D_LL_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_2_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__6265\,
            in1 => \N__6182\,
            in2 => \_gnd_net_\,
            in3 => \N__6055\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.N_158_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_0_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__5873\,
            in1 => \N__6771\,
            in2 => \N__5858\,
            in3 => \N__6645\,
            lcout => \U111_CYCLE_SM.N_130_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_4_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6847\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6717\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10590\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_1_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__6846\,
            in1 => \N__7471\,
            in2 => \N__5849\,
            in3 => \N__6441\,
            lcout => \U111_CYCLE_SM.TS_EN_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIC4111_3_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6848\,
            in2 => \_gnd_net_\,
            in3 => \N__6390\,
            lcout => \U111_CYCLE_SM.un1_CYCLE_STATE_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__6167\,
            in1 => \N__6266\,
            in2 => \_gnd_net_\,
            in3 => \N__6060\,
            lcout => \U111_CYCLE_SM.N_160\,
            ltout => \U111_CYCLE_SM.N_160_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_1_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010000000"
        )
    port map (
            in0 => \N__6718\,
            in1 => \N__6439\,
            in2 => \N__6119\,
            in3 => \N__6391\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10585\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_3_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6719\,
            in1 => \N__7448\,
            in2 => \_gnd_net_\,
            in3 => \N__6320\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10585\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.BURST_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__6115\,
            in1 => \N__6440\,
            in2 => \N__6092\,
            in3 => \N__6392\,
            lcout => \U111_CYCLE_SM.BURSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10582\,
            ce => 'H',
            sr => \N__10287\
        );

    \U111_CYCLE_SM.LW_TRANS_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__6393\,
            in1 => \N__6116\,
            in2 => \N__7538\,
            in3 => \N__6091\,
            lcout => \U111_CYCLE_SM.LW_TRANSZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10582\,
            ce => 'H',
            sr => \N__10287\
        );

    \U111_CYCLE_SM.TA_DIS_RNO_0_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7516\,
            in2 => \_gnd_net_\,
            in3 => \N__7533\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.PORT_MISMATCH_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_DIS_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__7822\,
            in1 => \N__6850\,
            in2 => \N__6065\,
            in3 => \N__7472\,
            lcout => \U111_CYCLE_SM.TA_DISZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10582\,
            ce => 'H',
            sr => \N__10287\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6062\,
            in2 => \_gnd_net_\,
            in3 => \N__6646\,
            lcout => \U111_CYCLE_SM.N_142_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__6337\,
            in1 => \N__6429\,
            in2 => \N__6023\,
            in3 => \N__6357\,
            lcout => \U111_CYCLE_SM.un7_CYCLE_STATE_0\,
            ltout => \U111_CYCLE_SM.un7_CYCLE_STATE_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__6276\,
            in1 => \N__7439\,
            in2 => \N__6452\,
            in3 => \N__6647\,
            lcout => \U111_CYCLE_SM.N_149\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.BURST_COUNT_RNO_0_1_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__6314\,
            in1 => \N__6442\,
            in2 => \_gnd_net_\,
            in3 => \N__6394\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.N_132_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.BURST_COUNT_1_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000010100000"
        )
    port map (
            in0 => \N__6338\,
            in1 => \N__6358\,
            in2 => \N__6341\,
            in3 => \N__6315\,
            lcout => \U111_CYCLE_SM.BURST_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10576\,
            ce => 'H',
            sr => \N__10291\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7392\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10572\,
            ce => \N__7903\,
            sr => \N__7861\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6285\,
            in1 => \N__6201\,
            in2 => \_gnd_net_\,
            in3 => \N__6635\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_RNIGD6KZ0Z_2\,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_RNIGD6KZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3B1_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6734\,
            in2 => \N__6326\,
            in3 => \N__7234\,
            lcout => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1\,
            ltout => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNI9Q9V1_2_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6323\,
            in3 => \N__6313\,
            lcout => \U111_CYCLE_SM.N_159_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100111111"
        )
    port map (
            in0 => \N__7447\,
            in1 => \N__6286\,
            in2 => \N__6206\,
            in3 => \N__6128\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_srsts_i_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_2_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010001000"
        )
    port map (
            in0 => \N__6733\,
            in1 => \N__7484\,
            in2 => \N__6650\,
            in3 => \N__6636\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_7_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6995\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10567\,
            ce => \N__7904\,
            sr => \N__7872\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7141\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10567\,
            ce => \N__7904\,
            sr => \N__7872\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_0_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7066\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10567\,
            ce => \N__7904\,
            sr => \N__7872\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6613\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10567\,
            ce => \N__7904\,
            sr => \N__7872\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_2_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6918\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10567\,
            ce => \N__7904\,
            sr => \N__7872\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7200\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10567\,
            ce => \N__7904\,
            sr => \N__7872\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6600\,
            in1 => \N__6575\,
            in2 => \_gnd_net_\,
            in3 => \N__8408\,
            lcout => \un1_D_UM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6548\,
            lcout => \GB_BUFFER_CLK80_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8487\,
            in1 => \N__6491\,
            in2 => \_gnd_net_\,
            in3 => \N__8975\,
            lcout => \un2_D_LM_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7223\,
            in1 => \N__7210\,
            in2 => \_gnd_net_\,
            in3 => \N__8442\,
            lcout => \un1_D_UM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7140\,
            in1 => \N__7106\,
            in2 => \_gnd_net_\,
            in3 => \N__8443\,
            lcout => \un1_D_UM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNISP6Q_0_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7065\,
            in1 => \N__7031\,
            in2 => \_gnd_net_\,
            in3 => \N__8446\,
            lcout => \un1_D_UU_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNIA87Q_7_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7007\,
            in1 => \N__6994\,
            in2 => \_gnd_net_\,
            in3 => \N__8445\,
            lcout => \un1_D_UU_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNI0U6Q_2_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8444\,
            in1 => \N__6935\,
            in2 => \_gnd_net_\,
            in3 => \N__6925\,
            lcout => \un1_D_UU_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011101110"
        )
    port map (
            in0 => \N__8763\,
            in1 => \N__6851\,
            in2 => \N__6866\,
            in3 => \N__7473\,
            lcout => \U111_CYCLE_SM.FLIP_WORDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10597\,
            ce => 'H',
            sr => \N__10296\
        );

    \U111_CYCLE_SM.A2_EN_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__6802\,
            in1 => \N__6849\,
            in2 => \_gnd_net_\,
            in3 => \N__6818\,
            lcout => \U111_CYCLE_SM.A2_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10592\,
            ce => 'H',
            sr => \N__10292\
        );

    \U111_CYCLE_SM.LATCH_EN_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__7238\,
            in1 => \N__6790\,
            in2 => \N__8384\,
            in3 => \N__6778\,
            lcout => \U111_CYCLE_SM.LATCH_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10592\,
            ce => 'H',
            sr => \N__10292\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7247\,
            in1 => \N__7282\,
            in2 => \_gnd_net_\,
            in3 => \N__8368\,
            lcout => \un1_D_UM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.PORT_MISMATCH_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__7443\,
            in1 => \N__7537\,
            in2 => \N__7520\,
            in3 => \N__7480\,
            lcout => \U111_CYCLE_SM.PORT_MISMATCHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10583\,
            ce => 'H',
            sr => \N__10293\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8385\,
            in1 => \N__7295\,
            in2 => \_gnd_net_\,
            in3 => \N__7324\,
            lcout => \un1_D_UM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7393\,
            in1 => \N__7358\,
            in2 => \_gnd_net_\,
            in3 => \N__8386\,
            lcout => \un1_D_UM_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7323\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10577\,
            ce => \N__7906\,
            sr => \N__7877\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7281\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10577\,
            ce => \N__7906\,
            sr => \N__7877\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__10823\,
            in1 => \N__12088\,
            in2 => \N__11553\,
            in3 => \N__12527\,
            lcout => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10574\,
            ce => \N__10429\,
            sr => \N__10299\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_6_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8492\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10571\,
            ce => \N__7907\,
            sr => \N__7876\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7637\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10571\,
            ce => \N__7907\,
            sr => \N__7876\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_4_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8544\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10571\,
            ce => \N__7907\,
            sr => \N__7876\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7703\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10571\,
            ce => \N__7907\,
            sr => \N__7876\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_3_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7784\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10571\,
            ce => \N__7907\,
            sr => \N__7876\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_5_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8618\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10571\,
            ce => \N__7907\,
            sr => \N__7876\
        );

    \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11554\,
            in2 => \_gnd_net_\,
            in3 => \N__7829\,
            lcout => \TAn_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNI207Q_3_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8407\,
            in1 => \N__7793\,
            in2 => \_gnd_net_\,
            in3 => \N__7773\,
            lcout => \un1_D_UU_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8437\,
            in1 => \N__7712\,
            in2 => \_gnd_net_\,
            in3 => \N__7698\,
            lcout => \un1_D_UM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7632\,
            in1 => \N__7592\,
            in2 => \_gnd_net_\,
            in3 => \N__8438\,
            lcout => \un1_D_UM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNI647Q_5_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8439\,
            in1 => \N__8630\,
            in2 => \_gnd_net_\,
            in3 => \N__8614\,
            lcout => \un1_D_UU_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNI427Q_4_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8440\,
            in1 => \N__8561\,
            in2 => \_gnd_net_\,
            in3 => \N__8551\,
            lcout => \un1_D_UU_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_esr_RNI867Q_6_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8491\,
            in1 => \N__8441\,
            in2 => \_gnd_net_\,
            in3 => \N__8342\,
            lcout => \un1_D_UU_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8308\,
            in1 => \N__8279\,
            in2 => \_gnd_net_\,
            in3 => \N__8997\,
            lcout => \un1_D_UU_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8240\,
            in1 => \N__8215\,
            in2 => \_gnd_net_\,
            in3 => \N__9008\,
            lcout => \un1_D_UM_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9006\,
            in1 => \N__8156\,
            in2 => \_gnd_net_\,
            in3 => \N__8111\,
            lcout => \un1_D_UM_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8075\,
            in1 => \N__8047\,
            in2 => \_gnd_net_\,
            in3 => \N__8998\,
            lcout => \un1_D_UM_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8974\,
            in1 => \N__7981\,
            in2 => \_gnd_net_\,
            in3 => \N__7946\,
            lcout => \un1_D_UM_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9512\,
            in1 => \N__9476\,
            in2 => \_gnd_net_\,
            in3 => \N__9000\,
            lcout => \un1_D_UU_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__9434\,
            in1 => \N__9412\,
            in2 => \_gnd_net_\,
            in3 => \N__8999\,
            lcout => \un1_D_UU_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9337\,
            in1 => \N__9302\,
            in2 => \_gnd_net_\,
            in3 => \N__9001\,
            lcout => \un1_D_UU_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9002\,
            in1 => \N__9260\,
            in2 => \_gnd_net_\,
            in3 => \N__9235\,
            lcout => \un1_D_UU_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__9185\,
            in1 => \N__9163\,
            in2 => \_gnd_net_\,
            in3 => \N__8984\,
            lcout => \un1_D_UM_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__9110\,
            in1 => \N__9091\,
            in2 => \_gnd_net_\,
            in3 => \N__9018\,
            lcout => \un1_D_UM_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9019\,
            in1 => \N__8716\,
            in2 => \_gnd_net_\,
            in3 => \N__8675\,
            lcout => \un1_D_UM_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep4_i_ess_LC_19_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__12526\,
            in1 => \N__11013\,
            in2 => \N__11932\,
            in3 => \N__11475\,
            lcout => \READ_CYCLE_ACTIVE_rep4_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10578\,
            ce => \N__10432\,
            sr => \N__10304\
        );

    \D_UU_040_iobuf_RNO_4_LC_19_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9620\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_184_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep2_i_ess_LC_20_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__12505\,
            in1 => \N__10930\,
            in2 => \N__11942\,
            in3 => \N__11476\,
            lcout => \READ_CYCLE_ACTIVE_rep2_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10581\,
            ce => \N__10434\,
            sr => \N__10305\
        );

    \D_UU_040_iobuf_RNO_2_LC_20_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9599\,
            lcout => \N_182_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep7_i_ess_LC_22_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__10867\,
            in1 => \N__12443\,
            in2 => \N__12094\,
            in3 => \N__11503\,
            lcout => \READ_CYCLE_ACTIVE_rep7_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10593\,
            ce => \N__10436\,
            sr => \N__10308\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep0_i_ess_LC_22_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__10821\,
            in1 => \N__12444\,
            in2 => \N__11943\,
            in3 => \N__11477\,
            lcout => \READ_CYCLE_ACTIVE_rep0_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10587\,
            ce => \N__10437\,
            sr => \N__10310\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep6_i_ess_LC_22_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__10822\,
            in1 => \N__12445\,
            in2 => \N__11944\,
            in3 => \N__11478\,
            lcout => \READ_CYCLE_ACTIVE_rep6_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10587\,
            ce => \N__10437\,
            sr => \N__10310\
        );

    \D_UU_040_iobuf_RNO_0_LC_22_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9578\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_180_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_040_iobuf_RNO_7_LC_22_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9554\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_187_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_040_iobuf_RNO_6_LC_22_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9533\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_186_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_040_iobuf_RNO_3_LC_23_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9713\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_207_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_040_iobuf_RNO_1_LC_23_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9707\,
            lcout => \N_205_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep27_i_ess_LC_23_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__11014\,
            in1 => \N__12132\,
            in2 => \N__11349\,
            in3 => \N__12705\,
            lcout => \READ_CYCLE_ACTIVE_rep27_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10626\,
            ce => \N__10443\,
            sr => \N__10309\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep25_i_ess_LC_23_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__12595\,
            in1 => \N__11001\,
            in2 => \N__12162\,
            in3 => \N__11465\,
            lcout => \READ_CYCLE_ACTIVE_rep25_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10623\,
            ce => \N__10438\,
            sr => \N__10306\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep30_i_ess_LC_23_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__11002\,
            in1 => \N__12131\,
            in2 => \N__11548\,
            in3 => \N__12596\,
            lcout => \READ_CYCLE_ACTIVE_rep30_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10623\,
            ce => \N__10438\,
            sr => \N__10306\
        );

    \D_LM_040_iobuf_RNO_0_LC_23_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9680\,
            lcout => \N_196_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep16_i_ess_LC_23_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__10925\,
            in1 => \N__12076\,
            in2 => \N__11549\,
            in3 => \N__12591\,
            lcout => \READ_CYCLE_ACTIVE_rep16_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10620\,
            ce => \N__10435\,
            sr => \N__10302\
        );

    \GB_BUFFER_CLK40_THRU_LUT4_0_LC_23_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10631\,
            lcout => \GB_BUFFER_CLK40_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep5_i_ess_LC_23_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__10866\,
            in1 => \N__11953\,
            in2 => \N__12504\,
            in3 => \N__11504\,
            lcout => \READ_CYCLE_ACTIVE_rep5_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10598\,
            ce => \N__10439\,
            sr => \N__10311\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep13_i_ess_LC_23_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__10931\,
            in1 => \N__11945\,
            in2 => \N__11550\,
            in3 => \N__12430\,
            lcout => \READ_CYCLE_ACTIVE_rep13_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10594\,
            ce => \N__10442\,
            sr => \N__10314\
        );

    \D_UU_040_iobuf_RNO_5_LC_23_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9887\,
            lcout => \N_185_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_040_iobuf_RNO_5_LC_23_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9863\,
            lcout => \N_193_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_040_iobuf_RNO_4_LC_24_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9827\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_208_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep28_i_ess_LC_24_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__10929\,
            in1 => \N__12133\,
            in2 => \N__12704\,
            in3 => \N__11358\,
            lcout => \READ_CYCLE_ACTIVE_rep28_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10627\,
            ce => \N__10445\,
            sr => \N__10313\
        );

    \D_LL_040_iobuf_RNO_0_LC_24_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9974\,
            lcout => \N_204_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_040_iobuf_RNO_6_LC_24_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9803\,
            lcout => \N_210_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_040_iobuf_RNO_2_LC_24_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9968\,
            lcout => \N_206_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_040_iobuf_RNO_5_LC_24_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9980\,
            lcout => \N_209_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep29_i_ess_LC_24_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__12594\,
            in1 => \N__10928\,
            in2 => \N__11913\,
            in3 => \N__11363\,
            lcout => \READ_CYCLE_ACTIVE_rep29_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10624\,
            ce => \N__10440\,
            sr => \N__10307\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep24_i_ess_LC_24_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__10926\,
            in1 => \N__11817\,
            in2 => \N__11472\,
            in3 => \N__12592\,
            lcout => \READ_CYCLE_ACTIVE_rep24_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10624\,
            ce => \N__10440\,
            sr => \N__10307\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep26_i_ess_LC_24_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__12593\,
            in1 => \N__10927\,
            in2 => \N__11912\,
            in3 => \N__11362\,
            lcout => \READ_CYCLE_ACTIVE_rep26_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10624\,
            ce => \N__10440\,
            sr => \N__10307\
        );

    \D_LM_040_iobuf_RNO_1_LC_24_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10064\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_197_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LL_040_iobuf_RNO_7_LC_24_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9902\,
            lcout => \N_211_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_040_iobuf_RNO_2_LC_24_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10070\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_198_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_040_iobuf_RNO_3_LC_24_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9893\,
            lcout => \N_199_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep21_i_ess_LC_24_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__12074\,
            in1 => \N__10848\,
            in2 => \N__12503\,
            in3 => \N__11369\,
            lcout => \READ_CYCLE_ACTIVE_rep21_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10618\,
            ce => \N__10433\,
            sr => \N__10301\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep31_i_ess_LC_24_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__10849\,
            in1 => \N__12426\,
            in2 => \N__11474\,
            in3 => \N__12075\,
            lcout => \READ_CYCLE_ACTIVE_rep31_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10618\,
            ce => \N__10433\,
            sr => \N__10301\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep19_i_ess_LC_24_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__12073\,
            in1 => \N__10847\,
            in2 => \N__12502\,
            in3 => \N__11368\,
            lcout => \READ_CYCLE_ACTIVE_rep19_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10618\,
            ce => \N__10433\,
            sr => \N__10301\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep18_i_ess_LC_24_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__10846\,
            in1 => \N__12419\,
            in2 => \N__11473\,
            in3 => \N__12072\,
            lcout => \READ_CYCLE_ACTIVE_rep18_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10618\,
            ce => \N__10433\,
            sr => \N__10301\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep17_i_ess_LC_24_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__12071\,
            in1 => \N__10845\,
            in2 => \N__12501\,
            in3 => \N__11364\,
            lcout => \READ_CYCLE_ACTIVE_rep17_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10618\,
            ce => \N__10433\,
            sr => \N__10301\
        );

    \D_LM_040_iobuf_RNO_4_LC_24_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10016\,
            lcout => \N_200_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_040_iobuf_RNO_0_LC_24_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10010\,
            lcout => \N_188_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_040_iobuf_RNO_5_LC_24_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10031\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_201_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep20_i_ess_LC_24_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__11373\,
            in1 => \N__10840\,
            in2 => \N__12069\,
            in3 => \N__12414\,
            lcout => \READ_CYCLE_ACTIVE_rep20_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10615\,
            ce => \N__10430\,
            sr => \N__10300\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep8_i_ess_LC_24_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__10841\,
            in1 => \N__12415\,
            in2 => \N__12070\,
            in3 => \N__11374\,
            lcout => \READ_CYCLE_ACTIVE_rep8_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10615\,
            ce => \N__10430\,
            sr => \N__10300\
        );

    \D_UM_040_iobuf_RNO_2_LC_24_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10115\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_190_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_040_iobuf_RNO_6_LC_24_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10121\,
            lcout => \N_194_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep22_i_ess_LC_24_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__10764\,
            in1 => \N__12327\,
            in2 => \N__11914\,
            in3 => \N__11377\,
            lcout => \READ_CYCLE_ACTIVE_rep22_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10608\,
            ce => \N__10431\,
            sr => \N__10303\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep23_i_ess_LC_24_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__11378\,
            in1 => \N__10765\,
            in2 => \N__12412\,
            in3 => \N__11829\,
            lcout => \READ_CYCLE_ACTIVE_rep23_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10608\,
            ce => \N__10431\,
            sr => \N__10303\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep14_i_ess_LC_24_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__11376\,
            in1 => \N__10763\,
            in2 => \N__12411\,
            in3 => \N__11825\,
            lcout => \READ_CYCLE_ACTIVE_rep14_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10608\,
            ce => \N__10431\,
            sr => \N__10303\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep10_i_ess_LC_24_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__11375\,
            in1 => \N__10762\,
            in2 => \N__12410\,
            in3 => \N__11824\,
            lcout => \READ_CYCLE_ACTIVE_rep10_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10608\,
            ce => \N__10431\,
            sr => \N__10303\
        );

    \D_LM_040_iobuf_RNO_6_LC_24_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10109\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_202_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_LM_040_iobuf_RNO_7_LC_24_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10091\,
            lcout => \N_203_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep15_i_ess_LC_24_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__10794\,
            in1 => \N__12334\,
            in2 => \N__11816\,
            in3 => \N__11483\,
            lcout => \READ_CYCLE_ACTIVE_rep15_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10602\,
            ce => \N__10441\,
            sr => \N__10312\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep9_i_ess_LC_24_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__10795\,
            in1 => \N__11746\,
            in2 => \N__11551\,
            in3 => \N__12335\,
            lcout => \READ_CYCLE_ACTIVE_rep9_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10602\,
            ce => \N__10441\,
            sr => \N__10312\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep11_i_ess_LC_24_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__11482\,
            in1 => \N__10793\,
            in2 => \N__12413\,
            in3 => \N__11742\,
            lcout => \READ_CYCLE_ACTIVE_rep11_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10602\,
            ce => \N__10441\,
            sr => \N__10312\
        );

    \D_UM_040_iobuf_RNO_1_LC_24_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12782\,
            lcout => \N_189_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_040_iobuf_RNO_3_LC_24_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12761\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_191_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_040_iobuf_RNO_7_LC_24_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12740\,
            lcout => \N_195_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep1_i_ess_LC_24_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__10864\,
            in1 => \N__12337\,
            in2 => \N__12030\,
            in3 => \N__11488\,
            lcout => \READ_CYCLE_ACTIVE_rep1_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10599\,
            ce => \N__10444\,
            sr => \N__10315\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep12_i_ess_LC_24_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__10863\,
            in1 => \N__12336\,
            in2 => \N__12029\,
            in3 => \N__11487\,
            lcout => \READ_CYCLE_ACTIVE_rep12_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10599\,
            ce => \N__10444\,
            sr => \N__10315\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep3_i_ess_LC_24_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__12338\,
            in1 => \N__11952\,
            in2 => \N__11552\,
            in3 => \N__10865\,
            lcout => \READ_CYCLE_ACTIVE_rep3_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10599\,
            ce => \N__10444\,
            sr => \N__10315\
        );

    \D_UU_040_iobuf_RNO_1_LC_24_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10163\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_181_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UM_040_iobuf_RNO_4_LC_24_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10142\,
            lcout => \N_192_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \D_UU_040_iobuf_RNO_3_LC_24_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12800\,
            lcout => \N_183_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 29 2025 20:48:25

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    CMA,
    SIZ,
    DRA,
    A,
    RAMENn,
    TSn,
    LMBEn,
    DMA_LATCH_EN,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    UUBEn,
    LDSn,
    LATCH_CLK,
    CASUn,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    UMBEn,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    RAMSPACEn,
    WEn,
    REGENn,
    LLBEn,
    DBRn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    output [10:0] CMA;
    input [1:0] SIZ;
    input [9:0] DRA;
    input [20:0] A;
    output RAMENn;
    input TSn;
    output LMBEn;
    output DMA_LATCH_EN;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output UUBEn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    output UMBEn;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    output LLBEn;
    input DBRn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__11587;
    wire N__11586;
    wire N__11585;
    wire N__11578;
    wire N__11577;
    wire N__11576;
    wire N__11569;
    wire N__11568;
    wire N__11567;
    wire N__11560;
    wire N__11559;
    wire N__11558;
    wire N__11551;
    wire N__11550;
    wire N__11549;
    wire N__11542;
    wire N__11541;
    wire N__11540;
    wire N__11533;
    wire N__11532;
    wire N__11531;
    wire N__11524;
    wire N__11523;
    wire N__11522;
    wire N__11515;
    wire N__11514;
    wire N__11513;
    wire N__11506;
    wire N__11505;
    wire N__11504;
    wire N__11497;
    wire N__11496;
    wire N__11495;
    wire N__11488;
    wire N__11487;
    wire N__11486;
    wire N__11479;
    wire N__11478;
    wire N__11477;
    wire N__11470;
    wire N__11469;
    wire N__11468;
    wire N__11461;
    wire N__11460;
    wire N__11459;
    wire N__11452;
    wire N__11451;
    wire N__11450;
    wire N__11443;
    wire N__11442;
    wire N__11441;
    wire N__11434;
    wire N__11433;
    wire N__11432;
    wire N__11425;
    wire N__11424;
    wire N__11423;
    wire N__11416;
    wire N__11415;
    wire N__11414;
    wire N__11407;
    wire N__11406;
    wire N__11405;
    wire N__11398;
    wire N__11397;
    wire N__11396;
    wire N__11389;
    wire N__11388;
    wire N__11387;
    wire N__11380;
    wire N__11379;
    wire N__11378;
    wire N__11371;
    wire N__11370;
    wire N__11369;
    wire N__11362;
    wire N__11361;
    wire N__11360;
    wire N__11353;
    wire N__11352;
    wire N__11351;
    wire N__11344;
    wire N__11343;
    wire N__11342;
    wire N__11335;
    wire N__11334;
    wire N__11333;
    wire N__11326;
    wire N__11325;
    wire N__11324;
    wire N__11317;
    wire N__11316;
    wire N__11315;
    wire N__11308;
    wire N__11307;
    wire N__11306;
    wire N__11299;
    wire N__11298;
    wire N__11297;
    wire N__11290;
    wire N__11289;
    wire N__11288;
    wire N__11281;
    wire N__11280;
    wire N__11279;
    wire N__11272;
    wire N__11271;
    wire N__11270;
    wire N__11263;
    wire N__11262;
    wire N__11261;
    wire N__11254;
    wire N__11253;
    wire N__11252;
    wire N__11245;
    wire N__11244;
    wire N__11243;
    wire N__11236;
    wire N__11235;
    wire N__11234;
    wire N__11227;
    wire N__11226;
    wire N__11225;
    wire N__11218;
    wire N__11217;
    wire N__11216;
    wire N__11209;
    wire N__11208;
    wire N__11207;
    wire N__11200;
    wire N__11199;
    wire N__11198;
    wire N__11191;
    wire N__11190;
    wire N__11189;
    wire N__11182;
    wire N__11181;
    wire N__11180;
    wire N__11173;
    wire N__11172;
    wire N__11171;
    wire N__11164;
    wire N__11163;
    wire N__11162;
    wire N__11155;
    wire N__11154;
    wire N__11153;
    wire N__11146;
    wire N__11145;
    wire N__11144;
    wire N__11137;
    wire N__11136;
    wire N__11135;
    wire N__11128;
    wire N__11127;
    wire N__11126;
    wire N__11119;
    wire N__11118;
    wire N__11117;
    wire N__11110;
    wire N__11109;
    wire N__11108;
    wire N__11101;
    wire N__11100;
    wire N__11099;
    wire N__11092;
    wire N__11091;
    wire N__11090;
    wire N__11083;
    wire N__11082;
    wire N__11081;
    wire N__11074;
    wire N__11073;
    wire N__11072;
    wire N__11065;
    wire N__11064;
    wire N__11063;
    wire N__11056;
    wire N__11055;
    wire N__11054;
    wire N__11047;
    wire N__11046;
    wire N__11045;
    wire N__11038;
    wire N__11037;
    wire N__11036;
    wire N__11029;
    wire N__11028;
    wire N__11027;
    wire N__11020;
    wire N__11019;
    wire N__11018;
    wire N__11011;
    wire N__11010;
    wire N__11009;
    wire N__11002;
    wire N__11001;
    wire N__11000;
    wire N__10993;
    wire N__10992;
    wire N__10991;
    wire N__10984;
    wire N__10983;
    wire N__10982;
    wire N__10975;
    wire N__10974;
    wire N__10973;
    wire N__10966;
    wire N__10965;
    wire N__10964;
    wire N__10957;
    wire N__10956;
    wire N__10955;
    wire N__10948;
    wire N__10947;
    wire N__10946;
    wire N__10939;
    wire N__10938;
    wire N__10937;
    wire N__10930;
    wire N__10929;
    wire N__10928;
    wire N__10921;
    wire N__10920;
    wire N__10919;
    wire N__10912;
    wire N__10911;
    wire N__10910;
    wire N__10903;
    wire N__10902;
    wire N__10901;
    wire N__10894;
    wire N__10893;
    wire N__10892;
    wire N__10885;
    wire N__10884;
    wire N__10883;
    wire N__10876;
    wire N__10875;
    wire N__10874;
    wire N__10867;
    wire N__10866;
    wire N__10865;
    wire N__10858;
    wire N__10857;
    wire N__10856;
    wire N__10849;
    wire N__10848;
    wire N__10847;
    wire N__10840;
    wire N__10839;
    wire N__10838;
    wire N__10831;
    wire N__10830;
    wire N__10829;
    wire N__10822;
    wire N__10821;
    wire N__10820;
    wire N__10813;
    wire N__10812;
    wire N__10811;
    wire N__10804;
    wire N__10803;
    wire N__10802;
    wire N__10795;
    wire N__10794;
    wire N__10793;
    wire N__10786;
    wire N__10785;
    wire N__10784;
    wire N__10767;
    wire N__10766;
    wire N__10763;
    wire N__10760;
    wire N__10757;
    wire N__10754;
    wire N__10753;
    wire N__10748;
    wire N__10745;
    wire N__10744;
    wire N__10741;
    wire N__10738;
    wire N__10735;
    wire N__10732;
    wire N__10727;
    wire N__10724;
    wire N__10721;
    wire N__10718;
    wire N__10715;
    wire N__10710;
    wire N__10709;
    wire N__10708;
    wire N__10707;
    wire N__10704;
    wire N__10703;
    wire N__10702;
    wire N__10699;
    wire N__10698;
    wire N__10697;
    wire N__10696;
    wire N__10695;
    wire N__10694;
    wire N__10693;
    wire N__10692;
    wire N__10689;
    wire N__10688;
    wire N__10685;
    wire N__10684;
    wire N__10681;
    wire N__10680;
    wire N__10679;
    wire N__10676;
    wire N__10665;
    wire N__10662;
    wire N__10661;
    wire N__10660;
    wire N__10657;
    wire N__10654;
    wire N__10653;
    wire N__10646;
    wire N__10641;
    wire N__10638;
    wire N__10635;
    wire N__10632;
    wire N__10627;
    wire N__10622;
    wire N__10621;
    wire N__10612;
    wire N__10607;
    wire N__10596;
    wire N__10593;
    wire N__10590;
    wire N__10583;
    wire N__10580;
    wire N__10577;
    wire N__10574;
    wire N__10571;
    wire N__10568;
    wire N__10565;
    wire N__10562;
    wire N__10559;
    wire N__10554;
    wire N__10553;
    wire N__10550;
    wire N__10547;
    wire N__10546;
    wire N__10541;
    wire N__10538;
    wire N__10537;
    wire N__10532;
    wire N__10529;
    wire N__10524;
    wire N__10521;
    wire N__10518;
    wire N__10515;
    wire N__10512;
    wire N__10509;
    wire N__10508;
    wire N__10507;
    wire N__10506;
    wire N__10505;
    wire N__10504;
    wire N__10503;
    wire N__10502;
    wire N__10485;
    wire N__10482;
    wire N__10479;
    wire N__10478;
    wire N__10477;
    wire N__10476;
    wire N__10475;
    wire N__10474;
    wire N__10473;
    wire N__10470;
    wire N__10465;
    wire N__10462;
    wire N__10459;
    wire N__10456;
    wire N__10453;
    wire N__10452;
    wire N__10451;
    wire N__10448;
    wire N__10447;
    wire N__10446;
    wire N__10445;
    wire N__10444;
    wire N__10443;
    wire N__10442;
    wire N__10439;
    wire N__10438;
    wire N__10437;
    wire N__10436;
    wire N__10435;
    wire N__10434;
    wire N__10431;
    wire N__10430;
    wire N__10429;
    wire N__10428;
    wire N__10427;
    wire N__10426;
    wire N__10425;
    wire N__10424;
    wire N__10423;
    wire N__10422;
    wire N__10421;
    wire N__10420;
    wire N__10417;
    wire N__10416;
    wire N__10415;
    wire N__10414;
    wire N__10413;
    wire N__10412;
    wire N__10411;
    wire N__10410;
    wire N__10409;
    wire N__10406;
    wire N__10405;
    wire N__10404;
    wire N__10403;
    wire N__10402;
    wire N__10401;
    wire N__10400;
    wire N__10399;
    wire N__10398;
    wire N__10395;
    wire N__10394;
    wire N__10299;
    wire N__10296;
    wire N__10293;
    wire N__10290;
    wire N__10287;
    wire N__10284;
    wire N__10283;
    wire N__10278;
    wire N__10277;
    wire N__10276;
    wire N__10273;
    wire N__10268;
    wire N__10263;
    wire N__10260;
    wire N__10257;
    wire N__10254;
    wire N__10251;
    wire N__10248;
    wire N__10245;
    wire N__10244;
    wire N__10239;
    wire N__10236;
    wire N__10235;
    wire N__10234;
    wire N__10231;
    wire N__10228;
    wire N__10225;
    wire N__10220;
    wire N__10217;
    wire N__10214;
    wire N__10211;
    wire N__10208;
    wire N__10205;
    wire N__10200;
    wire N__10199;
    wire N__10196;
    wire N__10193;
    wire N__10188;
    wire N__10185;
    wire N__10182;
    wire N__10179;
    wire N__10176;
    wire N__10173;
    wire N__10170;
    wire N__10167;
    wire N__10164;
    wire N__10161;
    wire N__10158;
    wire N__10155;
    wire N__10152;
    wire N__10149;
    wire N__10146;
    wire N__10143;
    wire N__10140;
    wire N__10137;
    wire N__10134;
    wire N__10133;
    wire N__10132;
    wire N__10131;
    wire N__10128;
    wire N__10125;
    wire N__10122;
    wire N__10119;
    wire N__10110;
    wire N__10107;
    wire N__10104;
    wire N__10101;
    wire N__10098;
    wire N__10095;
    wire N__10092;
    wire N__10089;
    wire N__10086;
    wire N__10085;
    wire N__10084;
    wire N__10079;
    wire N__10076;
    wire N__10075;
    wire N__10072;
    wire N__10069;
    wire N__10066;
    wire N__10063;
    wire N__10058;
    wire N__10055;
    wire N__10052;
    wire N__10049;
    wire N__10046;
    wire N__10041;
    wire N__10038;
    wire N__10035;
    wire N__10032;
    wire N__10029;
    wire N__10026;
    wire N__10023;
    wire N__10022;
    wire N__10021;
    wire N__10020;
    wire N__10017;
    wire N__10014;
    wire N__10011;
    wire N__10008;
    wire N__10005;
    wire N__9998;
    wire N__9995;
    wire N__9992;
    wire N__9987;
    wire N__9984;
    wire N__9981;
    wire N__9980;
    wire N__9979;
    wire N__9978;
    wire N__9975;
    wire N__9972;
    wire N__9967;
    wire N__9962;
    wire N__9957;
    wire N__9954;
    wire N__9951;
    wire N__9950;
    wire N__9945;
    wire N__9942;
    wire N__9939;
    wire N__9936;
    wire N__9935;
    wire N__9934;
    wire N__9933;
    wire N__9924;
    wire N__9921;
    wire N__9918;
    wire N__9915;
    wire N__9912;
    wire N__9909;
    wire N__9906;
    wire N__9903;
    wire N__9900;
    wire N__9897;
    wire N__9894;
    wire N__9891;
    wire N__9888;
    wire N__9885;
    wire N__9882;
    wire N__9881;
    wire N__9878;
    wire N__9875;
    wire N__9870;
    wire N__9867;
    wire N__9864;
    wire N__9863;
    wire N__9860;
    wire N__9857;
    wire N__9852;
    wire N__9851;
    wire N__9850;
    wire N__9849;
    wire N__9848;
    wire N__9843;
    wire N__9838;
    wire N__9835;
    wire N__9834;
    wire N__9833;
    wire N__9832;
    wire N__9831;
    wire N__9830;
    wire N__9827;
    wire N__9824;
    wire N__9821;
    wire N__9818;
    wire N__9813;
    wire N__9810;
    wire N__9807;
    wire N__9804;
    wire N__9801;
    wire N__9794;
    wire N__9789;
    wire N__9786;
    wire N__9781;
    wire N__9778;
    wire N__9775;
    wire N__9772;
    wire N__9769;
    wire N__9764;
    wire N__9759;
    wire N__9758;
    wire N__9755;
    wire N__9750;
    wire N__9749;
    wire N__9748;
    wire N__9747;
    wire N__9744;
    wire N__9743;
    wire N__9740;
    wire N__9737;
    wire N__9734;
    wire N__9733;
    wire N__9732;
    wire N__9729;
    wire N__9726;
    wire N__9723;
    wire N__9718;
    wire N__9713;
    wire N__9712;
    wire N__9707;
    wire N__9700;
    wire N__9697;
    wire N__9694;
    wire N__9691;
    wire N__9688;
    wire N__9685;
    wire N__9682;
    wire N__9679;
    wire N__9676;
    wire N__9673;
    wire N__9670;
    wire N__9665;
    wire N__9660;
    wire N__9657;
    wire N__9654;
    wire N__9651;
    wire N__9648;
    wire N__9645;
    wire N__9642;
    wire N__9639;
    wire N__9636;
    wire N__9633;
    wire N__9630;
    wire N__9627;
    wire N__9624;
    wire N__9621;
    wire N__9618;
    wire N__9615;
    wire N__9612;
    wire N__9609;
    wire N__9606;
    wire N__9603;
    wire N__9600;
    wire N__9599;
    wire N__9598;
    wire N__9597;
    wire N__9594;
    wire N__9591;
    wire N__9588;
    wire N__9585;
    wire N__9582;
    wire N__9577;
    wire N__9574;
    wire N__9571;
    wire N__9566;
    wire N__9563;
    wire N__9560;
    wire N__9557;
    wire N__9554;
    wire N__9549;
    wire N__9546;
    wire N__9543;
    wire N__9540;
    wire N__9537;
    wire N__9534;
    wire N__9531;
    wire N__9528;
    wire N__9525;
    wire N__9522;
    wire N__9519;
    wire N__9518;
    wire N__9517;
    wire N__9516;
    wire N__9515;
    wire N__9514;
    wire N__9513;
    wire N__9512;
    wire N__9511;
    wire N__9508;
    wire N__9505;
    wire N__9504;
    wire N__9503;
    wire N__9502;
    wire N__9501;
    wire N__9498;
    wire N__9495;
    wire N__9494;
    wire N__9491;
    wire N__9488;
    wire N__9487;
    wire N__9484;
    wire N__9483;
    wire N__9480;
    wire N__9477;
    wire N__9476;
    wire N__9475;
    wire N__9474;
    wire N__9473;
    wire N__9472;
    wire N__9467;
    wire N__9458;
    wire N__9455;
    wire N__9450;
    wire N__9447;
    wire N__9444;
    wire N__9439;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9424;
    wire N__9423;
    wire N__9422;
    wire N__9417;
    wire N__9414;
    wire N__9405;
    wire N__9400;
    wire N__9397;
    wire N__9396;
    wire N__9393;
    wire N__9388;
    wire N__9385;
    wire N__9382;
    wire N__9379;
    wire N__9378;
    wire N__9375;
    wire N__9372;
    wire N__9369;
    wire N__9366;
    wire N__9361;
    wire N__9358;
    wire N__9351;
    wire N__9348;
    wire N__9345;
    wire N__9342;
    wire N__9329;
    wire N__9326;
    wire N__9323;
    wire N__9312;
    wire N__9309;
    wire N__9306;
    wire N__9303;
    wire N__9300;
    wire N__9299;
    wire N__9296;
    wire N__9295;
    wire N__9294;
    wire N__9291;
    wire N__9288;
    wire N__9285;
    wire N__9284;
    wire N__9283;
    wire N__9282;
    wire N__9281;
    wire N__9280;
    wire N__9279;
    wire N__9278;
    wire N__9275;
    wire N__9274;
    wire N__9273;
    wire N__9272;
    wire N__9267;
    wire N__9264;
    wire N__9259;
    wire N__9252;
    wire N__9251;
    wire N__9250;
    wire N__9245;
    wire N__9244;
    wire N__9241;
    wire N__9236;
    wire N__9235;
    wire N__9232;
    wire N__9223;
    wire N__9218;
    wire N__9215;
    wire N__9214;
    wire N__9213;
    wire N__9210;
    wire N__9209;
    wire N__9206;
    wire N__9203;
    wire N__9200;
    wire N__9199;
    wire N__9198;
    wire N__9197;
    wire N__9194;
    wire N__9187;
    wire N__9180;
    wire N__9177;
    wire N__9170;
    wire N__9167;
    wire N__9162;
    wire N__9155;
    wire N__9150;
    wire N__9141;
    wire N__9138;
    wire N__9135;
    wire N__9132;
    wire N__9129;
    wire N__9126;
    wire N__9123;
    wire N__9120;
    wire N__9117;
    wire N__9114;
    wire N__9111;
    wire N__9108;
    wire N__9105;
    wire N__9102;
    wire N__9099;
    wire N__9096;
    wire N__9095;
    wire N__9094;
    wire N__9091;
    wire N__9086;
    wire N__9085;
    wire N__9084;
    wire N__9079;
    wire N__9076;
    wire N__9075;
    wire N__9074;
    wire N__9073;
    wire N__9070;
    wire N__9065;
    wire N__9062;
    wire N__9059;
    wire N__9056;
    wire N__9045;
    wire N__9044;
    wire N__9043;
    wire N__9042;
    wire N__9041;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9031;
    wire N__9028;
    wire N__9021;
    wire N__9018;
    wire N__9015;
    wire N__9012;
    wire N__9007;
    wire N__9004;
    wire N__8999;
    wire N__8994;
    wire N__8991;
    wire N__8988;
    wire N__8985;
    wire N__8982;
    wire N__8979;
    wire N__8976;
    wire N__8973;
    wire N__8970;
    wire N__8967;
    wire N__8966;
    wire N__8965;
    wire N__8964;
    wire N__8963;
    wire N__8962;
    wire N__8961;
    wire N__8960;
    wire N__8959;
    wire N__8958;
    wire N__8957;
    wire N__8956;
    wire N__8955;
    wire N__8954;
    wire N__8953;
    wire N__8952;
    wire N__8951;
    wire N__8950;
    wire N__8949;
    wire N__8948;
    wire N__8947;
    wire N__8946;
    wire N__8945;
    wire N__8944;
    wire N__8943;
    wire N__8940;
    wire N__8939;
    wire N__8938;
    wire N__8937;
    wire N__8936;
    wire N__8935;
    wire N__8934;
    wire N__8933;
    wire N__8932;
    wire N__8931;
    wire N__8930;
    wire N__8929;
    wire N__8928;
    wire N__8927;
    wire N__8926;
    wire N__8925;
    wire N__8844;
    wire N__8841;
    wire N__8838;
    wire N__8837;
    wire N__8836;
    wire N__8835;
    wire N__8832;
    wire N__8831;
    wire N__8828;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8815;
    wire N__8812;
    wire N__8807;
    wire N__8802;
    wire N__8799;
    wire N__8796;
    wire N__8793;
    wire N__8788;
    wire N__8781;
    wire N__8778;
    wire N__8775;
    wire N__8772;
    wire N__8769;
    wire N__8766;
    wire N__8763;
    wire N__8760;
    wire N__8759;
    wire N__8754;
    wire N__8751;
    wire N__8748;
    wire N__8745;
    wire N__8742;
    wire N__8739;
    wire N__8736;
    wire N__8733;
    wire N__8730;
    wire N__8727;
    wire N__8724;
    wire N__8721;
    wire N__8718;
    wire N__8715;
    wire N__8712;
    wire N__8709;
    wire N__8706;
    wire N__8703;
    wire N__8700;
    wire N__8697;
    wire N__8694;
    wire N__8691;
    wire N__8688;
    wire N__8685;
    wire N__8682;
    wire N__8679;
    wire N__8676;
    wire N__8673;
    wire N__8670;
    wire N__8667;
    wire N__8664;
    wire N__8661;
    wire N__8658;
    wire N__8655;
    wire N__8652;
    wire N__8649;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8631;
    wire N__8628;
    wire N__8625;
    wire N__8624;
    wire N__8621;
    wire N__8618;
    wire N__8615;
    wire N__8610;
    wire N__8607;
    wire N__8604;
    wire N__8601;
    wire N__8598;
    wire N__8595;
    wire N__8594;
    wire N__8593;
    wire N__8592;
    wire N__8587;
    wire N__8582;
    wire N__8581;
    wire N__8578;
    wire N__8575;
    wire N__8574;
    wire N__8571;
    wire N__8570;
    wire N__8567;
    wire N__8564;
    wire N__8561;
    wire N__8556;
    wire N__8553;
    wire N__8550;
    wire N__8545;
    wire N__8544;
    wire N__8541;
    wire N__8536;
    wire N__8533;
    wire N__8526;
    wire N__8523;
    wire N__8520;
    wire N__8517;
    wire N__8516;
    wire N__8515;
    wire N__8512;
    wire N__8509;
    wire N__8506;
    wire N__8505;
    wire N__8502;
    wire N__8499;
    wire N__8496;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8484;
    wire N__8479;
    wire N__8476;
    wire N__8473;
    wire N__8470;
    wire N__8463;
    wire N__8460;
    wire N__8457;
    wire N__8454;
    wire N__8451;
    wire N__8448;
    wire N__8445;
    wire N__8444;
    wire N__8441;
    wire N__8438;
    wire N__8437;
    wire N__8434;
    wire N__8433;
    wire N__8430;
    wire N__8427;
    wire N__8424;
    wire N__8423;
    wire N__8422;
    wire N__8419;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire N__8404;
    wire N__8401;
    wire N__8398;
    wire N__8391;
    wire N__8388;
    wire N__8379;
    wire N__8376;
    wire N__8373;
    wire N__8370;
    wire N__8367;
    wire N__8364;
    wire N__8361;
    wire N__8358;
    wire N__8357;
    wire N__8354;
    wire N__8351;
    wire N__8348;
    wire N__8347;
    wire N__8346;
    wire N__8341;
    wire N__8338;
    wire N__8337;
    wire N__8334;
    wire N__8329;
    wire N__8326;
    wire N__8319;
    wire N__8316;
    wire N__8313;
    wire N__8310;
    wire N__8307;
    wire N__8304;
    wire N__8301;
    wire N__8298;
    wire N__8295;
    wire N__8294;
    wire N__8289;
    wire N__8286;
    wire N__8285;
    wire N__8284;
    wire N__8281;
    wire N__8276;
    wire N__8273;
    wire N__8270;
    wire N__8265;
    wire N__8262;
    wire N__8259;
    wire N__8256;
    wire N__8253;
    wire N__8250;
    wire N__8247;
    wire N__8244;
    wire N__8241;
    wire N__8238;
    wire N__8235;
    wire N__8232;
    wire N__8229;
    wire N__8226;
    wire N__8223;
    wire N__8220;
    wire N__8217;
    wire N__8214;
    wire N__8211;
    wire N__8208;
    wire N__8205;
    wire N__8202;
    wire N__8199;
    wire N__8196;
    wire N__8193;
    wire N__8190;
    wire N__8187;
    wire N__8184;
    wire N__8181;
    wire N__8178;
    wire N__8175;
    wire N__8172;
    wire N__8169;
    wire N__8166;
    wire N__8163;
    wire N__8160;
    wire N__8157;
    wire N__8154;
    wire N__8151;
    wire N__8148;
    wire N__8147;
    wire N__8142;
    wire N__8139;
    wire N__8138;
    wire N__8137;
    wire N__8134;
    wire N__8129;
    wire N__8124;
    wire N__8121;
    wire N__8118;
    wire N__8115;
    wire N__8112;
    wire N__8109;
    wire N__8106;
    wire N__8103;
    wire N__8102;
    wire N__8101;
    wire N__8098;
    wire N__8097;
    wire N__8094;
    wire N__8093;
    wire N__8090;
    wire N__8089;
    wire N__8086;
    wire N__8083;
    wire N__8080;
    wire N__8077;
    wire N__8076;
    wire N__8073;
    wire N__8070;
    wire N__8065;
    wire N__8062;
    wire N__8059;
    wire N__8056;
    wire N__8053;
    wire N__8048;
    wire N__8043;
    wire N__8040;
    wire N__8031;
    wire N__8028;
    wire N__8025;
    wire N__8022;
    wire N__8019;
    wire N__8016;
    wire N__8013;
    wire N__8010;
    wire N__8007;
    wire N__8004;
    wire N__8001;
    wire N__7998;
    wire N__7995;
    wire N__7992;
    wire N__7989;
    wire N__7986;
    wire N__7983;
    wire N__7980;
    wire N__7977;
    wire N__7974;
    wire N__7971;
    wire N__7968;
    wire N__7965;
    wire N__7962;
    wire N__7959;
    wire N__7956;
    wire N__7953;
    wire N__7950;
    wire N__7947;
    wire N__7944;
    wire N__7941;
    wire N__7938;
    wire N__7935;
    wire N__7932;
    wire N__7929;
    wire N__7926;
    wire N__7923;
    wire N__7920;
    wire N__7917;
    wire N__7914;
    wire N__7911;
    wire N__7908;
    wire N__7905;
    wire N__7902;
    wire N__7901;
    wire N__7900;
    wire N__7899;
    wire N__7898;
    wire N__7897;
    wire N__7894;
    wire N__7889;
    wire N__7886;
    wire N__7883;
    wire N__7880;
    wire N__7877;
    wire N__7876;
    wire N__7871;
    wire N__7868;
    wire N__7865;
    wire N__7864;
    wire N__7861;
    wire N__7858;
    wire N__7853;
    wire N__7850;
    wire N__7847;
    wire N__7836;
    wire N__7833;
    wire N__7832;
    wire N__7831;
    wire N__7828;
    wire N__7827;
    wire N__7824;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7814;
    wire N__7811;
    wire N__7808;
    wire N__7805;
    wire N__7800;
    wire N__7797;
    wire N__7794;
    wire N__7793;
    wire N__7790;
    wire N__7787;
    wire N__7782;
    wire N__7779;
    wire N__7776;
    wire N__7773;
    wire N__7770;
    wire N__7767;
    wire N__7764;
    wire N__7761;
    wire N__7758;
    wire N__7755;
    wire N__7752;
    wire N__7749;
    wire N__7744;
    wire N__7737;
    wire N__7734;
    wire N__7733;
    wire N__7730;
    wire N__7727;
    wire N__7726;
    wire N__7725;
    wire N__7724;
    wire N__7721;
    wire N__7718;
    wire N__7713;
    wire N__7710;
    wire N__7707;
    wire N__7700;
    wire N__7697;
    wire N__7694;
    wire N__7693;
    wire N__7688;
    wire N__7685;
    wire N__7680;
    wire N__7677;
    wire N__7674;
    wire N__7671;
    wire N__7668;
    wire N__7665;
    wire N__7662;
    wire N__7659;
    wire N__7656;
    wire N__7653;
    wire N__7650;
    wire N__7647;
    wire N__7644;
    wire N__7641;
    wire N__7638;
    wire N__7635;
    wire N__7632;
    wire N__7629;
    wire N__7626;
    wire N__7623;
    wire N__7620;
    wire N__7617;
    wire N__7614;
    wire N__7611;
    wire N__7608;
    wire N__7605;
    wire N__7602;
    wire N__7599;
    wire N__7596;
    wire N__7593;
    wire N__7590;
    wire N__7587;
    wire N__7584;
    wire N__7581;
    wire N__7578;
    wire N__7575;
    wire N__7572;
    wire N__7569;
    wire N__7566;
    wire N__7563;
    wire N__7560;
    wire N__7557;
    wire N__7554;
    wire N__7553;
    wire N__7552;
    wire N__7551;
    wire N__7550;
    wire N__7547;
    wire N__7544;
    wire N__7541;
    wire N__7536;
    wire N__7531;
    wire N__7528;
    wire N__7527;
    wire N__7524;
    wire N__7521;
    wire N__7518;
    wire N__7515;
    wire N__7512;
    wire N__7507;
    wire N__7504;
    wire N__7501;
    wire N__7498;
    wire N__7495;
    wire N__7492;
    wire N__7489;
    wire N__7486;
    wire N__7481;
    wire N__7476;
    wire N__7473;
    wire N__7470;
    wire N__7467;
    wire N__7464;
    wire N__7461;
    wire N__7458;
    wire N__7455;
    wire N__7452;
    wire N__7449;
    wire N__7446;
    wire N__7443;
    wire N__7440;
    wire N__7437;
    wire N__7434;
    wire N__7431;
    wire N__7428;
    wire N__7425;
    wire N__7422;
    wire N__7419;
    wire N__7416;
    wire N__7413;
    wire N__7410;
    wire N__7407;
    wire N__7404;
    wire N__7401;
    wire N__7398;
    wire N__7395;
    wire N__7392;
    wire N__7389;
    wire N__7386;
    wire N__7383;
    wire N__7380;
    wire N__7377;
    wire N__7376;
    wire N__7375;
    wire N__7374;
    wire N__7373;
    wire N__7372;
    wire N__7367;
    wire N__7362;
    wire N__7357;
    wire N__7356;
    wire N__7355;
    wire N__7354;
    wire N__7353;
    wire N__7346;
    wire N__7343;
    wire N__7342;
    wire N__7339;
    wire N__7336;
    wire N__7333;
    wire N__7332;
    wire N__7331;
    wire N__7330;
    wire N__7329;
    wire N__7324;
    wire N__7321;
    wire N__7318;
    wire N__7315;
    wire N__7312;
    wire N__7307;
    wire N__7304;
    wire N__7301;
    wire N__7296;
    wire N__7293;
    wire N__7282;
    wire N__7281;
    wire N__7278;
    wire N__7273;
    wire N__7270;
    wire N__7263;
    wire N__7260;
    wire N__7257;
    wire N__7254;
    wire N__7251;
    wire N__7248;
    wire N__7245;
    wire N__7242;
    wire N__7239;
    wire N__7236;
    wire N__7233;
    wire N__7230;
    wire N__7227;
    wire N__7224;
    wire N__7221;
    wire N__7218;
    wire N__7215;
    wire N__7212;
    wire N__7209;
    wire N__7206;
    wire N__7203;
    wire N__7200;
    wire N__7197;
    wire N__7194;
    wire N__7191;
    wire N__7188;
    wire N__7187;
    wire N__7184;
    wire N__7181;
    wire N__7176;
    wire N__7175;
    wire N__7172;
    wire N__7169;
    wire N__7164;
    wire N__7163;
    wire N__7160;
    wire N__7157;
    wire N__7152;
    wire N__7149;
    wire N__7146;
    wire N__7143;
    wire N__7140;
    wire N__7137;
    wire N__7136;
    wire N__7133;
    wire N__7130;
    wire N__7127;
    wire N__7124;
    wire N__7121;
    wire N__7118;
    wire N__7113;
    wire N__7110;
    wire N__7107;
    wire N__7104;
    wire N__7101;
    wire N__7098;
    wire N__7095;
    wire N__7092;
    wire N__7091;
    wire N__7086;
    wire N__7083;
    wire N__7080;
    wire N__7077;
    wire N__7074;
    wire N__7071;
    wire N__7068;
    wire N__7067;
    wire N__7064;
    wire N__7063;
    wire N__7062;
    wire N__7059;
    wire N__7056;
    wire N__7051;
    wire N__7044;
    wire N__7041;
    wire N__7038;
    wire N__7035;
    wire N__7032;
    wire N__7029;
    wire N__7026;
    wire N__7025;
    wire N__7022;
    wire N__7019;
    wire N__7018;
    wire N__7013;
    wire N__7010;
    wire N__7007;
    wire N__7004;
    wire N__7001;
    wire N__6998;
    wire N__6995;
    wire N__6992;
    wire N__6989;
    wire N__6986;
    wire N__6983;
    wire N__6980;
    wire N__6975;
    wire N__6974;
    wire N__6973;
    wire N__6968;
    wire N__6965;
    wire N__6960;
    wire N__6959;
    wire N__6956;
    wire N__6953;
    wire N__6950;
    wire N__6945;
    wire N__6942;
    wire N__6939;
    wire N__6936;
    wire N__6933;
    wire N__6930;
    wire N__6927;
    wire N__6924;
    wire N__6921;
    wire N__6918;
    wire N__6915;
    wire N__6912;
    wire N__6911;
    wire N__6908;
    wire N__6905;
    wire N__6900;
    wire N__6897;
    wire N__6896;
    wire N__6893;
    wire N__6890;
    wire N__6885;
    wire N__6882;
    wire N__6879;
    wire N__6876;
    wire N__6875;
    wire N__6872;
    wire N__6869;
    wire N__6864;
    wire N__6863;
    wire N__6862;
    wire N__6861;
    wire N__6860;
    wire N__6859;
    wire N__6846;
    wire N__6843;
    wire N__6840;
    wire N__6839;
    wire N__6836;
    wire N__6833;
    wire N__6830;
    wire N__6827;
    wire N__6822;
    wire N__6819;
    wire N__6816;
    wire N__6813;
    wire N__6812;
    wire N__6809;
    wire N__6806;
    wire N__6803;
    wire N__6798;
    wire N__6797;
    wire N__6794;
    wire N__6793;
    wire N__6792;
    wire N__6791;
    wire N__6790;
    wire N__6787;
    wire N__6786;
    wire N__6785;
    wire N__6784;
    wire N__6781;
    wire N__6778;
    wire N__6775;
    wire N__6770;
    wire N__6769;
    wire N__6768;
    wire N__6765;
    wire N__6762;
    wire N__6759;
    wire N__6756;
    wire N__6755;
    wire N__6754;
    wire N__6747;
    wire N__6746;
    wire N__6743;
    wire N__6742;
    wire N__6741;
    wire N__6740;
    wire N__6737;
    wire N__6734;
    wire N__6729;
    wire N__6724;
    wire N__6721;
    wire N__6718;
    wire N__6715;
    wire N__6712;
    wire N__6709;
    wire N__6702;
    wire N__6681;
    wire N__6680;
    wire N__6675;
    wire N__6672;
    wire N__6669;
    wire N__6666;
    wire N__6665;
    wire N__6664;
    wire N__6661;
    wire N__6658;
    wire N__6655;
    wire N__6648;
    wire N__6647;
    wire N__6644;
    wire N__6643;
    wire N__6640;
    wire N__6637;
    wire N__6636;
    wire N__6633;
    wire N__6630;
    wire N__6627;
    wire N__6624;
    wire N__6615;
    wire N__6614;
    wire N__6611;
    wire N__6610;
    wire N__6607;
    wire N__6604;
    wire N__6601;
    wire N__6596;
    wire N__6593;
    wire N__6590;
    wire N__6585;
    wire N__6584;
    wire N__6583;
    wire N__6582;
    wire N__6579;
    wire N__6572;
    wire N__6567;
    wire N__6564;
    wire N__6561;
    wire N__6558;
    wire N__6557;
    wire N__6554;
    wire N__6551;
    wire N__6546;
    wire N__6543;
    wire N__6542;
    wire N__6539;
    wire N__6536;
    wire N__6531;
    wire N__6530;
    wire N__6527;
    wire N__6524;
    wire N__6519;
    wire N__6516;
    wire N__6515;
    wire N__6512;
    wire N__6509;
    wire N__6506;
    wire N__6501;
    wire N__6500;
    wire N__6499;
    wire N__6498;
    wire N__6497;
    wire N__6496;
    wire N__6493;
    wire N__6490;
    wire N__6487;
    wire N__6484;
    wire N__6479;
    wire N__6468;
    wire N__6467;
    wire N__6464;
    wire N__6461;
    wire N__6456;
    wire N__6455;
    wire N__6454;
    wire N__6453;
    wire N__6452;
    wire N__6451;
    wire N__6448;
    wire N__6445;
    wire N__6442;
    wire N__6435;
    wire N__6426;
    wire N__6425;
    wire N__6422;
    wire N__6419;
    wire N__6414;
    wire N__6411;
    wire N__6410;
    wire N__6409;
    wire N__6406;
    wire N__6405;
    wire N__6400;
    wire N__6399;
    wire N__6398;
    wire N__6397;
    wire N__6394;
    wire N__6393;
    wire N__6392;
    wire N__6391;
    wire N__6390;
    wire N__6387;
    wire N__6384;
    wire N__6381;
    wire N__6376;
    wire N__6373;
    wire N__6368;
    wire N__6363;
    wire N__6358;
    wire N__6355;
    wire N__6342;
    wire N__6339;
    wire N__6338;
    wire N__6335;
    wire N__6332;
    wire N__6329;
    wire N__6326;
    wire N__6323;
    wire N__6320;
    wire N__6317;
    wire N__6314;
    wire N__6309;
    wire N__6306;
    wire N__6303;
    wire N__6300;
    wire N__6299;
    wire N__6298;
    wire N__6295;
    wire N__6292;
    wire N__6289;
    wire N__6284;
    wire N__6283;
    wire N__6280;
    wire N__6277;
    wire N__6274;
    wire N__6271;
    wire N__6266;
    wire N__6263;
    wire N__6260;
    wire N__6257;
    wire N__6254;
    wire N__6249;
    wire N__6246;
    wire N__6243;
    wire N__6242;
    wire N__6239;
    wire N__6238;
    wire N__6237;
    wire N__6236;
    wire N__6235;
    wire N__6232;
    wire N__6229;
    wire N__6226;
    wire N__6223;
    wire N__6218;
    wire N__6217;
    wire N__6214;
    wire N__6209;
    wire N__6206;
    wire N__6203;
    wire N__6200;
    wire N__6197;
    wire N__6188;
    wire N__6183;
    wire N__6180;
    wire N__6177;
    wire N__6174;
    wire N__6171;
    wire N__6168;
    wire N__6165;
    wire N__6162;
    wire N__6159;
    wire N__6158;
    wire N__6157;
    wire N__6156;
    wire N__6155;
    wire N__6154;
    wire N__6151;
    wire N__6148;
    wire N__6147;
    wire N__6144;
    wire N__6141;
    wire N__6136;
    wire N__6131;
    wire N__6128;
    wire N__6123;
    wire N__6114;
    wire N__6111;
    wire N__6108;
    wire N__6105;
    wire N__6102;
    wire N__6099;
    wire N__6096;
    wire N__6093;
    wire N__6090;
    wire N__6087;
    wire N__6084;
    wire N__6081;
    wire N__6078;
    wire N__6077;
    wire N__6074;
    wire N__6071;
    wire N__6066;
    wire N__6065;
    wire N__6062;
    wire N__6059;
    wire N__6054;
    wire N__6053;
    wire N__6048;
    wire N__6045;
    wire N__6042;
    wire N__6041;
    wire N__6040;
    wire N__6037;
    wire N__6036;
    wire N__6035;
    wire N__6034;
    wire N__6033;
    wire N__6032;
    wire N__6031;
    wire N__6026;
    wire N__6023;
    wire N__6022;
    wire N__6021;
    wire N__6018;
    wire N__6015;
    wire N__6014;
    wire N__6013;
    wire N__6012;
    wire N__6011;
    wire N__6008;
    wire N__6007;
    wire N__6006;
    wire N__6005;
    wire N__6002;
    wire N__6001;
    wire N__5996;
    wire N__5995;
    wire N__5992;
    wire N__5989;
    wire N__5986;
    wire N__5983;
    wire N__5978;
    wire N__5975;
    wire N__5968;
    wire N__5961;
    wire N__5954;
    wire N__5951;
    wire N__5948;
    wire N__5925;
    wire N__5924;
    wire N__5923;
    wire N__5922;
    wire N__5921;
    wire N__5918;
    wire N__5911;
    wire N__5910;
    wire N__5909;
    wire N__5908;
    wire N__5907;
    wire N__5904;
    wire N__5899;
    wire N__5896;
    wire N__5891;
    wire N__5888;
    wire N__5877;
    wire N__5876;
    wire N__5875;
    wire N__5874;
    wire N__5873;
    wire N__5872;
    wire N__5867;
    wire N__5864;
    wire N__5863;
    wire N__5862;
    wire N__5861;
    wire N__5860;
    wire N__5857;
    wire N__5856;
    wire N__5851;
    wire N__5848;
    wire N__5845;
    wire N__5840;
    wire N__5835;
    wire N__5834;
    wire N__5831;
    wire N__5828;
    wire N__5819;
    wire N__5816;
    wire N__5813;
    wire N__5810;
    wire N__5799;
    wire N__5798;
    wire N__5797;
    wire N__5794;
    wire N__5793;
    wire N__5790;
    wire N__5789;
    wire N__5786;
    wire N__5785;
    wire N__5784;
    wire N__5783;
    wire N__5782;
    wire N__5779;
    wire N__5776;
    wire N__5775;
    wire N__5772;
    wire N__5769;
    wire N__5766;
    wire N__5763;
    wire N__5762;
    wire N__5761;
    wire N__5760;
    wire N__5757;
    wire N__5752;
    wire N__5751;
    wire N__5750;
    wire N__5747;
    wire N__5744;
    wire N__5741;
    wire N__5734;
    wire N__5729;
    wire N__5722;
    wire N__5719;
    wire N__5714;
    wire N__5697;
    wire N__5696;
    wire N__5693;
    wire N__5692;
    wire N__5691;
    wire N__5688;
    wire N__5685;
    wire N__5684;
    wire N__5683;
    wire N__5680;
    wire N__5677;
    wire N__5672;
    wire N__5671;
    wire N__5670;
    wire N__5667;
    wire N__5666;
    wire N__5665;
    wire N__5664;
    wire N__5663;
    wire N__5660;
    wire N__5657;
    wire N__5652;
    wire N__5643;
    wire N__5638;
    wire N__5635;
    wire N__5622;
    wire N__5619;
    wire N__5618;
    wire N__5615;
    wire N__5612;
    wire N__5607;
    wire N__5604;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5592;
    wire N__5589;
    wire N__5586;
    wire N__5583;
    wire N__5582;
    wire N__5581;
    wire N__5578;
    wire N__5577;
    wire N__5576;
    wire N__5575;
    wire N__5574;
    wire N__5573;
    wire N__5572;
    wire N__5567;
    wire N__5564;
    wire N__5561;
    wire N__5558;
    wire N__5555;
    wire N__5552;
    wire N__5547;
    wire N__5532;
    wire N__5529;
    wire N__5526;
    wire N__5523;
    wire N__5520;
    wire N__5517;
    wire N__5514;
    wire N__5511;
    wire N__5510;
    wire N__5507;
    wire N__5504;
    wire N__5501;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5489;
    wire N__5486;
    wire N__5483;
    wire N__5480;
    wire N__5475;
    wire N__5472;
    wire N__5469;
    wire N__5466;
    wire N__5463;
    wire N__5460;
    wire N__5457;
    wire N__5454;
    wire N__5451;
    wire N__5448;
    wire N__5447;
    wire N__5444;
    wire N__5443;
    wire N__5442;
    wire N__5439;
    wire N__5436;
    wire N__5433;
    wire N__5430;
    wire N__5421;
    wire N__5418;
    wire N__5415;
    wire N__5412;
    wire N__5409;
    wire N__5406;
    wire N__5403;
    wire N__5400;
    wire N__5399;
    wire N__5398;
    wire N__5397;
    wire N__5396;
    wire N__5393;
    wire N__5392;
    wire N__5391;
    wire N__5388;
    wire N__5385;
    wire N__5384;
    wire N__5379;
    wire N__5376;
    wire N__5375;
    wire N__5370;
    wire N__5367;
    wire N__5364;
    wire N__5361;
    wire N__5358;
    wire N__5355;
    wire N__5352;
    wire N__5349;
    wire N__5334;
    wire N__5333;
    wire N__5332;
    wire N__5331;
    wire N__5328;
    wire N__5327;
    wire N__5324;
    wire N__5321;
    wire N__5318;
    wire N__5315;
    wire N__5312;
    wire N__5307;
    wire N__5304;
    wire N__5297;
    wire N__5294;
    wire N__5291;
    wire N__5286;
    wire N__5283;
    wire N__5280;
    wire N__5277;
    wire N__5276;
    wire N__5273;
    wire N__5270;
    wire N__5267;
    wire N__5262;
    wire N__5261;
    wire N__5260;
    wire N__5257;
    wire N__5254;
    wire N__5251;
    wire N__5248;
    wire N__5245;
    wire N__5238;
    wire N__5235;
    wire N__5232;
    wire N__5229;
    wire N__5226;
    wire N__5223;
    wire N__5220;
    wire N__5217;
    wire N__5216;
    wire N__5215;
    wire N__5214;
    wire N__5213;
    wire N__5212;
    wire N__5211;
    wire N__5208;
    wire N__5201;
    wire N__5194;
    wire N__5187;
    wire N__5184;
    wire N__5181;
    wire N__5180;
    wire N__5177;
    wire N__5176;
    wire N__5173;
    wire N__5170;
    wire N__5167;
    wire N__5160;
    wire N__5159;
    wire N__5156;
    wire N__5153;
    wire N__5148;
    wire N__5147;
    wire N__5144;
    wire N__5141;
    wire N__5136;
    wire N__5133;
    wire N__5132;
    wire N__5129;
    wire N__5126;
    wire N__5123;
    wire N__5118;
    wire N__5117;
    wire N__5114;
    wire N__5111;
    wire N__5106;
    wire N__5103;
    wire N__5100;
    wire N__5097;
    wire N__5094;
    wire N__5091;
    wire N__5088;
    wire N__5085;
    wire N__5082;
    wire N__5079;
    wire N__5076;
    wire N__5073;
    wire N__5070;
    wire N__5069;
    wire N__5066;
    wire N__5063;
    wire N__5058;
    wire N__5057;
    wire N__5056;
    wire N__5055;
    wire N__5052;
    wire N__5049;
    wire N__5046;
    wire N__5043;
    wire N__5040;
    wire N__5033;
    wire N__5032;
    wire N__5031;
    wire N__5026;
    wire N__5021;
    wire N__5016;
    wire N__5013;
    wire N__5010;
    wire N__5007;
    wire N__5006;
    wire N__5005;
    wire N__5004;
    wire N__5001;
    wire N__4996;
    wire N__4993;
    wire N__4986;
    wire N__4983;
    wire N__4982;
    wire N__4979;
    wire N__4976;
    wire N__4971;
    wire N__4968;
    wire N__4965;
    wire N__4962;
    wire N__4959;
    wire N__4956;
    wire N__4953;
    wire N__4950;
    wire N__4947;
    wire N__4944;
    wire N__4943;
    wire N__4940;
    wire N__4937;
    wire N__4932;
    wire N__4929;
    wire N__4926;
    wire N__4923;
    wire N__4920;
    wire N__4917;
    wire N__4916;
    wire N__4913;
    wire N__4910;
    wire N__4905;
    wire N__4902;
    wire N__4899;
    wire N__4896;
    wire N__4893;
    wire N__4890;
    wire N__4887;
    wire N__4884;
    wire N__4881;
    wire N__4880;
    wire N__4877;
    wire N__4876;
    wire N__4875;
    wire N__4872;
    wire N__4869;
    wire N__4864;
    wire N__4857;
    wire N__4854;
    wire N__4851;
    wire N__4850;
    wire N__4849;
    wire N__4846;
    wire N__4841;
    wire N__4836;
    wire N__4833;
    wire N__4830;
    wire N__4827;
    wire N__4824;
    wire N__4821;
    wire N__4820;
    wire N__4817;
    wire N__4814;
    wire N__4813;
    wire N__4812;
    wire N__4811;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4799;
    wire N__4796;
    wire N__4785;
    wire N__4782;
    wire N__4779;
    wire N__4776;
    wire N__4773;
    wire N__4770;
    wire N__4767;
    wire N__4764;
    wire N__4763;
    wire N__4762;
    wire N__4759;
    wire N__4756;
    wire N__4753;
    wire N__4746;
    wire N__4745;
    wire N__4740;
    wire N__4737;
    wire N__4734;
    wire N__4731;
    wire N__4728;
    wire N__4725;
    wire N__4722;
    wire N__4719;
    wire N__4718;
    wire N__4717;
    wire N__4714;
    wire N__4711;
    wire N__4708;
    wire N__4705;
    wire N__4702;
    wire N__4699;
    wire N__4698;
    wire N__4697;
    wire N__4694;
    wire N__4689;
    wire N__4684;
    wire N__4677;
    wire N__4674;
    wire N__4671;
    wire N__4668;
    wire N__4665;
    wire N__4662;
    wire N__4659;
    wire N__4656;
    wire N__4653;
    wire N__4650;
    wire N__4647;
    wire N__4644;
    wire N__4641;
    wire N__4638;
    wire N__4635;
    wire N__4632;
    wire N__4629;
    wire N__4626;
    wire N__4623;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4613;
    wire N__4608;
    wire N__4607;
    wire N__4606;
    wire N__4605;
    wire N__4602;
    wire N__4599;
    wire N__4592;
    wire N__4587;
    wire N__4584;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4573;
    wire N__4572;
    wire N__4569;
    wire N__4566;
    wire N__4561;
    wire N__4554;
    wire N__4551;
    wire N__4548;
    wire N__4545;
    wire N__4542;
    wire N__4539;
    wire N__4536;
    wire N__4533;
    wire N__4530;
    wire N__4527;
    wire N__4526;
    wire N__4523;
    wire N__4522;
    wire N__4519;
    wire N__4516;
    wire N__4515;
    wire N__4514;
    wire N__4511;
    wire N__4506;
    wire N__4503;
    wire N__4500;
    wire N__4491;
    wire N__4488;
    wire N__4485;
    wire N__4482;
    wire N__4479;
    wire N__4476;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4461;
    wire N__4458;
    wire N__4455;
    wire N__4452;
    wire N__4449;
    wire N__4448;
    wire N__4445;
    wire N__4442;
    wire N__4437;
    wire N__4434;
    wire N__4431;
    wire N__4428;
    wire N__4425;
    wire N__4422;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4402;
    wire N__4401;
    wire N__4398;
    wire N__4395;
    wire N__4392;
    wire N__4389;
    wire N__4380;
    wire N__4379;
    wire N__4376;
    wire N__4373;
    wire N__4370;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire N__4355;
    wire N__4350;
    wire N__4347;
    wire N__4344;
    wire N__4341;
    wire N__4338;
    wire N__4335;
    wire N__4332;
    wire N__4329;
    wire N__4326;
    wire N__4323;
    wire N__4320;
    wire N__4317;
    wire N__4314;
    wire N__4311;
    wire N__4308;
    wire N__4305;
    wire N__4302;
    wire N__4299;
    wire N__4298;
    wire N__4295;
    wire N__4292;
    wire N__4287;
    wire N__4284;
    wire N__4281;
    wire N__4278;
    wire N__4275;
    wire N__4274;
    wire N__4271;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4256;
    wire N__4253;
    wire N__4250;
    wire N__4247;
    wire N__4242;
    wire N__4239;
    wire N__4236;
    wire N__4233;
    wire N__4230;
    wire N__4227;
    wire N__4224;
    wire N__4221;
    wire N__4218;
    wire N__4217;
    wire N__4214;
    wire N__4211;
    wire N__4206;
    wire N__4203;
    wire N__4200;
    wire N__4197;
    wire N__4196;
    wire N__4195;
    wire N__4192;
    wire N__4187;
    wire N__4182;
    wire N__4179;
    wire N__4176;
    wire N__4173;
    wire N__4172;
    wire N__4169;
    wire N__4166;
    wire N__4163;
    wire N__4160;
    wire N__4155;
    wire N__4152;
    wire N__4149;
    wire N__4146;
    wire N__4143;
    wire N__4140;
    wire N__4139;
    wire N__4138;
    wire N__4137;
    wire N__4134;
    wire N__4127;
    wire N__4124;
    wire N__4119;
    wire N__4116;
    wire N__4113;
    wire N__4110;
    wire N__4107;
    wire N__4104;
    wire N__4101;
    wire N__4098;
    wire N__4095;
    wire N__4092;
    wire N__4089;
    wire N__4086;
    wire N__4083;
    wire N__4080;
    wire N__4077;
    wire N__4074;
    wire N__4071;
    wire N__4068;
    wire N__4065;
    wire N__4062;
    wire N__4059;
    wire N__4056;
    wire N__4053;
    wire N__4050;
    wire N__4047;
    wire N__4044;
    wire N__4041;
    wire N__4038;
    wire N__4035;
    wire N__4032;
    wire N__4029;
    wire N__4026;
    wire N__4023;
    wire N__4020;
    wire N__4017;
    wire N__4014;
    wire N__4011;
    wire N__4008;
    wire N__4005;
    wire N__4002;
    wire N__3999;
    wire N__3996;
    wire N__3993;
    wire N__3990;
    wire N__3987;
    wire N__3984;
    wire N__3981;
    wire N__3978;
    wire N__3975;
    wire N__3972;
    wire N__3969;
    wire N__3966;
    wire N__3963;
    wire N__3962;
    wire N__3959;
    wire N__3956;
    wire N__3951;
    wire N__3948;
    wire N__3945;
    wire N__3942;
    wire N__3939;
    wire N__3936;
    wire N__3933;
    wire N__3930;
    wire N__3927;
    wire N__3924;
    wire N__3921;
    wire N__3918;
    wire N__3915;
    wire N__3912;
    wire N__3909;
    wire N__3906;
    wire N__3903;
    wire N__3900;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire CLK80_PLL_i_i;
    wire DBRn_c_i_0;
    wire DBRn_c;
    wire DBR_SYNCZ0Z_0;
    wire RAMSPACEn_c;
    wire A_c_18;
    wire A_c_16;
    wire N_848_i;
    wire N_336;
    wire VBENn_c;
    wire \U712_CHIP_RAM.SDRAM_COUNTER18_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_0 ;
    wire \U712_CHIP_RAM.N_371_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0 ;
    wire \U712_CHIP_RAM.N_321 ;
    wire AWEn_c;
    wire \U712_CHIP_RAM.N_371 ;
    wire DBDIR_c;
    wire \U712_CHIP_RAM.N_285_cascade_ ;
    wire \U712_CHIP_RAM.N_309_cascade_ ;
    wire \U712_CHIP_RAM.N_311 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_55_i_a2_0_0_cascade_ ;
    wire \U712_CHIP_RAM.N_212 ;
    wire \U712_CHIP_RAM.N_326_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0_cascade_ ;
    wire A_c_12;
    wire A_c_5;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire TACK_EN_i_ess;
    wire \U712_REG_SM.N_294_cascade_ ;
    wire TSn_c;
    wire REGSPACEn_c;
    wire REG_CYCLEm;
    wire DRDENn_c;
    wire \U712_CHIP_RAM.LATCH_CLK_8_i_0_0_cascade_ ;
    wire \U712_CHIP_RAM.N_368_cascade_ ;
    wire \U712_CHIP_RAM.N_323_cascade_ ;
    wire \U712_CHIP_RAM.N_359_cascade_ ;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_ ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_ ;
    wire A_c_20;
    wire \U712_CHIP_RAM.SDRAM_COUNTER15 ;
    wire \U712_CHIP_RAM.N_330_cascade_ ;
    wire \U712_CHIP_RAM.N_331 ;
    wire \U712_CHIP_RAM.BANK0_9_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ;
    wire BANK0_c;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_0 ;
    wire \U712_CHIP_RAM.N_16 ;
    wire \U712_CHIP_RAM.N_49_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_55_i_a2_0_a2_0_0 ;
    wire A_c_15;
    wire A_c_8;
    wire \U712_CHIP_RAM.N_217 ;
    wire \U712_CHIP_RAM.N_361 ;
    wire \U712_CHIP_RAM.N_217_cascade_ ;
    wire \U712_CHIP_RAM.N_222 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ;
    wire \U712_CHIP_RAM.N_262 ;
    wire \U712_CHIP_RAM.N_354_cascade_ ;
    wire \U712_CHIP_RAM.N_408 ;
    wire \U712_CHIP_RAM.N_408_cascade_ ;
    wire \U712_CHIP_RAM.N_359 ;
    wire \U712_CHIP_RAM.N_305 ;
    wire \U712_CYCLE_TERM.N_236_i_0_en_cascade_ ;
    wire \U712_CYCLE_TERM.N_236_i_0_en_0 ;
    wire \U712_REG_SM.STATE_COUNTc_1_0 ;
    wire DBR_SYNCZ0Z_1;
    wire \U712_REG_SM.N_255 ;
    wire C3_c;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_REG_SM.STATE_COUNT_srsts_i_0_a2_0_0_0 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_1 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_0 ;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.N_264 ;
    wire \U712_REG_SM.N_24 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_2 ;
    wire \U712_CHIP_RAM.N_323 ;
    wire \U712_CHIP_RAM.N_63 ;
    wire LATCH_CLK_c;
    wire \U712_CHIP_RAM.N_363 ;
    wire \U712_CHIP_RAM.N_363_cascade_ ;
    wire \U712_CHIP_RAM.N_369 ;
    wire \U712_CHIP_RAM.N_397 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0 ;
    wire \U712_CHIP_RAM.N_306 ;
    wire bfn_10_6_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.N_49 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.N_352_cascade_ ;
    wire \U712_CHIP_RAM.N_328_cascade_ ;
    wire \U712_CHIP_RAM.un3_DMA_CYCLE_START ;
    wire \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_0 ;
    wire \U712_CHIP_RAM.N_207 ;
    wire \U712_CHIP_RAM.CLK_EN_5_0_a2_1_a2_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0_1 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_370 ;
    wire \U712_CHIP_RAM.N_307 ;
    wire \U712_CHIP_RAM.N_411 ;
    wire \U712_CHIP_RAM.N_403 ;
    wire \U712_CHIP_RAM.N_411_cascade_ ;
    wire \U712_CHIP_RAM.N_308 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.N_352 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_REG_SM.N_232 ;
    wire REG_TACK;
    wire \U712_REG_SM.N_289 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.N_254 ;
    wire \U712_REG_SM.N_254_cascade_ ;
    wire \U712_REG_SM.N_26 ;
    wire C1_c;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire \U712_REG_SM.N_216 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire \U712_REG_SM.N_239 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire ASn_c;
    wire \U712_REG_SM.N_239_0_0 ;
    wire RnW_c;
    wire WRITE_CYCLEm;
    wire N_259;
    wire \U712_CHIP_RAM.N_360 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0_0 ;
    wire \U712_CHIP_RAM.CLK_EN_5_0 ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.N_404 ;
    wire \U712_CHIP_RAM.N_313_2 ;
    wire \U712_CHIP_RAM.N_312_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.N_314 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_cascade_ ;
    wire \U712_CHIP_RAM.N_37 ;
    wire CPU_TACKm;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.N_396 ;
    wire \U712_CHIP_RAM.N_400 ;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire TACK_OUTn;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ;
    wire bfn_11_10_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire C1_c_g;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH5lto2 ;
    wire \U712_CHIP_RAM.REFRESH5lt7 ;
    wire CONSTANT_ONE_NET;
    wire A_c_7;
    wire \U712_CHIP_RAM.N_231_cascade_ ;
    wire A_c_14;
    wire CLK40_PLL_i;
    wire CLK40_PLL_i_i;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_2 ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ;
    wire A_c_3;
    wire A_c_10;
    wire N_180_i;
    wire RESETn_c;
    wire RESETn_c_i;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire CMA_c_3;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1_cascade_ ;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ;
    wire CMA_c_5;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ;
    wire A_c_2;
    wire A_c_9;
    wire CASLn_c;
    wire \U712_BYTE_ENABLE.N_342 ;
    wire \U712_BYTE_ENABLE.N_341_cascade_ ;
    wire N_55_i;
    wire \U712_BYTE_ENABLE.N_320 ;
    wire \U712_BYTE_ENABLE.N_318_cascade_ ;
    wire N_105_i;
    wire CMA_c_2;
    wire \U712_CHIP_RAM.un1_CMA28_0_i ;
    wire A_c_4;
    wire A_c_11;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ;
    wire DMA_CYCLEm;
    wire CASUn_c;
    wire DBENn_c;
    wire N_57_i;
    wire \U712_BYTE_ENABLE.N_339 ;
    wire \U712_BYTE_ENABLE.N_206_i ;
    wire \U712_BYTE_ENABLE.N_316 ;
    wire N_277_i;
    wire LLBE_i_o2_i;
    wire WEn_c;
    wire A_c_17;
    wire CMA_c_8;
    wire A_c_19;
    wire \U712_CHIP_RAM.CMA_5_0_8 ;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire CMA_c_10;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ;
    wire CMA_c_0;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ;
    wire A_c_13;
    wire A_c_6;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ;
    wire DBRn_c_i;
    wire \U712_CHIP_RAM.DMA_AZ0Z20 ;
    wire \INVU712_CHIP_RAM.DMA_A20C_net ;
    wire UMBEn_c;
    wire A_c_1;
    wire SIZ_c_1;
    wire N_276_i;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire RASn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CRCSn_c;
    wire CASn_c;
    wire CPU_CYCLEm;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ;
    wire CMA_c_4;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ;
    wire CMA_c_7;
    wire \U712_CHIP_RAM.CMA_5_sn_N_5_mux ;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNIHMEAZ0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ;
    wire CMA_c_6;
    wire CLK80_PLL;
    wire \U712_CHIP_RAM.un1_CMA28_0_i_0 ;
    wire RAS0n_c;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ;
    wire un1_LDSn_i_0;
    wire DS_ENm;
    wire A_c_0;
    wire SIZ_c_0;
    wire N_87;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire DRA_c_1;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire DRA_c_6;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire C3_c_g;
    wire DRA_c_9;
    wire AGNUS_REV_c;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire _gnd_net_;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ;
    wire DBRn_c_i_0_g;
    wire RESETn_c_i_g;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL_i),
            .REFERENCECLK(N__3921),
            .RESETB(N__7143),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__11587),
            .DIN(N__11586),
            .DOUT(N__11585),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__11587),
            .PADOUT(N__11586),
            .PADIN(N__11585),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7737),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__11578),
            .DIN(N__11577),
            .DOUT(N__11576),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__11578),
            .PADOUT(N__11577),
            .PADIN(N__11576),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__11569),
            .DIN(N__11568),
            .DOUT(N__11567),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__11569),
            .PADOUT(N__11568),
            .PADIN(N__11567),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9540),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__11560),
            .DIN(N__11559),
            .DOUT(N__11558),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__11560),
            .PADOUT(N__11559),
            .PADIN(N__11558),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6183),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__11551),
            .DIN(N__11550),
            .DOUT(N__11549),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__11551),
            .PADOUT(N__11550),
            .PADIN(N__11549),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__11542),
            .DIN(N__11541),
            .DOUT(N__11540),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__11542),
            .PADOUT(N__11541),
            .PADIN(N__11540),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__11533),
            .DIN(N__11532),
            .DOUT(N__11531),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__11533),
            .PADOUT(N__11532),
            .PADIN(N__11531),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__11524),
            .DIN(N__11523),
            .DOUT(N__11522),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__11524),
            .PADOUT(N__11523),
            .PADIN(N__11522),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__11515),
            .DIN(N__11514),
            .DOUT(N__11513),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__11515),
            .PADOUT(N__11514),
            .PADIN(N__11513),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__11506),
            .DIN(N__11505),
            .DOUT(N__11504),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__11506),
            .PADOUT(N__11505),
            .PADIN(N__11504),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__11497),
            .DIN(N__11496),
            .DOUT(N__11495),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__11497),
            .PADOUT(N__11496),
            .PADIN(N__11495),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9114),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__11488),
            .DIN(N__11487),
            .DOUT(N__11486),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__11488),
            .PADOUT(N__11487),
            .PADIN(N__11486),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8253),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__11479),
            .DIN(N__11478),
            .DOUT(N__11477),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__11479),
            .PADOUT(N__11478),
            .PADIN(N__11477),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMENn_obuf_iopad (
            .OE(N__11470),
            .DIN(N__11469),
            .DOUT(N__11468),
            .PACKAGEPIN(RAMENn));
    defparam RAMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMENn_obuf_preio (
            .PADOEN(N__11470),
            .PADOUT(N__11469),
            .PADIN(N__11468),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4379),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__11461),
            .DIN(N__11460),
            .DOUT(N__11459),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__11461),
            .PADOUT(N__11460),
            .PADIN(N__11459),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__11452),
            .DIN(N__11451),
            .DOUT(N__11450),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__11452),
            .PADOUT(N__11451),
            .PADIN(N__11450),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__11443),
            .DIN(N__11442),
            .DOUT(N__11441),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__11443),
            .PADOUT(N__11442),
            .PADIN(N__11441),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4014),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__11434),
            .DIN(N__11433),
            .DOUT(N__11432),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__11434),
            .PADOUT(N__11433),
            .PADIN(N__11432),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__11425),
            .DIN(N__11424),
            .DOUT(N__11423),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__11425),
            .PADOUT(N__11424),
            .PADIN(N__11423),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__11416),
            .DIN(N__11415),
            .DOUT(N__11414),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__11416),
            .PADOUT(N__11415),
            .PADIN(N__11414),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8727),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__11407),
            .DIN(N__11406),
            .DOUT(N__11405),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__11407),
            .PADOUT(N__11406),
            .PADIN(N__11405),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__11398),
            .DIN(N__11397),
            .DOUT(N__11396),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__11398),
            .PADOUT(N__11397),
            .PADIN(N__11396),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8319),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__11389),
            .DIN(N__11388),
            .DOUT(N__11387),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__11389),
            .PADOUT(N__11388),
            .PADIN(N__11387),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__11380),
            .DIN(N__11379),
            .DOUT(N__11378),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__11380),
            .PADOUT(N__11379),
            .PADIN(N__11378),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8241),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__11371),
            .DIN(N__11370),
            .DOUT(N__11369),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__11371),
            .PADOUT(N__11370),
            .PADIN(N__11369),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__11362),
            .DIN(N__11361),
            .DOUT(N__11360),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__11362),
            .PADOUT(N__11361),
            .PADIN(N__11360),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__11353),
            .DIN(N__11352),
            .DOUT(N__11351),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__11353),
            .PADOUT(N__11352),
            .PADIN(N__11351),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__11344),
            .DIN(N__11343),
            .DOUT(N__11342),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__11344),
            .PADOUT(N__11343),
            .PADIN(N__11342),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__11335),
            .DIN(N__11334),
            .DOUT(N__11333),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__11335),
            .PADOUT(N__11334),
            .PADIN(N__11333),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_EN_obuf_iopad (
            .OE(N__11326),
            .DIN(N__11325),
            .DOUT(N__11324),
            .PACKAGEPIN(DMA_LATCH_EN));
    defparam DMA_LATCH_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_EN_obuf_preio (
            .PADOEN(N__11326),
            .PADOUT(N__11325),
            .PADIN(N__11324),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4026),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__11317),
            .DIN(N__11316),
            .DOUT(N__11315),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__11317),
            .PADOUT(N__11316),
            .PADIN(N__11315),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__11308),
            .DIN(N__11307),
            .DOUT(N__11306),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__11308),
            .PADOUT(N__11307),
            .PADIN(N__11306),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__11299),
            .DIN(N__11298),
            .DOUT(N__11297),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__11299),
            .PADOUT(N__11298),
            .PADIN(N__11297),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__11290),
            .DIN(N__11289),
            .DOUT(N__11288),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__11290),
            .PADOUT(N__11289),
            .PADIN(N__11288),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__11281),
            .DIN(N__11280),
            .DOUT(N__11279),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__11281),
            .PADOUT(N__11280),
            .PADIN(N__11279),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__11272),
            .DIN(N__11271),
            .DOUT(N__11270),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__11272),
            .PADOUT(N__11271),
            .PADIN(N__11270),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5088),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__11263),
            .DIN(N__11262),
            .DOUT(N__11261),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__11263),
            .PADOUT(N__11262),
            .PADIN(N__11261),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9900),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__11254),
            .DIN(N__11253),
            .DOUT(N__11252),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__11254),
            .PADOUT(N__11253),
            .PADIN(N__11252),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7029),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__11245),
            .DIN(N__11244),
            .DOUT(N__11243),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__11245),
            .PADOUT(N__11244),
            .PADIN(N__11243),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__11236),
            .DIN(N__11235),
            .DOUT(N__11234),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__11236),
            .PADOUT(N__11235),
            .PADIN(N__11234),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8379),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__11227),
            .DIN(N__11226),
            .DOUT(N__11225),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__11227),
            .PADOUT(N__11226),
            .PADIN(N__11225),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__11218),
            .DIN(N__11217),
            .DOUT(N__11216),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__11218),
            .PADOUT(N__11217),
            .PADIN(N__11216),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4461),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__11209),
            .DIN(N__11208),
            .DOUT(N__11207),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__11209),
            .PADOUT(N__11208),
            .PADIN(N__11207),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7025),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__11200),
            .DIN(N__11199),
            .DOUT(N__11198),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__11200),
            .PADOUT(N__11199),
            .PADIN(N__11198),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3999),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__11191),
            .DIN(N__11190),
            .DOUT(N__11189),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__11191),
            .PADOUT(N__11190),
            .PADIN(N__11189),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__11182),
            .DIN(N__11181),
            .DOUT(N__11180),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__11182),
            .PADOUT(N__11181),
            .PADIN(N__11180),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6342),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__11173),
            .DIN(N__11172),
            .DOUT(N__11171),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__11173),
            .PADOUT(N__11172),
            .PADIN(N__11171),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7236),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__11164),
            .DIN(N__11163),
            .DOUT(N__11162),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__11164),
            .PADOUT(N__11163),
            .PADIN(N__11162),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__11155),
            .DIN(N__11154),
            .DOUT(N__11153),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__11155),
            .PADOUT(N__11154),
            .PADIN(N__11153),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__11146),
            .DIN(N__11145),
            .DOUT(N__11144),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__11146),
            .PADOUT(N__11145),
            .PADIN(N__11144),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__11137),
            .DIN(N__11136),
            .DOUT(N__11135),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__11137),
            .PADOUT(N__11136),
            .PADIN(N__11135),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__11128),
            .DIN(N__11127),
            .DOUT(N__11126),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__11128),
            .PADOUT(N__11127),
            .PADIN(N__11126),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8031),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__11119),
            .DIN(N__11118),
            .DOUT(N__11117),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__11119),
            .PADOUT(N__11118),
            .PADIN(N__11117),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__11110),
            .DIN(N__11109),
            .DOUT(N__11108),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__11110),
            .PADOUT(N__11109),
            .PADIN(N__11108),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7018),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__11101),
            .DIN(N__11100),
            .DOUT(N__11099),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__11101),
            .PADOUT(N__11100),
            .PADIN(N__11099),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9135),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__11092),
            .DIN(N__11091),
            .DOUT(N__11090),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__11092),
            .PADOUT(N__11091),
            .PADIN(N__11090),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4380),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__11083),
            .DIN(N__11082),
            .DOUT(N__11081),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__11083),
            .PADOUT(N__11082),
            .PADIN(N__11081),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7467),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__11074),
            .DIN(N__11073),
            .DOUT(N__11072),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__11074),
            .PADOUT(N__11073),
            .PADIN(N__11072),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8124),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__11065),
            .DIN(N__11064),
            .DOUT(N__11063),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__11065),
            .PADOUT(N__11064),
            .PADIN(N__11063),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6338),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__11056),
            .DIN(N__11055),
            .DOUT(N__11054),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__11056),
            .PADOUT(N__11055),
            .PADIN(N__11054),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__11047),
            .DIN(N__11046),
            .DOUT(N__11045),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__11047),
            .PADOUT(N__11046),
            .PADIN(N__11045),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__11038),
            .DIN(N__11037),
            .DOUT(N__11036),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__11038),
            .PADOUT(N__11037),
            .PADIN(N__11036),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7680),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__11029),
            .DIN(N__11028),
            .DOUT(N__11027),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__11029),
            .PADOUT(N__11028),
            .PADIN(N__11027),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8226),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__11020),
            .DIN(N__11019),
            .DOUT(N__11018),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__11020),
            .PADOUT(N__11019),
            .PADIN(N__11018),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4182),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__11011),
            .DIN(N__11010),
            .DOUT(N__11009),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__11011),
            .PADOUT(N__11010),
            .PADIN(N__11009),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8001),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__11002),
            .DIN(N__11001),
            .DOUT(N__11000),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__11002),
            .PADOUT(N__11001),
            .PADIN(N__11000),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__10993),
            .DIN(N__10992),
            .DOUT(N__10991),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__10993),
            .PADOUT(N__10992),
            .PADIN(N__10991),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__10984),
            .DIN(N__10983),
            .DOUT(N__10982),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__10984),
            .PADOUT(N__10983),
            .PADIN(N__10982),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__10975),
            .DIN(N__10974),
            .DOUT(N__10973),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__10975),
            .PADOUT(N__10974),
            .PADIN(N__10973),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__10966),
            .DIN(N__10965),
            .DOUT(N__10964),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__10966),
            .PADOUT(N__10965),
            .PADIN(N__10964),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7212),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__10957),
            .DIN(N__10956),
            .DOUT(N__10955),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__10957),
            .PADOUT(N__10956),
            .PADIN(N__10955),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8457),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__10948),
            .DIN(N__10947),
            .DOUT(N__10946),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__10948),
            .PADOUT(N__10947),
            .PADIN(N__10946),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__10939),
            .DIN(N__10938),
            .DOUT(N__10937),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__10939),
            .PADOUT(N__10938),
            .PADIN(N__10937),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7398),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__10930),
            .DIN(N__10929),
            .DOUT(N__10928),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__10930),
            .PADOUT(N__10929),
            .PADIN(N__10928),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4044),
            .DIN0(),
            .DOUT0(N__6567),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__10921),
            .DIN(N__10920),
            .DOUT(N__10919),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__10921),
            .PADOUT(N__10920),
            .PADIN(N__10919),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7977),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__10912),
            .DIN(N__10911),
            .DOUT(N__10910),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__10912),
            .PADOUT(N__10911),
            .PADIN(N__10910),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__10903),
            .DIN(N__10902),
            .DOUT(N__10901),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__10903),
            .PADOUT(N__10902),
            .PADIN(N__10901),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__10894),
            .DIN(N__10893),
            .DOUT(N__10892),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__10894),
            .PADOUT(N__10893),
            .PADIN(N__10892),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8187),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__10885),
            .DIN(N__10884),
            .DOUT(N__10883),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__10885),
            .PADOUT(N__10884),
            .PADIN(N__10883),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__10876),
            .DIN(N__10875),
            .DOUT(N__10874),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__10876),
            .PADOUT(N__10875),
            .PADIN(N__10874),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__10867),
            .DIN(N__10866),
            .DOUT(N__10865),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__10867),
            .PADOUT(N__10866),
            .PADIN(N__10865),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__10858),
            .DIN(N__10857),
            .DOUT(N__10856),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__10858),
            .PADOUT(N__10857),
            .PADIN(N__10856),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__10849),
            .DIN(N__10848),
            .DOUT(N__10847),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__10849),
            .PADOUT(N__10848),
            .PADIN(N__10847),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7632),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__10840),
            .DIN(N__10839),
            .DOUT(N__10838),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__10840),
            .PADOUT(N__10839),
            .PADIN(N__10838),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9660),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__10831),
            .DIN(N__10830),
            .DOUT(N__10829),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__10831),
            .PADOUT(N__10830),
            .PADIN(N__10829),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8610),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__10822),
            .DIN(N__10821),
            .DOUT(N__10820),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__10822),
            .PADOUT(N__10821),
            .PADIN(N__10820),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6093),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__10813),
            .DIN(N__10812),
            .DOUT(N__10811),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__10813),
            .PADOUT(N__10812),
            .PADIN(N__10811),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__10804),
            .DIN(N__10803),
            .DOUT(N__10802),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__10804),
            .PADOUT(N__10803),
            .PADIN(N__10802),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__10795),
            .DIN(N__10794),
            .DOUT(N__10793),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__10795),
            .PADOUT(N__10794),
            .PADIN(N__10793),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8988),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__10786),
            .DIN(N__10785),
            .DOUT(N__10784),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__10786),
            .PADOUT(N__10785),
            .PADIN(N__10784),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2625 (
            .O(N__10767),
            .I(N__10763));
    CascadeMux I__2624 (
            .O(N__10766),
            .I(N__10760));
    LocalMux I__2623 (
            .O(N__10763),
            .I(N__10757));
    InMux I__2622 (
            .O(N__10760),
            .I(N__10754));
    Span4Mux_h I__2621 (
            .O(N__10757),
            .I(N__10748));
    LocalMux I__2620 (
            .O(N__10754),
            .I(N__10748));
    InMux I__2619 (
            .O(N__10753),
            .I(N__10745));
    Span4Mux_v I__2618 (
            .O(N__10748),
            .I(N__10741));
    LocalMux I__2617 (
            .O(N__10745),
            .I(N__10738));
    InMux I__2616 (
            .O(N__10744),
            .I(N__10735));
    Sp12to4 I__2615 (
            .O(N__10741),
            .I(N__10732));
    Sp12to4 I__2614 (
            .O(N__10738),
            .I(N__10727));
    LocalMux I__2613 (
            .O(N__10735),
            .I(N__10727));
    Span12Mux_h I__2612 (
            .O(N__10732),
            .I(N__10724));
    Span12Mux_v I__2611 (
            .O(N__10727),
            .I(N__10721));
    Span12Mux_v I__2610 (
            .O(N__10724),
            .I(N__10718));
    Span12Mux_v I__2609 (
            .O(N__10721),
            .I(N__10715));
    Odrv12 I__2608 (
            .O(N__10718),
            .I(DRA_c_9));
    Odrv12 I__2607 (
            .O(N__10715),
            .I(DRA_c_9));
    InMux I__2606 (
            .O(N__10710),
            .I(N__10704));
    CascadeMux I__2605 (
            .O(N__10709),
            .I(N__10699));
    CascadeMux I__2604 (
            .O(N__10708),
            .I(N__10689));
    CascadeMux I__2603 (
            .O(N__10707),
            .I(N__10685));
    LocalMux I__2602 (
            .O(N__10704),
            .I(N__10681));
    InMux I__2601 (
            .O(N__10703),
            .I(N__10676));
    InMux I__2600 (
            .O(N__10702),
            .I(N__10665));
    InMux I__2599 (
            .O(N__10699),
            .I(N__10665));
    InMux I__2598 (
            .O(N__10698),
            .I(N__10665));
    InMux I__2597 (
            .O(N__10697),
            .I(N__10665));
    InMux I__2596 (
            .O(N__10696),
            .I(N__10665));
    CascadeMux I__2595 (
            .O(N__10695),
            .I(N__10662));
    CascadeMux I__2594 (
            .O(N__10694),
            .I(N__10657));
    CascadeMux I__2593 (
            .O(N__10693),
            .I(N__10654));
    InMux I__2592 (
            .O(N__10692),
            .I(N__10646));
    InMux I__2591 (
            .O(N__10689),
            .I(N__10646));
    InMux I__2590 (
            .O(N__10688),
            .I(N__10646));
    InMux I__2589 (
            .O(N__10685),
            .I(N__10641));
    InMux I__2588 (
            .O(N__10684),
            .I(N__10641));
    Span4Mux_v I__2587 (
            .O(N__10681),
            .I(N__10638));
    InMux I__2586 (
            .O(N__10680),
            .I(N__10635));
    InMux I__2585 (
            .O(N__10679),
            .I(N__10632));
    LocalMux I__2584 (
            .O(N__10676),
            .I(N__10627));
    LocalMux I__2583 (
            .O(N__10665),
            .I(N__10627));
    InMux I__2582 (
            .O(N__10662),
            .I(N__10622));
    InMux I__2581 (
            .O(N__10661),
            .I(N__10622));
    InMux I__2580 (
            .O(N__10660),
            .I(N__10612));
    InMux I__2579 (
            .O(N__10657),
            .I(N__10612));
    InMux I__2578 (
            .O(N__10654),
            .I(N__10612));
    InMux I__2577 (
            .O(N__10653),
            .I(N__10612));
    LocalMux I__2576 (
            .O(N__10646),
            .I(N__10607));
    LocalMux I__2575 (
            .O(N__10641),
            .I(N__10607));
    Span4Mux_h I__2574 (
            .O(N__10638),
            .I(N__10596));
    LocalMux I__2573 (
            .O(N__10635),
            .I(N__10596));
    LocalMux I__2572 (
            .O(N__10632),
            .I(N__10596));
    Span4Mux_v I__2571 (
            .O(N__10627),
            .I(N__10596));
    LocalMux I__2570 (
            .O(N__10622),
            .I(N__10596));
    InMux I__2569 (
            .O(N__10621),
            .I(N__10593));
    LocalMux I__2568 (
            .O(N__10612),
            .I(N__10590));
    Span4Mux_v I__2567 (
            .O(N__10607),
            .I(N__10583));
    Span4Mux_h I__2566 (
            .O(N__10596),
            .I(N__10583));
    LocalMux I__2565 (
            .O(N__10593),
            .I(N__10583));
    Span4Mux_v I__2564 (
            .O(N__10590),
            .I(N__10580));
    Span4Mux_h I__2563 (
            .O(N__10583),
            .I(N__10577));
    Span4Mux_v I__2562 (
            .O(N__10580),
            .I(N__10574));
    Span4Mux_h I__2561 (
            .O(N__10577),
            .I(N__10571));
    Sp12to4 I__2560 (
            .O(N__10574),
            .I(N__10568));
    Sp12to4 I__2559 (
            .O(N__10571),
            .I(N__10565));
    Span12Mux_h I__2558 (
            .O(N__10568),
            .I(N__10562));
    Span12Mux_v I__2557 (
            .O(N__10565),
            .I(N__10559));
    Odrv12 I__2556 (
            .O(N__10562),
            .I(AGNUS_REV_c));
    Odrv12 I__2555 (
            .O(N__10559),
            .I(AGNUS_REV_c));
    InMux I__2554 (
            .O(N__10554),
            .I(N__10550));
    InMux I__2553 (
            .O(N__10553),
            .I(N__10547));
    LocalMux I__2552 (
            .O(N__10550),
            .I(N__10541));
    LocalMux I__2551 (
            .O(N__10547),
            .I(N__10541));
    InMux I__2550 (
            .O(N__10546),
            .I(N__10538));
    Span4Mux_v I__2549 (
            .O(N__10541),
            .I(N__10532));
    LocalMux I__2548 (
            .O(N__10538),
            .I(N__10532));
    InMux I__2547 (
            .O(N__10537),
            .I(N__10529));
    Sp12to4 I__2546 (
            .O(N__10532),
            .I(N__10524));
    LocalMux I__2545 (
            .O(N__10529),
            .I(N__10524));
    Odrv12 I__2544 (
            .O(N__10524),
            .I(DRA_c_8));
    InMux I__2543 (
            .O(N__10521),
            .I(N__10518));
    LocalMux I__2542 (
            .O(N__10518),
            .I(N__10515));
    Span4Mux_h I__2541 (
            .O(N__10515),
            .I(N__10512));
    Odrv4 I__2540 (
            .O(N__10512),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    CEMux I__2539 (
            .O(N__10509),
            .I(N__10485));
    CEMux I__2538 (
            .O(N__10508),
            .I(N__10485));
    CEMux I__2537 (
            .O(N__10507),
            .I(N__10485));
    CEMux I__2536 (
            .O(N__10506),
            .I(N__10485));
    CEMux I__2535 (
            .O(N__10505),
            .I(N__10485));
    CEMux I__2534 (
            .O(N__10504),
            .I(N__10485));
    CEMux I__2533 (
            .O(N__10503),
            .I(N__10485));
    CEMux I__2532 (
            .O(N__10502),
            .I(N__10485));
    GlobalMux I__2531 (
            .O(N__10485),
            .I(N__10482));
    gio2CtrlBuf I__2530 (
            .O(N__10482),
            .I(DBRn_c_i_0_g));
    InMux I__2529 (
            .O(N__10479),
            .I(N__10470));
    InMux I__2528 (
            .O(N__10478),
            .I(N__10465));
    InMux I__2527 (
            .O(N__10477),
            .I(N__10465));
    InMux I__2526 (
            .O(N__10476),
            .I(N__10462));
    InMux I__2525 (
            .O(N__10475),
            .I(N__10459));
    InMux I__2524 (
            .O(N__10474),
            .I(N__10456));
    InMux I__2523 (
            .O(N__10473),
            .I(N__10453));
    LocalMux I__2522 (
            .O(N__10470),
            .I(N__10448));
    LocalMux I__2521 (
            .O(N__10465),
            .I(N__10439));
    LocalMux I__2520 (
            .O(N__10462),
            .I(N__10431));
    LocalMux I__2519 (
            .O(N__10459),
            .I(N__10417));
    LocalMux I__2518 (
            .O(N__10456),
            .I(N__10406));
    LocalMux I__2517 (
            .O(N__10453),
            .I(N__10395));
    SRMux I__2516 (
            .O(N__10452),
            .I(N__10299));
    SRMux I__2515 (
            .O(N__10451),
            .I(N__10299));
    Glb2LocalMux I__2514 (
            .O(N__10448),
            .I(N__10299));
    SRMux I__2513 (
            .O(N__10447),
            .I(N__10299));
    SRMux I__2512 (
            .O(N__10446),
            .I(N__10299));
    SRMux I__2511 (
            .O(N__10445),
            .I(N__10299));
    SRMux I__2510 (
            .O(N__10444),
            .I(N__10299));
    SRMux I__2509 (
            .O(N__10443),
            .I(N__10299));
    SRMux I__2508 (
            .O(N__10442),
            .I(N__10299));
    Glb2LocalMux I__2507 (
            .O(N__10439),
            .I(N__10299));
    SRMux I__2506 (
            .O(N__10438),
            .I(N__10299));
    SRMux I__2505 (
            .O(N__10437),
            .I(N__10299));
    SRMux I__2504 (
            .O(N__10436),
            .I(N__10299));
    SRMux I__2503 (
            .O(N__10435),
            .I(N__10299));
    SRMux I__2502 (
            .O(N__10434),
            .I(N__10299));
    Glb2LocalMux I__2501 (
            .O(N__10431),
            .I(N__10299));
    SRMux I__2500 (
            .O(N__10430),
            .I(N__10299));
    SRMux I__2499 (
            .O(N__10429),
            .I(N__10299));
    SRMux I__2498 (
            .O(N__10428),
            .I(N__10299));
    SRMux I__2497 (
            .O(N__10427),
            .I(N__10299));
    SRMux I__2496 (
            .O(N__10426),
            .I(N__10299));
    SRMux I__2495 (
            .O(N__10425),
            .I(N__10299));
    SRMux I__2494 (
            .O(N__10424),
            .I(N__10299));
    SRMux I__2493 (
            .O(N__10423),
            .I(N__10299));
    SRMux I__2492 (
            .O(N__10422),
            .I(N__10299));
    SRMux I__2491 (
            .O(N__10421),
            .I(N__10299));
    SRMux I__2490 (
            .O(N__10420),
            .I(N__10299));
    Glb2LocalMux I__2489 (
            .O(N__10417),
            .I(N__10299));
    SRMux I__2488 (
            .O(N__10416),
            .I(N__10299));
    SRMux I__2487 (
            .O(N__10415),
            .I(N__10299));
    SRMux I__2486 (
            .O(N__10414),
            .I(N__10299));
    SRMux I__2485 (
            .O(N__10413),
            .I(N__10299));
    SRMux I__2484 (
            .O(N__10412),
            .I(N__10299));
    SRMux I__2483 (
            .O(N__10411),
            .I(N__10299));
    SRMux I__2482 (
            .O(N__10410),
            .I(N__10299));
    SRMux I__2481 (
            .O(N__10409),
            .I(N__10299));
    Glb2LocalMux I__2480 (
            .O(N__10406),
            .I(N__10299));
    SRMux I__2479 (
            .O(N__10405),
            .I(N__10299));
    SRMux I__2478 (
            .O(N__10404),
            .I(N__10299));
    SRMux I__2477 (
            .O(N__10403),
            .I(N__10299));
    SRMux I__2476 (
            .O(N__10402),
            .I(N__10299));
    SRMux I__2475 (
            .O(N__10401),
            .I(N__10299));
    SRMux I__2474 (
            .O(N__10400),
            .I(N__10299));
    SRMux I__2473 (
            .O(N__10399),
            .I(N__10299));
    SRMux I__2472 (
            .O(N__10398),
            .I(N__10299));
    Glb2LocalMux I__2471 (
            .O(N__10395),
            .I(N__10299));
    SRMux I__2470 (
            .O(N__10394),
            .I(N__10299));
    GlobalMux I__2469 (
            .O(N__10299),
            .I(N__10296));
    gio2CtrlBuf I__2468 (
            .O(N__10296),
            .I(RESETn_c_i_g));
    InMux I__2467 (
            .O(N__10293),
            .I(N__10290));
    LocalMux I__2466 (
            .O(N__10290),
            .I(N__10287));
    Odrv12 I__2465 (
            .O(N__10287),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__2464 (
            .O(N__10284),
            .I(N__10278));
    InMux I__2463 (
            .O(N__10283),
            .I(N__10278));
    LocalMux I__2462 (
            .O(N__10278),
            .I(N__10273));
    InMux I__2461 (
            .O(N__10277),
            .I(N__10268));
    InMux I__2460 (
            .O(N__10276),
            .I(N__10268));
    Span4Mux_h I__2459 (
            .O(N__10273),
            .I(N__10263));
    LocalMux I__2458 (
            .O(N__10268),
            .I(N__10263));
    Sp12to4 I__2457 (
            .O(N__10263),
            .I(N__10260));
    Span12Mux_v I__2456 (
            .O(N__10260),
            .I(N__10257));
    Odrv12 I__2455 (
            .O(N__10257),
            .I(DRA_c_3));
    InMux I__2454 (
            .O(N__10254),
            .I(N__10251));
    LocalMux I__2453 (
            .O(N__10251),
            .I(N__10248));
    Odrv4 I__2452 (
            .O(N__10248),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__2451 (
            .O(N__10245),
            .I(N__10239));
    InMux I__2450 (
            .O(N__10244),
            .I(N__10239));
    LocalMux I__2449 (
            .O(N__10239),
            .I(N__10236));
    Span4Mux_v I__2448 (
            .O(N__10236),
            .I(N__10231));
    InMux I__2447 (
            .O(N__10235),
            .I(N__10228));
    InMux I__2446 (
            .O(N__10234),
            .I(N__10225));
    Sp12to4 I__2445 (
            .O(N__10231),
            .I(N__10220));
    LocalMux I__2444 (
            .O(N__10228),
            .I(N__10220));
    LocalMux I__2443 (
            .O(N__10225),
            .I(N__10217));
    Span12Mux_h I__2442 (
            .O(N__10220),
            .I(N__10214));
    Sp12to4 I__2441 (
            .O(N__10217),
            .I(N__10211));
    Span12Mux_v I__2440 (
            .O(N__10214),
            .I(N__10208));
    Span12Mux_v I__2439 (
            .O(N__10211),
            .I(N__10205));
    Odrv12 I__2438 (
            .O(N__10208),
            .I(DRA_c_1));
    Odrv12 I__2437 (
            .O(N__10205),
            .I(DRA_c_1));
    InMux I__2436 (
            .O(N__10200),
            .I(N__10196));
    InMux I__2435 (
            .O(N__10199),
            .I(N__10193));
    LocalMux I__2434 (
            .O(N__10196),
            .I(N__10188));
    LocalMux I__2433 (
            .O(N__10193),
            .I(N__10188));
    Span4Mux_h I__2432 (
            .O(N__10188),
            .I(N__10185));
    Sp12to4 I__2431 (
            .O(N__10185),
            .I(N__10182));
    Span12Mux_v I__2430 (
            .O(N__10182),
            .I(N__10179));
    Odrv12 I__2429 (
            .O(N__10179),
            .I(DRA_c_0));
    InMux I__2428 (
            .O(N__10176),
            .I(N__10173));
    LocalMux I__2427 (
            .O(N__10173),
            .I(N__10170));
    Span4Mux_v I__2426 (
            .O(N__10170),
            .I(N__10167));
    Sp12to4 I__2425 (
            .O(N__10167),
            .I(N__10164));
    Odrv12 I__2424 (
            .O(N__10164),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    InMux I__2423 (
            .O(N__10161),
            .I(N__10158));
    LocalMux I__2422 (
            .O(N__10158),
            .I(N__10155));
    Span4Mux_h I__2421 (
            .O(N__10155),
            .I(N__10152));
    Span4Mux_h I__2420 (
            .O(N__10152),
            .I(N__10149));
    Odrv4 I__2419 (
            .O(N__10149),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__2418 (
            .O(N__10146),
            .I(N__10143));
    LocalMux I__2417 (
            .O(N__10143),
            .I(N__10140));
    Span4Mux_v I__2416 (
            .O(N__10140),
            .I(N__10137));
    Odrv4 I__2415 (
            .O(N__10137),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__2414 (
            .O(N__10134),
            .I(N__10128));
    InMux I__2413 (
            .O(N__10133),
            .I(N__10125));
    InMux I__2412 (
            .O(N__10132),
            .I(N__10122));
    InMux I__2411 (
            .O(N__10131),
            .I(N__10119));
    LocalMux I__2410 (
            .O(N__10128),
            .I(N__10110));
    LocalMux I__2409 (
            .O(N__10125),
            .I(N__10110));
    LocalMux I__2408 (
            .O(N__10122),
            .I(N__10110));
    LocalMux I__2407 (
            .O(N__10119),
            .I(N__10110));
    Span4Mux_v I__2406 (
            .O(N__10110),
            .I(N__10107));
    Sp12to4 I__2405 (
            .O(N__10107),
            .I(N__10104));
    Span12Mux_h I__2404 (
            .O(N__10104),
            .I(N__10101));
    Odrv12 I__2403 (
            .O(N__10101),
            .I(DRA_c_7));
    InMux I__2402 (
            .O(N__10098),
            .I(N__10095));
    LocalMux I__2401 (
            .O(N__10095),
            .I(N__10092));
    Span4Mux_h I__2400 (
            .O(N__10092),
            .I(N__10089));
    Odrv4 I__2399 (
            .O(N__10089),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__2398 (
            .O(N__10086),
            .I(N__10079));
    InMux I__2397 (
            .O(N__10085),
            .I(N__10079));
    InMux I__2396 (
            .O(N__10084),
            .I(N__10076));
    LocalMux I__2395 (
            .O(N__10079),
            .I(N__10072));
    LocalMux I__2394 (
            .O(N__10076),
            .I(N__10069));
    InMux I__2393 (
            .O(N__10075),
            .I(N__10066));
    Span4Mux_v I__2392 (
            .O(N__10072),
            .I(N__10063));
    Span4Mux_h I__2391 (
            .O(N__10069),
            .I(N__10058));
    LocalMux I__2390 (
            .O(N__10066),
            .I(N__10058));
    Span4Mux_v I__2389 (
            .O(N__10063),
            .I(N__10055));
    Span4Mux_v I__2388 (
            .O(N__10058),
            .I(N__10052));
    Span4Mux_h I__2387 (
            .O(N__10055),
            .I(N__10049));
    Span4Mux_v I__2386 (
            .O(N__10052),
            .I(N__10046));
    Sp12to4 I__2385 (
            .O(N__10049),
            .I(N__10041));
    Sp12to4 I__2384 (
            .O(N__10046),
            .I(N__10041));
    Odrv12 I__2383 (
            .O(N__10041),
            .I(DRA_c_4));
    InMux I__2382 (
            .O(N__10038),
            .I(N__10035));
    LocalMux I__2381 (
            .O(N__10035),
            .I(N__10032));
    Span4Mux_v I__2380 (
            .O(N__10032),
            .I(N__10029));
    Odrv4 I__2379 (
            .O(N__10029),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__2378 (
            .O(N__10026),
            .I(N__10023));
    LocalMux I__2377 (
            .O(N__10023),
            .I(N__10017));
    InMux I__2376 (
            .O(N__10022),
            .I(N__10014));
    InMux I__2375 (
            .O(N__10021),
            .I(N__10011));
    InMux I__2374 (
            .O(N__10020),
            .I(N__10008));
    Span4Mux_v I__2373 (
            .O(N__10017),
            .I(N__10005));
    LocalMux I__2372 (
            .O(N__10014),
            .I(N__9998));
    LocalMux I__2371 (
            .O(N__10011),
            .I(N__9998));
    LocalMux I__2370 (
            .O(N__10008),
            .I(N__9998));
    Span4Mux_v I__2369 (
            .O(N__10005),
            .I(N__9995));
    Sp12to4 I__2368 (
            .O(N__9998),
            .I(N__9992));
    Sp12to4 I__2367 (
            .O(N__9995),
            .I(N__9987));
    Span12Mux_v I__2366 (
            .O(N__9992),
            .I(N__9987));
    Odrv12 I__2365 (
            .O(N__9987),
            .I(DRA_c_6));
    InMux I__2364 (
            .O(N__9984),
            .I(N__9981));
    LocalMux I__2363 (
            .O(N__9981),
            .I(N__9975));
    InMux I__2362 (
            .O(N__9980),
            .I(N__9972));
    InMux I__2361 (
            .O(N__9979),
            .I(N__9967));
    InMux I__2360 (
            .O(N__9978),
            .I(N__9967));
    Span4Mux_h I__2359 (
            .O(N__9975),
            .I(N__9962));
    LocalMux I__2358 (
            .O(N__9972),
            .I(N__9962));
    LocalMux I__2357 (
            .O(N__9967),
            .I(N__9957));
    Sp12to4 I__2356 (
            .O(N__9962),
            .I(N__9957));
    Span12Mux_v I__2355 (
            .O(N__9957),
            .I(N__9954));
    Odrv12 I__2354 (
            .O(N__9954),
            .I(DRA_c_5));
    InMux I__2353 (
            .O(N__9951),
            .I(N__9945));
    InMux I__2352 (
            .O(N__9950),
            .I(N__9945));
    LocalMux I__2351 (
            .O(N__9945),
            .I(N__9942));
    Span12Mux_v I__2350 (
            .O(N__9942),
            .I(N__9939));
    Odrv12 I__2349 (
            .O(N__9939),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    ClkMux I__2348 (
            .O(N__9936),
            .I(N__9924));
    ClkMux I__2347 (
            .O(N__9935),
            .I(N__9924));
    ClkMux I__2346 (
            .O(N__9934),
            .I(N__9924));
    ClkMux I__2345 (
            .O(N__9933),
            .I(N__9924));
    GlobalMux I__2344 (
            .O(N__9924),
            .I(N__9921));
    gio2CtrlBuf I__2343 (
            .O(N__9921),
            .I(C3_c_g));
    InMux I__2342 (
            .O(N__9918),
            .I(N__9915));
    LocalMux I__2341 (
            .O(N__9915),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__2340 (
            .O(N__9912),
            .I(N__9909));
    LocalMux I__2339 (
            .O(N__9909),
            .I(N__9906));
    Span4Mux_h I__2338 (
            .O(N__9906),
            .I(N__9903));
    Odrv4 I__2337 (
            .O(N__9903),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    IoInMux I__2336 (
            .O(N__9900),
            .I(N__9897));
    LocalMux I__2335 (
            .O(N__9897),
            .I(N__9894));
    Span4Mux_s3_v I__2334 (
            .O(N__9894),
            .I(N__9891));
    Span4Mux_h I__2333 (
            .O(N__9891),
            .I(N__9888));
    Span4Mux_v I__2332 (
            .O(N__9888),
            .I(N__9885));
    Odrv4 I__2331 (
            .O(N__9885),
            .I(un1_LDSn_i_0));
    InMux I__2330 (
            .O(N__9882),
            .I(N__9878));
    InMux I__2329 (
            .O(N__9881),
            .I(N__9875));
    LocalMux I__2328 (
            .O(N__9878),
            .I(N__9870));
    LocalMux I__2327 (
            .O(N__9875),
            .I(N__9870));
    Span4Mux_v I__2326 (
            .O(N__9870),
            .I(N__9867));
    Span4Mux_h I__2325 (
            .O(N__9867),
            .I(N__9864));
    Span4Mux_v I__2324 (
            .O(N__9864),
            .I(N__9860));
    InMux I__2323 (
            .O(N__9863),
            .I(N__9857));
    Odrv4 I__2322 (
            .O(N__9860),
            .I(DS_ENm));
    LocalMux I__2321 (
            .O(N__9857),
            .I(DS_ENm));
    InMux I__2320 (
            .O(N__9852),
            .I(N__9843));
    InMux I__2319 (
            .O(N__9851),
            .I(N__9843));
    InMux I__2318 (
            .O(N__9850),
            .I(N__9838));
    InMux I__2317 (
            .O(N__9849),
            .I(N__9838));
    CascadeMux I__2316 (
            .O(N__9848),
            .I(N__9835));
    LocalMux I__2315 (
            .O(N__9843),
            .I(N__9827));
    LocalMux I__2314 (
            .O(N__9838),
            .I(N__9824));
    InMux I__2313 (
            .O(N__9835),
            .I(N__9821));
    InMux I__2312 (
            .O(N__9834),
            .I(N__9818));
    InMux I__2311 (
            .O(N__9833),
            .I(N__9813));
    InMux I__2310 (
            .O(N__9832),
            .I(N__9813));
    InMux I__2309 (
            .O(N__9831),
            .I(N__9810));
    InMux I__2308 (
            .O(N__9830),
            .I(N__9807));
    Span4Mux_v I__2307 (
            .O(N__9827),
            .I(N__9804));
    Span4Mux_v I__2306 (
            .O(N__9824),
            .I(N__9801));
    LocalMux I__2305 (
            .O(N__9821),
            .I(N__9794));
    LocalMux I__2304 (
            .O(N__9818),
            .I(N__9794));
    LocalMux I__2303 (
            .O(N__9813),
            .I(N__9794));
    LocalMux I__2302 (
            .O(N__9810),
            .I(N__9789));
    LocalMux I__2301 (
            .O(N__9807),
            .I(N__9789));
    Span4Mux_v I__2300 (
            .O(N__9804),
            .I(N__9786));
    Span4Mux_v I__2299 (
            .O(N__9801),
            .I(N__9781));
    Span4Mux_v I__2298 (
            .O(N__9794),
            .I(N__9781));
    Span12Mux_s10_v I__2297 (
            .O(N__9789),
            .I(N__9778));
    Span4Mux_h I__2296 (
            .O(N__9786),
            .I(N__9775));
    Sp12to4 I__2295 (
            .O(N__9781),
            .I(N__9772));
    Span12Mux_h I__2294 (
            .O(N__9778),
            .I(N__9769));
    Sp12to4 I__2293 (
            .O(N__9775),
            .I(N__9764));
    Span12Mux_h I__2292 (
            .O(N__9772),
            .I(N__9764));
    Odrv12 I__2291 (
            .O(N__9769),
            .I(A_c_0));
    Odrv12 I__2290 (
            .O(N__9764),
            .I(A_c_0));
    CascadeMux I__2289 (
            .O(N__9759),
            .I(N__9755));
    InMux I__2288 (
            .O(N__9758),
            .I(N__9750));
    InMux I__2287 (
            .O(N__9755),
            .I(N__9750));
    LocalMux I__2286 (
            .O(N__9750),
            .I(N__9744));
    InMux I__2285 (
            .O(N__9749),
            .I(N__9740));
    InMux I__2284 (
            .O(N__9748),
            .I(N__9737));
    InMux I__2283 (
            .O(N__9747),
            .I(N__9734));
    Span4Mux_v I__2282 (
            .O(N__9744),
            .I(N__9729));
    InMux I__2281 (
            .O(N__9743),
            .I(N__9726));
    LocalMux I__2280 (
            .O(N__9740),
            .I(N__9723));
    LocalMux I__2279 (
            .O(N__9737),
            .I(N__9718));
    LocalMux I__2278 (
            .O(N__9734),
            .I(N__9718));
    InMux I__2277 (
            .O(N__9733),
            .I(N__9713));
    InMux I__2276 (
            .O(N__9732),
            .I(N__9713));
    Span4Mux_v I__2275 (
            .O(N__9729),
            .I(N__9707));
    LocalMux I__2274 (
            .O(N__9726),
            .I(N__9707));
    Span4Mux_v I__2273 (
            .O(N__9723),
            .I(N__9700));
    Span4Mux_h I__2272 (
            .O(N__9718),
            .I(N__9700));
    LocalMux I__2271 (
            .O(N__9713),
            .I(N__9700));
    InMux I__2270 (
            .O(N__9712),
            .I(N__9697));
    Span4Mux_v I__2269 (
            .O(N__9707),
            .I(N__9694));
    Span4Mux_h I__2268 (
            .O(N__9700),
            .I(N__9691));
    LocalMux I__2267 (
            .O(N__9697),
            .I(N__9688));
    Span4Mux_v I__2266 (
            .O(N__9694),
            .I(N__9685));
    Span4Mux_v I__2265 (
            .O(N__9691),
            .I(N__9682));
    Span12Mux_v I__2264 (
            .O(N__9688),
            .I(N__9679));
    Span4Mux_h I__2263 (
            .O(N__9685),
            .I(N__9676));
    Span4Mux_h I__2262 (
            .O(N__9682),
            .I(N__9673));
    Span12Mux_h I__2261 (
            .O(N__9679),
            .I(N__9670));
    Sp12to4 I__2260 (
            .O(N__9676),
            .I(N__9665));
    Sp12to4 I__2259 (
            .O(N__9673),
            .I(N__9665));
    Odrv12 I__2258 (
            .O(N__9670),
            .I(SIZ_c_0));
    Odrv12 I__2257 (
            .O(N__9665),
            .I(SIZ_c_0));
    IoInMux I__2256 (
            .O(N__9660),
            .I(N__9657));
    LocalMux I__2255 (
            .O(N__9657),
            .I(N__9654));
    Span4Mux_s2_v I__2254 (
            .O(N__9654),
            .I(N__9651));
    Span4Mux_h I__2253 (
            .O(N__9651),
            .I(N__9648));
    Span4Mux_v I__2252 (
            .O(N__9648),
            .I(N__9645));
    Odrv4 I__2251 (
            .O(N__9645),
            .I(N_87));
    InMux I__2250 (
            .O(N__9642),
            .I(N__9639));
    LocalMux I__2249 (
            .O(N__9639),
            .I(N__9636));
    Odrv4 I__2248 (
            .O(N__9636),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__2247 (
            .O(N__9633),
            .I(N__9630));
    LocalMux I__2246 (
            .O(N__9630),
            .I(N__9627));
    Span4Mux_h I__2245 (
            .O(N__9627),
            .I(N__9624));
    Odrv4 I__2244 (
            .O(N__9624),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__2243 (
            .O(N__9621),
            .I(N__9618));
    LocalMux I__2242 (
            .O(N__9618),
            .I(N__9615));
    Span4Mux_h I__2241 (
            .O(N__9615),
            .I(N__9612));
    Odrv4 I__2240 (
            .O(N__9612),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__2239 (
            .O(N__9609),
            .I(N__9606));
    LocalMux I__2238 (
            .O(N__9606),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__2237 (
            .O(N__9603),
            .I(N__9600));
    LocalMux I__2236 (
            .O(N__9600),
            .I(N__9594));
    InMux I__2235 (
            .O(N__9599),
            .I(N__9591));
    InMux I__2234 (
            .O(N__9598),
            .I(N__9588));
    InMux I__2233 (
            .O(N__9597),
            .I(N__9585));
    Span4Mux_v I__2232 (
            .O(N__9594),
            .I(N__9582));
    LocalMux I__2231 (
            .O(N__9591),
            .I(N__9577));
    LocalMux I__2230 (
            .O(N__9588),
            .I(N__9577));
    LocalMux I__2229 (
            .O(N__9585),
            .I(N__9574));
    Sp12to4 I__2228 (
            .O(N__9582),
            .I(N__9571));
    Span4Mux_v I__2227 (
            .O(N__9577),
            .I(N__9566));
    Span4Mux_h I__2226 (
            .O(N__9574),
            .I(N__9566));
    Span12Mux_h I__2225 (
            .O(N__9571),
            .I(N__9563));
    Sp12to4 I__2224 (
            .O(N__9566),
            .I(N__9560));
    Span12Mux_v I__2223 (
            .O(N__9563),
            .I(N__9557));
    Span12Mux_v I__2222 (
            .O(N__9560),
            .I(N__9554));
    Odrv12 I__2221 (
            .O(N__9557),
            .I(DRA_c_2));
    Odrv12 I__2220 (
            .O(N__9554),
            .I(DRA_c_2));
    InMux I__2219 (
            .O(N__9549),
            .I(N__9546));
    LocalMux I__2218 (
            .O(N__9546),
            .I(N__9543));
    Odrv12 I__2217 (
            .O(N__9543),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    IoInMux I__2216 (
            .O(N__9540),
            .I(N__9537));
    LocalMux I__2215 (
            .O(N__9537),
            .I(N__9534));
    Span4Mux_s2_v I__2214 (
            .O(N__9534),
            .I(N__9531));
    Span4Mux_v I__2213 (
            .O(N__9531),
            .I(N__9528));
    Span4Mux_v I__2212 (
            .O(N__9528),
            .I(N__9525));
    Span4Mux_h I__2211 (
            .O(N__9525),
            .I(N__9522));
    Odrv4 I__2210 (
            .O(N__9522),
            .I(CASn_c));
    CascadeMux I__2209 (
            .O(N__9519),
            .I(N__9508));
    CascadeMux I__2208 (
            .O(N__9518),
            .I(N__9505));
    CascadeMux I__2207 (
            .O(N__9517),
            .I(N__9498));
    CascadeMux I__2206 (
            .O(N__9516),
            .I(N__9495));
    CascadeMux I__2205 (
            .O(N__9515),
            .I(N__9491));
    CascadeMux I__2204 (
            .O(N__9514),
            .I(N__9488));
    CascadeMux I__2203 (
            .O(N__9513),
            .I(N__9484));
    CascadeMux I__2202 (
            .O(N__9512),
            .I(N__9480));
    CascadeMux I__2201 (
            .O(N__9511),
            .I(N__9477));
    InMux I__2200 (
            .O(N__9508),
            .I(N__9467));
    InMux I__2199 (
            .O(N__9505),
            .I(N__9467));
    InMux I__2198 (
            .O(N__9504),
            .I(N__9458));
    InMux I__2197 (
            .O(N__9503),
            .I(N__9458));
    InMux I__2196 (
            .O(N__9502),
            .I(N__9458));
    InMux I__2195 (
            .O(N__9501),
            .I(N__9458));
    InMux I__2194 (
            .O(N__9498),
            .I(N__9455));
    InMux I__2193 (
            .O(N__9495),
            .I(N__9450));
    InMux I__2192 (
            .O(N__9494),
            .I(N__9450));
    InMux I__2191 (
            .O(N__9491),
            .I(N__9447));
    InMux I__2190 (
            .O(N__9488),
            .I(N__9444));
    InMux I__2189 (
            .O(N__9487),
            .I(N__9439));
    InMux I__2188 (
            .O(N__9484),
            .I(N__9439));
    InMux I__2187 (
            .O(N__9483),
            .I(N__9434));
    InMux I__2186 (
            .O(N__9480),
            .I(N__9434));
    InMux I__2185 (
            .O(N__9477),
            .I(N__9431));
    InMux I__2184 (
            .O(N__9476),
            .I(N__9428));
    InMux I__2183 (
            .O(N__9475),
            .I(N__9425));
    InMux I__2182 (
            .O(N__9474),
            .I(N__9417));
    InMux I__2181 (
            .O(N__9473),
            .I(N__9417));
    InMux I__2180 (
            .O(N__9472),
            .I(N__9414));
    LocalMux I__2179 (
            .O(N__9467),
            .I(N__9405));
    LocalMux I__2178 (
            .O(N__9458),
            .I(N__9405));
    LocalMux I__2177 (
            .O(N__9455),
            .I(N__9405));
    LocalMux I__2176 (
            .O(N__9450),
            .I(N__9405));
    LocalMux I__2175 (
            .O(N__9447),
            .I(N__9400));
    LocalMux I__2174 (
            .O(N__9444),
            .I(N__9400));
    LocalMux I__2173 (
            .O(N__9439),
            .I(N__9397));
    LocalMux I__2172 (
            .O(N__9434),
            .I(N__9393));
    LocalMux I__2171 (
            .O(N__9431),
            .I(N__9388));
    LocalMux I__2170 (
            .O(N__9428),
            .I(N__9388));
    LocalMux I__2169 (
            .O(N__9425),
            .I(N__9385));
    InMux I__2168 (
            .O(N__9424),
            .I(N__9382));
    InMux I__2167 (
            .O(N__9423),
            .I(N__9379));
    InMux I__2166 (
            .O(N__9422),
            .I(N__9375));
    LocalMux I__2165 (
            .O(N__9417),
            .I(N__9372));
    LocalMux I__2164 (
            .O(N__9414),
            .I(N__9369));
    Span4Mux_v I__2163 (
            .O(N__9405),
            .I(N__9366));
    Span4Mux_h I__2162 (
            .O(N__9400),
            .I(N__9361));
    Span4Mux_v I__2161 (
            .O(N__9397),
            .I(N__9361));
    InMux I__2160 (
            .O(N__9396),
            .I(N__9358));
    Span4Mux_v I__2159 (
            .O(N__9393),
            .I(N__9351));
    Span4Mux_h I__2158 (
            .O(N__9388),
            .I(N__9351));
    Span4Mux_h I__2157 (
            .O(N__9385),
            .I(N__9351));
    LocalMux I__2156 (
            .O(N__9382),
            .I(N__9348));
    LocalMux I__2155 (
            .O(N__9379),
            .I(N__9345));
    InMux I__2154 (
            .O(N__9378),
            .I(N__9342));
    LocalMux I__2153 (
            .O(N__9375),
            .I(N__9329));
    Span12Mux_v I__2152 (
            .O(N__9372),
            .I(N__9329));
    Span12Mux_h I__2151 (
            .O(N__9369),
            .I(N__9329));
    Sp12to4 I__2150 (
            .O(N__9366),
            .I(N__9329));
    Sp12to4 I__2149 (
            .O(N__9361),
            .I(N__9329));
    LocalMux I__2148 (
            .O(N__9358),
            .I(N__9329));
    Span4Mux_h I__2147 (
            .O(N__9351),
            .I(N__9326));
    Span4Mux_v I__2146 (
            .O(N__9348),
            .I(N__9323));
    Odrv4 I__2145 (
            .O(N__9345),
            .I(CPU_CYCLEm));
    LocalMux I__2144 (
            .O(N__9342),
            .I(CPU_CYCLEm));
    Odrv12 I__2143 (
            .O(N__9329),
            .I(CPU_CYCLEm));
    Odrv4 I__2142 (
            .O(N__9326),
            .I(CPU_CYCLEm));
    Odrv4 I__2141 (
            .O(N__9323),
            .I(CPU_CYCLEm));
    InMux I__2140 (
            .O(N__9312),
            .I(N__9309));
    LocalMux I__2139 (
            .O(N__9309),
            .I(N__9306));
    Span12Mux_h I__2138 (
            .O(N__9306),
            .I(N__9303));
    Odrv12 I__2137 (
            .O(N__9303),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ));
    CascadeMux I__2136 (
            .O(N__9300),
            .I(N__9296));
    InMux I__2135 (
            .O(N__9299),
            .I(N__9291));
    InMux I__2134 (
            .O(N__9296),
            .I(N__9288));
    CascadeMux I__2133 (
            .O(N__9295),
            .I(N__9285));
    InMux I__2132 (
            .O(N__9294),
            .I(N__9275));
    LocalMux I__2131 (
            .O(N__9291),
            .I(N__9267));
    LocalMux I__2130 (
            .O(N__9288),
            .I(N__9267));
    InMux I__2129 (
            .O(N__9285),
            .I(N__9264));
    InMux I__2128 (
            .O(N__9284),
            .I(N__9259));
    InMux I__2127 (
            .O(N__9283),
            .I(N__9259));
    InMux I__2126 (
            .O(N__9282),
            .I(N__9252));
    InMux I__2125 (
            .O(N__9281),
            .I(N__9252));
    InMux I__2124 (
            .O(N__9280),
            .I(N__9252));
    InMux I__2123 (
            .O(N__9279),
            .I(N__9245));
    InMux I__2122 (
            .O(N__9278),
            .I(N__9245));
    LocalMux I__2121 (
            .O(N__9275),
            .I(N__9241));
    InMux I__2120 (
            .O(N__9274),
            .I(N__9236));
    InMux I__2119 (
            .O(N__9273),
            .I(N__9236));
    CascadeMux I__2118 (
            .O(N__9272),
            .I(N__9232));
    Span4Mux_v I__2117 (
            .O(N__9267),
            .I(N__9223));
    LocalMux I__2116 (
            .O(N__9264),
            .I(N__9223));
    LocalMux I__2115 (
            .O(N__9259),
            .I(N__9223));
    LocalMux I__2114 (
            .O(N__9252),
            .I(N__9223));
    InMux I__2113 (
            .O(N__9251),
            .I(N__9218));
    InMux I__2112 (
            .O(N__9250),
            .I(N__9218));
    LocalMux I__2111 (
            .O(N__9245),
            .I(N__9215));
    CascadeMux I__2110 (
            .O(N__9244),
            .I(N__9210));
    Span4Mux_v I__2109 (
            .O(N__9241),
            .I(N__9206));
    LocalMux I__2108 (
            .O(N__9236),
            .I(N__9203));
    InMux I__2107 (
            .O(N__9235),
            .I(N__9200));
    InMux I__2106 (
            .O(N__9232),
            .I(N__9194));
    Span4Mux_h I__2105 (
            .O(N__9223),
            .I(N__9187));
    LocalMux I__2104 (
            .O(N__9218),
            .I(N__9187));
    Span4Mux_v I__2103 (
            .O(N__9215),
            .I(N__9187));
    InMux I__2102 (
            .O(N__9214),
            .I(N__9180));
    InMux I__2101 (
            .O(N__9213),
            .I(N__9180));
    InMux I__2100 (
            .O(N__9210),
            .I(N__9180));
    InMux I__2099 (
            .O(N__9209),
            .I(N__9177));
    Span4Mux_h I__2098 (
            .O(N__9206),
            .I(N__9170));
    Span4Mux_v I__2097 (
            .O(N__9203),
            .I(N__9170));
    LocalMux I__2096 (
            .O(N__9200),
            .I(N__9170));
    InMux I__2095 (
            .O(N__9199),
            .I(N__9167));
    InMux I__2094 (
            .O(N__9198),
            .I(N__9162));
    InMux I__2093 (
            .O(N__9197),
            .I(N__9162));
    LocalMux I__2092 (
            .O(N__9194),
            .I(N__9155));
    Sp12to4 I__2091 (
            .O(N__9187),
            .I(N__9155));
    LocalMux I__2090 (
            .O(N__9180),
            .I(N__9155));
    LocalMux I__2089 (
            .O(N__9177),
            .I(N__9150));
    Span4Mux_h I__2088 (
            .O(N__9170),
            .I(N__9150));
    LocalMux I__2087 (
            .O(N__9167),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2086 (
            .O(N__9162),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv12 I__2085 (
            .O(N__9155),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2084 (
            .O(N__9150),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    InMux I__2083 (
            .O(N__9141),
            .I(N__9138));
    LocalMux I__2082 (
            .O(N__9138),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ));
    IoInMux I__2081 (
            .O(N__9135),
            .I(N__9132));
    LocalMux I__2080 (
            .O(N__9132),
            .I(N__9129));
    Sp12to4 I__2079 (
            .O(N__9129),
            .I(N__9126));
    Span12Mux_h I__2078 (
            .O(N__9126),
            .I(N__9123));
    Odrv12 I__2077 (
            .O(N__9123),
            .I(CMA_c_4));
    InMux I__2076 (
            .O(N__9120),
            .I(N__9117));
    LocalMux I__2075 (
            .O(N__9117),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ));
    IoInMux I__2074 (
            .O(N__9114),
            .I(N__9111));
    LocalMux I__2073 (
            .O(N__9111),
            .I(N__9108));
    Span4Mux_s2_h I__2072 (
            .O(N__9108),
            .I(N__9105));
    Sp12to4 I__2071 (
            .O(N__9105),
            .I(N__9102));
    Span12Mux_v I__2070 (
            .O(N__9102),
            .I(N__9099));
    Odrv12 I__2069 (
            .O(N__9099),
            .I(CMA_c_7));
    InMux I__2068 (
            .O(N__9096),
            .I(N__9091));
    InMux I__2067 (
            .O(N__9095),
            .I(N__9086));
    InMux I__2066 (
            .O(N__9094),
            .I(N__9086));
    LocalMux I__2065 (
            .O(N__9091),
            .I(N__9079));
    LocalMux I__2064 (
            .O(N__9086),
            .I(N__9079));
    InMux I__2063 (
            .O(N__9085),
            .I(N__9076));
    InMux I__2062 (
            .O(N__9084),
            .I(N__9070));
    Span4Mux_h I__2061 (
            .O(N__9079),
            .I(N__9065));
    LocalMux I__2060 (
            .O(N__9076),
            .I(N__9065));
    InMux I__2059 (
            .O(N__9075),
            .I(N__9062));
    InMux I__2058 (
            .O(N__9074),
            .I(N__9059));
    InMux I__2057 (
            .O(N__9073),
            .I(N__9056));
    LocalMux I__2056 (
            .O(N__9070),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__2055 (
            .O(N__9065),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__2054 (
            .O(N__9062),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__2053 (
            .O(N__9059),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__2052 (
            .O(N__9056),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    CascadeMux I__2051 (
            .O(N__9045),
            .I(N__9038));
    CascadeMux I__2050 (
            .O(N__9044),
            .I(N__9035));
    CascadeMux I__2049 (
            .O(N__9043),
            .I(N__9032));
    CascadeMux I__2048 (
            .O(N__9042),
            .I(N__9028));
    InMux I__2047 (
            .O(N__9041),
            .I(N__9021));
    InMux I__2046 (
            .O(N__9038),
            .I(N__9021));
    InMux I__2045 (
            .O(N__9035),
            .I(N__9021));
    InMux I__2044 (
            .O(N__9032),
            .I(N__9018));
    CascadeMux I__2043 (
            .O(N__9031),
            .I(N__9015));
    InMux I__2042 (
            .O(N__9028),
            .I(N__9012));
    LocalMux I__2041 (
            .O(N__9021),
            .I(N__9007));
    LocalMux I__2040 (
            .O(N__9018),
            .I(N__9007));
    InMux I__2039 (
            .O(N__9015),
            .I(N__9004));
    LocalMux I__2038 (
            .O(N__9012),
            .I(N__8999));
    Span4Mux_v I__2037 (
            .O(N__9007),
            .I(N__8999));
    LocalMux I__2036 (
            .O(N__9004),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNIHMEAZ0Z_1 ));
    Odrv4 I__2035 (
            .O(N__8999),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNIHMEAZ0Z_1 ));
    InMux I__2034 (
            .O(N__8994),
            .I(N__8991));
    LocalMux I__2033 (
            .O(N__8991),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ));
    IoInMux I__2032 (
            .O(N__8988),
            .I(N__8985));
    LocalMux I__2031 (
            .O(N__8985),
            .I(N__8982));
    Span4Mux_s3_h I__2030 (
            .O(N__8982),
            .I(N__8979));
    Sp12to4 I__2029 (
            .O(N__8979),
            .I(N__8976));
    Span12Mux_v I__2028 (
            .O(N__8976),
            .I(N__8973));
    Odrv12 I__2027 (
            .O(N__8973),
            .I(CMA_c_6));
    InMux I__2026 (
            .O(N__8970),
            .I(N__8967));
    LocalMux I__2025 (
            .O(N__8967),
            .I(N__8940));
    ClkMux I__2024 (
            .O(N__8966),
            .I(N__8844));
    ClkMux I__2023 (
            .O(N__8965),
            .I(N__8844));
    ClkMux I__2022 (
            .O(N__8964),
            .I(N__8844));
    ClkMux I__2021 (
            .O(N__8963),
            .I(N__8844));
    ClkMux I__2020 (
            .O(N__8962),
            .I(N__8844));
    ClkMux I__2019 (
            .O(N__8961),
            .I(N__8844));
    ClkMux I__2018 (
            .O(N__8960),
            .I(N__8844));
    ClkMux I__2017 (
            .O(N__8959),
            .I(N__8844));
    ClkMux I__2016 (
            .O(N__8958),
            .I(N__8844));
    ClkMux I__2015 (
            .O(N__8957),
            .I(N__8844));
    ClkMux I__2014 (
            .O(N__8956),
            .I(N__8844));
    ClkMux I__2013 (
            .O(N__8955),
            .I(N__8844));
    ClkMux I__2012 (
            .O(N__8954),
            .I(N__8844));
    ClkMux I__2011 (
            .O(N__8953),
            .I(N__8844));
    ClkMux I__2010 (
            .O(N__8952),
            .I(N__8844));
    ClkMux I__2009 (
            .O(N__8951),
            .I(N__8844));
    ClkMux I__2008 (
            .O(N__8950),
            .I(N__8844));
    ClkMux I__2007 (
            .O(N__8949),
            .I(N__8844));
    ClkMux I__2006 (
            .O(N__8948),
            .I(N__8844));
    ClkMux I__2005 (
            .O(N__8947),
            .I(N__8844));
    ClkMux I__2004 (
            .O(N__8946),
            .I(N__8844));
    ClkMux I__2003 (
            .O(N__8945),
            .I(N__8844));
    ClkMux I__2002 (
            .O(N__8944),
            .I(N__8844));
    ClkMux I__2001 (
            .O(N__8943),
            .I(N__8844));
    Glb2LocalMux I__2000 (
            .O(N__8940),
            .I(N__8844));
    ClkMux I__1999 (
            .O(N__8939),
            .I(N__8844));
    ClkMux I__1998 (
            .O(N__8938),
            .I(N__8844));
    ClkMux I__1997 (
            .O(N__8937),
            .I(N__8844));
    ClkMux I__1996 (
            .O(N__8936),
            .I(N__8844));
    ClkMux I__1995 (
            .O(N__8935),
            .I(N__8844));
    ClkMux I__1994 (
            .O(N__8934),
            .I(N__8844));
    ClkMux I__1993 (
            .O(N__8933),
            .I(N__8844));
    ClkMux I__1992 (
            .O(N__8932),
            .I(N__8844));
    ClkMux I__1991 (
            .O(N__8931),
            .I(N__8844));
    ClkMux I__1990 (
            .O(N__8930),
            .I(N__8844));
    ClkMux I__1989 (
            .O(N__8929),
            .I(N__8844));
    ClkMux I__1988 (
            .O(N__8928),
            .I(N__8844));
    ClkMux I__1987 (
            .O(N__8927),
            .I(N__8844));
    ClkMux I__1986 (
            .O(N__8926),
            .I(N__8844));
    ClkMux I__1985 (
            .O(N__8925),
            .I(N__8844));
    GlobalMux I__1984 (
            .O(N__8844),
            .I(CLK80_PLL));
    CEMux I__1983 (
            .O(N__8841),
            .I(N__8838));
    LocalMux I__1982 (
            .O(N__8838),
            .I(N__8832));
    CEMux I__1981 (
            .O(N__8837),
            .I(N__8828));
    CEMux I__1980 (
            .O(N__8836),
            .I(N__8825));
    CEMux I__1979 (
            .O(N__8835),
            .I(N__8822));
    Span4Mux_h I__1978 (
            .O(N__8832),
            .I(N__8819));
    CEMux I__1977 (
            .O(N__8831),
            .I(N__8816));
    LocalMux I__1976 (
            .O(N__8828),
            .I(N__8812));
    LocalMux I__1975 (
            .O(N__8825),
            .I(N__8807));
    LocalMux I__1974 (
            .O(N__8822),
            .I(N__8807));
    Span4Mux_h I__1973 (
            .O(N__8819),
            .I(N__8802));
    LocalMux I__1972 (
            .O(N__8816),
            .I(N__8802));
    CEMux I__1971 (
            .O(N__8815),
            .I(N__8799));
    Span4Mux_v I__1970 (
            .O(N__8812),
            .I(N__8796));
    Sp12to4 I__1969 (
            .O(N__8807),
            .I(N__8793));
    Sp12to4 I__1968 (
            .O(N__8802),
            .I(N__8788));
    LocalMux I__1967 (
            .O(N__8799),
            .I(N__8788));
    Odrv4 I__1966 (
            .O(N__8796),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv12 I__1965 (
            .O(N__8793),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv12 I__1964 (
            .O(N__8788),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    InMux I__1963 (
            .O(N__8781),
            .I(N__8778));
    LocalMux I__1962 (
            .O(N__8778),
            .I(N__8775));
    Span12Mux_h I__1961 (
            .O(N__8775),
            .I(N__8772));
    Odrv12 I__1960 (
            .O(N__8772),
            .I(RAS0n_c));
    InMux I__1959 (
            .O(N__8769),
            .I(N__8766));
    LocalMux I__1958 (
            .O(N__8766),
            .I(N__8763));
    Odrv4 I__1957 (
            .O(N__8763),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    InMux I__1956 (
            .O(N__8760),
            .I(N__8754));
    InMux I__1955 (
            .O(N__8759),
            .I(N__8754));
    LocalMux I__1954 (
            .O(N__8754),
            .I(N__8751));
    Span4Mux_v I__1953 (
            .O(N__8751),
            .I(N__8748));
    Span4Mux_h I__1952 (
            .O(N__8748),
            .I(N__8745));
    Odrv4 I__1951 (
            .O(N__8745),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    CascadeMux I__1950 (
            .O(N__8742),
            .I(N__8739));
    InMux I__1949 (
            .O(N__8739),
            .I(N__8736));
    LocalMux I__1948 (
            .O(N__8736),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__1947 (
            .O(N__8733),
            .I(N__8730));
    LocalMux I__1946 (
            .O(N__8730),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ));
    IoInMux I__1945 (
            .O(N__8727),
            .I(N__8724));
    LocalMux I__1944 (
            .O(N__8724),
            .I(N__8721));
    Span4Mux_s0_v I__1943 (
            .O(N__8721),
            .I(N__8718));
    Span4Mux_v I__1942 (
            .O(N__8718),
            .I(N__8715));
    Span4Mux_v I__1941 (
            .O(N__8715),
            .I(N__8712));
    Span4Mux_v I__1940 (
            .O(N__8712),
            .I(N__8709));
    Odrv4 I__1939 (
            .O(N__8709),
            .I(CMA_c_0));
    InMux I__1938 (
            .O(N__8706),
            .I(N__8703));
    LocalMux I__1937 (
            .O(N__8703),
            .I(N__8700));
    Span4Mux_h I__1936 (
            .O(N__8700),
            .I(N__8697));
    Odrv4 I__1935 (
            .O(N__8697),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ));
    InMux I__1934 (
            .O(N__8694),
            .I(N__8691));
    LocalMux I__1933 (
            .O(N__8691),
            .I(N__8688));
    Span4Mux_v I__1932 (
            .O(N__8688),
            .I(N__8685));
    Sp12to4 I__1931 (
            .O(N__8685),
            .I(N__8682));
    Span12Mux_h I__1930 (
            .O(N__8682),
            .I(N__8679));
    Odrv12 I__1929 (
            .O(N__8679),
            .I(A_c_13));
    InMux I__1928 (
            .O(N__8676),
            .I(N__8673));
    LocalMux I__1927 (
            .O(N__8673),
            .I(N__8670));
    Span4Mux_h I__1926 (
            .O(N__8670),
            .I(N__8667));
    Span4Mux_v I__1925 (
            .O(N__8667),
            .I(N__8664));
    Sp12to4 I__1924 (
            .O(N__8664),
            .I(N__8661));
    Span12Mux_h I__1923 (
            .O(N__8661),
            .I(N__8658));
    Odrv12 I__1922 (
            .O(N__8658),
            .I(A_c_6));
    CascadeMux I__1921 (
            .O(N__8655),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ));
    InMux I__1920 (
            .O(N__8652),
            .I(N__8649));
    LocalMux I__1919 (
            .O(N__8649),
            .I(N__8645));
    InMux I__1918 (
            .O(N__8648),
            .I(N__8642));
    Span4Mux_h I__1917 (
            .O(N__8645),
            .I(N__8639));
    LocalMux I__1916 (
            .O(N__8642),
            .I(N__8636));
    Span4Mux_h I__1915 (
            .O(N__8639),
            .I(N__8631));
    Span4Mux_v I__1914 (
            .O(N__8636),
            .I(N__8631));
    Odrv4 I__1913 (
            .O(N__8631),
            .I(DBRn_c_i));
    InMux I__1912 (
            .O(N__8628),
            .I(N__8625));
    LocalMux I__1911 (
            .O(N__8625),
            .I(N__8621));
    InMux I__1910 (
            .O(N__8624),
            .I(N__8618));
    Span12Mux_h I__1909 (
            .O(N__8621),
            .I(N__8615));
    LocalMux I__1908 (
            .O(N__8618),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    Odrv12 I__1907 (
            .O(N__8615),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    IoInMux I__1906 (
            .O(N__8610),
            .I(N__8607));
    LocalMux I__1905 (
            .O(N__8607),
            .I(N__8604));
    Span12Mux_s7_v I__1904 (
            .O(N__8604),
            .I(N__8601));
    Odrv12 I__1903 (
            .O(N__8601),
            .I(UMBEn_c));
    CascadeMux I__1902 (
            .O(N__8598),
            .I(N__8595));
    InMux I__1901 (
            .O(N__8595),
            .I(N__8587));
    InMux I__1900 (
            .O(N__8594),
            .I(N__8587));
    InMux I__1899 (
            .O(N__8593),
            .I(N__8582));
    InMux I__1898 (
            .O(N__8592),
            .I(N__8582));
    LocalMux I__1897 (
            .O(N__8587),
            .I(N__8578));
    LocalMux I__1896 (
            .O(N__8582),
            .I(N__8575));
    CascadeMux I__1895 (
            .O(N__8581),
            .I(N__8571));
    Span4Mux_v I__1894 (
            .O(N__8578),
            .I(N__8567));
    Span4Mux_v I__1893 (
            .O(N__8575),
            .I(N__8564));
    InMux I__1892 (
            .O(N__8574),
            .I(N__8561));
    InMux I__1891 (
            .O(N__8571),
            .I(N__8556));
    InMux I__1890 (
            .O(N__8570),
            .I(N__8556));
    Span4Mux_v I__1889 (
            .O(N__8567),
            .I(N__8553));
    Span4Mux_v I__1888 (
            .O(N__8564),
            .I(N__8550));
    LocalMux I__1887 (
            .O(N__8561),
            .I(N__8545));
    LocalMux I__1886 (
            .O(N__8556),
            .I(N__8545));
    Span4Mux_v I__1885 (
            .O(N__8553),
            .I(N__8541));
    Span4Mux_v I__1884 (
            .O(N__8550),
            .I(N__8536));
    Span4Mux_v I__1883 (
            .O(N__8545),
            .I(N__8536));
    InMux I__1882 (
            .O(N__8544),
            .I(N__8533));
    Sp12to4 I__1881 (
            .O(N__8541),
            .I(N__8526));
    Sp12to4 I__1880 (
            .O(N__8536),
            .I(N__8526));
    LocalMux I__1879 (
            .O(N__8533),
            .I(N__8526));
    Span12Mux_h I__1878 (
            .O(N__8526),
            .I(N__8523));
    Odrv12 I__1877 (
            .O(N__8523),
            .I(A_c_1));
    CascadeMux I__1876 (
            .O(N__8520),
            .I(N__8517));
    InMux I__1875 (
            .O(N__8517),
            .I(N__8512));
    InMux I__1874 (
            .O(N__8516),
            .I(N__8509));
    InMux I__1873 (
            .O(N__8515),
            .I(N__8506));
    LocalMux I__1872 (
            .O(N__8512),
            .I(N__8502));
    LocalMux I__1871 (
            .O(N__8509),
            .I(N__8499));
    LocalMux I__1870 (
            .O(N__8506),
            .I(N__8496));
    CascadeMux I__1869 (
            .O(N__8505),
            .I(N__8492));
    Span4Mux_v I__1868 (
            .O(N__8502),
            .I(N__8489));
    Span4Mux_v I__1867 (
            .O(N__8499),
            .I(N__8484));
    Span4Mux_h I__1866 (
            .O(N__8496),
            .I(N__8484));
    InMux I__1865 (
            .O(N__8495),
            .I(N__8479));
    InMux I__1864 (
            .O(N__8492),
            .I(N__8479));
    Span4Mux_v I__1863 (
            .O(N__8489),
            .I(N__8476));
    Span4Mux_v I__1862 (
            .O(N__8484),
            .I(N__8473));
    LocalMux I__1861 (
            .O(N__8479),
            .I(N__8470));
    Sp12to4 I__1860 (
            .O(N__8476),
            .I(N__8463));
    Sp12to4 I__1859 (
            .O(N__8473),
            .I(N__8463));
    Span12Mux_v I__1858 (
            .O(N__8470),
            .I(N__8463));
    Span12Mux_h I__1857 (
            .O(N__8463),
            .I(N__8460));
    Odrv12 I__1856 (
            .O(N__8460),
            .I(SIZ_c_1));
    IoInMux I__1855 (
            .O(N__8457),
            .I(N__8454));
    LocalMux I__1854 (
            .O(N__8454),
            .I(N__8451));
    Span4Mux_s3_v I__1853 (
            .O(N__8451),
            .I(N__8448));
    Odrv4 I__1852 (
            .O(N__8448),
            .I(N_276_i));
    InMux I__1851 (
            .O(N__8445),
            .I(N__8441));
    InMux I__1850 (
            .O(N__8444),
            .I(N__8438));
    LocalMux I__1849 (
            .O(N__8441),
            .I(N__8434));
    LocalMux I__1848 (
            .O(N__8438),
            .I(N__8430));
    InMux I__1847 (
            .O(N__8437),
            .I(N__8427));
    Span4Mux_h I__1846 (
            .O(N__8434),
            .I(N__8424));
    CascadeMux I__1845 (
            .O(N__8433),
            .I(N__8419));
    Span4Mux_h I__1844 (
            .O(N__8430),
            .I(N__8414));
    LocalMux I__1843 (
            .O(N__8427),
            .I(N__8414));
    Span4Mux_v I__1842 (
            .O(N__8424),
            .I(N__8411));
    InMux I__1841 (
            .O(N__8423),
            .I(N__8408));
    InMux I__1840 (
            .O(N__8422),
            .I(N__8405));
    InMux I__1839 (
            .O(N__8419),
            .I(N__8401));
    Span4Mux_h I__1838 (
            .O(N__8414),
            .I(N__8398));
    Sp12to4 I__1837 (
            .O(N__8411),
            .I(N__8391));
    LocalMux I__1836 (
            .O(N__8408),
            .I(N__8391));
    LocalMux I__1835 (
            .O(N__8405),
            .I(N__8391));
    InMux I__1834 (
            .O(N__8404),
            .I(N__8388));
    LocalMux I__1833 (
            .O(N__8401),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1832 (
            .O(N__8398),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv12 I__1831 (
            .O(N__8391),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1830 (
            .O(N__8388),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    IoInMux I__1829 (
            .O(N__8379),
            .I(N__8376));
    LocalMux I__1828 (
            .O(N__8376),
            .I(N__8373));
    Span4Mux_s2_v I__1827 (
            .O(N__8373),
            .I(N__8370));
    Span4Mux_v I__1826 (
            .O(N__8370),
            .I(N__8367));
    Span4Mux_h I__1825 (
            .O(N__8367),
            .I(N__8364));
    Odrv4 I__1824 (
            .O(N__8364),
            .I(RASn_c));
    CascadeMux I__1823 (
            .O(N__8361),
            .I(N__8358));
    InMux I__1822 (
            .O(N__8358),
            .I(N__8354));
    InMux I__1821 (
            .O(N__8357),
            .I(N__8351));
    LocalMux I__1820 (
            .O(N__8354),
            .I(N__8348));
    LocalMux I__1819 (
            .O(N__8351),
            .I(N__8341));
    Sp12to4 I__1818 (
            .O(N__8348),
            .I(N__8341));
    InMux I__1817 (
            .O(N__8347),
            .I(N__8338));
    InMux I__1816 (
            .O(N__8346),
            .I(N__8334));
    Span12Mux_v I__1815 (
            .O(N__8341),
            .I(N__8329));
    LocalMux I__1814 (
            .O(N__8338),
            .I(N__8329));
    InMux I__1813 (
            .O(N__8337),
            .I(N__8326));
    LocalMux I__1812 (
            .O(N__8334),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv12 I__1811 (
            .O(N__8329),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__1810 (
            .O(N__8326),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__1809 (
            .O(N__8319),
            .I(N__8316));
    LocalMux I__1808 (
            .O(N__8316),
            .I(N__8313));
    Span4Mux_s2_v I__1807 (
            .O(N__8313),
            .I(N__8310));
    Span4Mux_v I__1806 (
            .O(N__8310),
            .I(N__8307));
    Span4Mux_h I__1805 (
            .O(N__8307),
            .I(N__8304));
    Odrv4 I__1804 (
            .O(N__8304),
            .I(CRCSn_c));
    InMux I__1803 (
            .O(N__8301),
            .I(N__8298));
    LocalMux I__1802 (
            .O(N__8298),
            .I(\U712_BYTE_ENABLE.N_339 ));
    InMux I__1801 (
            .O(N__8295),
            .I(N__8289));
    InMux I__1800 (
            .O(N__8294),
            .I(N__8289));
    LocalMux I__1799 (
            .O(N__8289),
            .I(N__8286));
    Span4Mux_v I__1798 (
            .O(N__8286),
            .I(N__8281));
    InMux I__1797 (
            .O(N__8285),
            .I(N__8276));
    InMux I__1796 (
            .O(N__8284),
            .I(N__8276));
    Span4Mux_v I__1795 (
            .O(N__8281),
            .I(N__8273));
    LocalMux I__1794 (
            .O(N__8276),
            .I(N__8270));
    Odrv4 I__1793 (
            .O(N__8273),
            .I(\U712_BYTE_ENABLE.N_206_i ));
    Odrv12 I__1792 (
            .O(N__8270),
            .I(\U712_BYTE_ENABLE.N_206_i ));
    InMux I__1791 (
            .O(N__8265),
            .I(N__8262));
    LocalMux I__1790 (
            .O(N__8262),
            .I(N__8259));
    Span4Mux_h I__1789 (
            .O(N__8259),
            .I(N__8256));
    Odrv4 I__1788 (
            .O(N__8256),
            .I(\U712_BYTE_ENABLE.N_316 ));
    IoInMux I__1787 (
            .O(N__8253),
            .I(N__8250));
    LocalMux I__1786 (
            .O(N__8250),
            .I(N__8247));
    Span4Mux_s3_v I__1785 (
            .O(N__8247),
            .I(N__8244));
    Odrv4 I__1784 (
            .O(N__8244),
            .I(N_277_i));
    IoInMux I__1783 (
            .O(N__8241),
            .I(N__8238));
    LocalMux I__1782 (
            .O(N__8238),
            .I(N__8235));
    Span4Mux_s2_v I__1781 (
            .O(N__8235),
            .I(N__8232));
    Span4Mux_v I__1780 (
            .O(N__8232),
            .I(N__8229));
    Odrv4 I__1779 (
            .O(N__8229),
            .I(LLBE_i_o2_i));
    IoInMux I__1778 (
            .O(N__8226),
            .I(N__8223));
    LocalMux I__1777 (
            .O(N__8223),
            .I(N__8220));
    IoSpan4Mux I__1776 (
            .O(N__8220),
            .I(N__8217));
    Sp12to4 I__1775 (
            .O(N__8217),
            .I(N__8214));
    Span12Mux_s7_v I__1774 (
            .O(N__8214),
            .I(N__8211));
    Span12Mux_h I__1773 (
            .O(N__8211),
            .I(N__8208));
    Odrv12 I__1772 (
            .O(N__8208),
            .I(WEn_c));
    InMux I__1771 (
            .O(N__8205),
            .I(N__8202));
    LocalMux I__1770 (
            .O(N__8202),
            .I(N__8199));
    Sp12to4 I__1769 (
            .O(N__8199),
            .I(N__8196));
    Span12Mux_v I__1768 (
            .O(N__8196),
            .I(N__8193));
    Span12Mux_h I__1767 (
            .O(N__8193),
            .I(N__8190));
    Odrv12 I__1766 (
            .O(N__8190),
            .I(A_c_17));
    IoInMux I__1765 (
            .O(N__8187),
            .I(N__8184));
    LocalMux I__1764 (
            .O(N__8184),
            .I(N__8181));
    IoSpan4Mux I__1763 (
            .O(N__8181),
            .I(N__8178));
    IoSpan4Mux I__1762 (
            .O(N__8178),
            .I(N__8175));
    Span4Mux_s2_h I__1761 (
            .O(N__8175),
            .I(N__8172));
    Sp12to4 I__1760 (
            .O(N__8172),
            .I(N__8169));
    Odrv12 I__1759 (
            .O(N__8169),
            .I(CMA_c_8));
    InMux I__1758 (
            .O(N__8166),
            .I(N__8163));
    LocalMux I__1757 (
            .O(N__8163),
            .I(N__8160));
    Sp12to4 I__1756 (
            .O(N__8160),
            .I(N__8157));
    Span12Mux_v I__1755 (
            .O(N__8157),
            .I(N__8154));
    Span12Mux_h I__1754 (
            .O(N__8154),
            .I(N__8151));
    Odrv12 I__1753 (
            .O(N__8151),
            .I(A_c_19));
    InMux I__1752 (
            .O(N__8148),
            .I(N__8142));
    InMux I__1751 (
            .O(N__8147),
            .I(N__8142));
    LocalMux I__1750 (
            .O(N__8142),
            .I(N__8139));
    Span4Mux_h I__1749 (
            .O(N__8139),
            .I(N__8134));
    InMux I__1748 (
            .O(N__8138),
            .I(N__8129));
    InMux I__1747 (
            .O(N__8137),
            .I(N__8129));
    Odrv4 I__1746 (
            .O(N__8134),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    LocalMux I__1745 (
            .O(N__8129),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    IoInMux I__1744 (
            .O(N__8124),
            .I(N__8121));
    LocalMux I__1743 (
            .O(N__8121),
            .I(N__8118));
    IoSpan4Mux I__1742 (
            .O(N__8118),
            .I(N__8115));
    Span4Mux_s3_h I__1741 (
            .O(N__8115),
            .I(N__8112));
    Sp12to4 I__1740 (
            .O(N__8112),
            .I(N__8109));
    Span12Mux_h I__1739 (
            .O(N__8109),
            .I(N__8106));
    Odrv12 I__1738 (
            .O(N__8106),
            .I(CMA_c_9));
    InMux I__1737 (
            .O(N__8103),
            .I(N__8098));
    InMux I__1736 (
            .O(N__8102),
            .I(N__8094));
    CascadeMux I__1735 (
            .O(N__8101),
            .I(N__8090));
    LocalMux I__1734 (
            .O(N__8098),
            .I(N__8086));
    InMux I__1733 (
            .O(N__8097),
            .I(N__8083));
    LocalMux I__1732 (
            .O(N__8094),
            .I(N__8080));
    InMux I__1731 (
            .O(N__8093),
            .I(N__8077));
    InMux I__1730 (
            .O(N__8090),
            .I(N__8073));
    InMux I__1729 (
            .O(N__8089),
            .I(N__8070));
    Span4Mux_h I__1728 (
            .O(N__8086),
            .I(N__8065));
    LocalMux I__1727 (
            .O(N__8083),
            .I(N__8065));
    Span4Mux_v I__1726 (
            .O(N__8080),
            .I(N__8062));
    LocalMux I__1725 (
            .O(N__8077),
            .I(N__8059));
    CascadeMux I__1724 (
            .O(N__8076),
            .I(N__8056));
    LocalMux I__1723 (
            .O(N__8073),
            .I(N__8053));
    LocalMux I__1722 (
            .O(N__8070),
            .I(N__8048));
    Span4Mux_v I__1721 (
            .O(N__8065),
            .I(N__8048));
    Span4Mux_h I__1720 (
            .O(N__8062),
            .I(N__8043));
    Span4Mux_h I__1719 (
            .O(N__8059),
            .I(N__8043));
    InMux I__1718 (
            .O(N__8056),
            .I(N__8040));
    Odrv4 I__1717 (
            .O(N__8053),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1716 (
            .O(N__8048),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1715 (
            .O(N__8043),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1714 (
            .O(N__8040),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    IoInMux I__1713 (
            .O(N__8031),
            .I(N__8028));
    LocalMux I__1712 (
            .O(N__8028),
            .I(N__8025));
    Span4Mux_s3_v I__1711 (
            .O(N__8025),
            .I(N__8022));
    Span4Mux_v I__1710 (
            .O(N__8022),
            .I(N__8019));
    Span4Mux_v I__1709 (
            .O(N__8019),
            .I(N__8016));
    Span4Mux_h I__1708 (
            .O(N__8016),
            .I(N__8013));
    Odrv4 I__1707 (
            .O(N__8013),
            .I(CMA_c_10));
    InMux I__1706 (
            .O(N__8010),
            .I(N__8007));
    LocalMux I__1705 (
            .O(N__8007),
            .I(\U712_BYTE_ENABLE.N_320 ));
    CascadeMux I__1704 (
            .O(N__8004),
            .I(\U712_BYTE_ENABLE.N_318_cascade_ ));
    IoInMux I__1703 (
            .O(N__8001),
            .I(N__7998));
    LocalMux I__1702 (
            .O(N__7998),
            .I(N__7995));
    IoSpan4Mux I__1701 (
            .O(N__7995),
            .I(N__7992));
    Span4Mux_s3_h I__1700 (
            .O(N__7992),
            .I(N__7989));
    Sp12to4 I__1699 (
            .O(N__7989),
            .I(N__7986));
    Span12Mux_s10_v I__1698 (
            .O(N__7986),
            .I(N__7983));
    Span12Mux_h I__1697 (
            .O(N__7983),
            .I(N__7980));
    Odrv12 I__1696 (
            .O(N__7980),
            .I(N_105_i));
    IoInMux I__1695 (
            .O(N__7977),
            .I(N__7974));
    LocalMux I__1694 (
            .O(N__7974),
            .I(N__7971));
    Span4Mux_s3_v I__1693 (
            .O(N__7971),
            .I(N__7968));
    Span4Mux_v I__1692 (
            .O(N__7968),
            .I(N__7965));
    Span4Mux_v I__1691 (
            .O(N__7965),
            .I(N__7962));
    Odrv4 I__1690 (
            .O(N__7962),
            .I(CMA_c_2));
    InMux I__1689 (
            .O(N__7959),
            .I(N__7956));
    LocalMux I__1688 (
            .O(N__7956),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i ));
    InMux I__1687 (
            .O(N__7953),
            .I(N__7950));
    LocalMux I__1686 (
            .O(N__7950),
            .I(N__7947));
    Span12Mux_v I__1685 (
            .O(N__7947),
            .I(N__7944));
    Span12Mux_h I__1684 (
            .O(N__7944),
            .I(N__7941));
    Odrv12 I__1683 (
            .O(N__7941),
            .I(A_c_4));
    InMux I__1682 (
            .O(N__7938),
            .I(N__7935));
    LocalMux I__1681 (
            .O(N__7935),
            .I(N__7932));
    Span4Mux_v I__1680 (
            .O(N__7932),
            .I(N__7929));
    Sp12to4 I__1679 (
            .O(N__7929),
            .I(N__7926));
    Span12Mux_h I__1678 (
            .O(N__7926),
            .I(N__7923));
    Odrv12 I__1677 (
            .O(N__7923),
            .I(A_c_11));
    CascadeMux I__1676 (
            .O(N__7920),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ));
    InMux I__1675 (
            .O(N__7917),
            .I(N__7914));
    LocalMux I__1674 (
            .O(N__7914),
            .I(N__7911));
    Odrv4 I__1673 (
            .O(N__7911),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ));
    InMux I__1672 (
            .O(N__7908),
            .I(N__7905));
    LocalMux I__1671 (
            .O(N__7905),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ));
    InMux I__1670 (
            .O(N__7902),
            .I(N__7894));
    InMux I__1669 (
            .O(N__7901),
            .I(N__7889));
    InMux I__1668 (
            .O(N__7900),
            .I(N__7889));
    InMux I__1667 (
            .O(N__7899),
            .I(N__7886));
    InMux I__1666 (
            .O(N__7898),
            .I(N__7883));
    InMux I__1665 (
            .O(N__7897),
            .I(N__7880));
    LocalMux I__1664 (
            .O(N__7894),
            .I(N__7877));
    LocalMux I__1663 (
            .O(N__7889),
            .I(N__7871));
    LocalMux I__1662 (
            .O(N__7886),
            .I(N__7871));
    LocalMux I__1661 (
            .O(N__7883),
            .I(N__7868));
    LocalMux I__1660 (
            .O(N__7880),
            .I(N__7865));
    Span4Mux_v I__1659 (
            .O(N__7877),
            .I(N__7861));
    InMux I__1658 (
            .O(N__7876),
            .I(N__7858));
    Span4Mux_v I__1657 (
            .O(N__7871),
            .I(N__7853));
    Span4Mux_v I__1656 (
            .O(N__7868),
            .I(N__7853));
    Span4Mux_h I__1655 (
            .O(N__7865),
            .I(N__7850));
    InMux I__1654 (
            .O(N__7864),
            .I(N__7847));
    Odrv4 I__1653 (
            .O(N__7861),
            .I(DMA_CYCLEm));
    LocalMux I__1652 (
            .O(N__7858),
            .I(DMA_CYCLEm));
    Odrv4 I__1651 (
            .O(N__7853),
            .I(DMA_CYCLEm));
    Odrv4 I__1650 (
            .O(N__7850),
            .I(DMA_CYCLEm));
    LocalMux I__1649 (
            .O(N__7847),
            .I(DMA_CYCLEm));
    InMux I__1648 (
            .O(N__7836),
            .I(N__7833));
    LocalMux I__1647 (
            .O(N__7833),
            .I(N__7828));
    CascadeMux I__1646 (
            .O(N__7832),
            .I(N__7824));
    CascadeMux I__1645 (
            .O(N__7831),
            .I(N__7820));
    Span4Mux_v I__1644 (
            .O(N__7828),
            .I(N__7817));
    InMux I__1643 (
            .O(N__7827),
            .I(N__7814));
    InMux I__1642 (
            .O(N__7824),
            .I(N__7811));
    InMux I__1641 (
            .O(N__7823),
            .I(N__7808));
    InMux I__1640 (
            .O(N__7820),
            .I(N__7805));
    Span4Mux_v I__1639 (
            .O(N__7817),
            .I(N__7800));
    LocalMux I__1638 (
            .O(N__7814),
            .I(N__7800));
    LocalMux I__1637 (
            .O(N__7811),
            .I(N__7797));
    LocalMux I__1636 (
            .O(N__7808),
            .I(N__7794));
    LocalMux I__1635 (
            .O(N__7805),
            .I(N__7790));
    Span4Mux_v I__1634 (
            .O(N__7800),
            .I(N__7787));
    Span4Mux_v I__1633 (
            .O(N__7797),
            .I(N__7782));
    Span4Mux_v I__1632 (
            .O(N__7794),
            .I(N__7782));
    InMux I__1631 (
            .O(N__7793),
            .I(N__7779));
    Span12Mux_v I__1630 (
            .O(N__7790),
            .I(N__7776));
    Span4Mux_v I__1629 (
            .O(N__7787),
            .I(N__7773));
    Sp12to4 I__1628 (
            .O(N__7782),
            .I(N__7770));
    LocalMux I__1627 (
            .O(N__7779),
            .I(N__7767));
    Span12Mux_h I__1626 (
            .O(N__7776),
            .I(N__7764));
    Sp12to4 I__1625 (
            .O(N__7773),
            .I(N__7761));
    Span12Mux_h I__1624 (
            .O(N__7770),
            .I(N__7758));
    Span12Mux_v I__1623 (
            .O(N__7767),
            .I(N__7755));
    Span12Mux_v I__1622 (
            .O(N__7764),
            .I(N__7752));
    Span12Mux_h I__1621 (
            .O(N__7761),
            .I(N__7749));
    Span12Mux_v I__1620 (
            .O(N__7758),
            .I(N__7744));
    Span12Mux_h I__1619 (
            .O(N__7755),
            .I(N__7744));
    Odrv12 I__1618 (
            .O(N__7752),
            .I(CASUn_c));
    Odrv12 I__1617 (
            .O(N__7749),
            .I(CASUn_c));
    Odrv12 I__1616 (
            .O(N__7744),
            .I(CASUn_c));
    IoInMux I__1615 (
            .O(N__7737),
            .I(N__7734));
    LocalMux I__1614 (
            .O(N__7734),
            .I(N__7730));
    InMux I__1613 (
            .O(N__7733),
            .I(N__7727));
    IoSpan4Mux I__1612 (
            .O(N__7730),
            .I(N__7721));
    LocalMux I__1611 (
            .O(N__7727),
            .I(N__7718));
    InMux I__1610 (
            .O(N__7726),
            .I(N__7713));
    InMux I__1609 (
            .O(N__7725),
            .I(N__7713));
    InMux I__1608 (
            .O(N__7724),
            .I(N__7710));
    Span4Mux_s2_v I__1607 (
            .O(N__7721),
            .I(N__7707));
    Span4Mux_v I__1606 (
            .O(N__7718),
            .I(N__7700));
    LocalMux I__1605 (
            .O(N__7713),
            .I(N__7700));
    LocalMux I__1604 (
            .O(N__7710),
            .I(N__7700));
    Span4Mux_v I__1603 (
            .O(N__7707),
            .I(N__7697));
    Span4Mux_h I__1602 (
            .O(N__7700),
            .I(N__7694));
    Span4Mux_v I__1601 (
            .O(N__7697),
            .I(N__7688));
    Span4Mux_v I__1600 (
            .O(N__7694),
            .I(N__7688));
    InMux I__1599 (
            .O(N__7693),
            .I(N__7685));
    Odrv4 I__1598 (
            .O(N__7688),
            .I(DBENn_c));
    LocalMux I__1597 (
            .O(N__7685),
            .I(DBENn_c));
    IoInMux I__1596 (
            .O(N__7680),
            .I(N__7677));
    LocalMux I__1595 (
            .O(N__7677),
            .I(N__7674));
    IoSpan4Mux I__1594 (
            .O(N__7674),
            .I(N__7671));
    Span4Mux_s3_h I__1593 (
            .O(N__7671),
            .I(N__7668));
    Sp12to4 I__1592 (
            .O(N__7668),
            .I(N__7665));
    Span12Mux_h I__1591 (
            .O(N__7665),
            .I(N__7662));
    Odrv12 I__1590 (
            .O(N__7662),
            .I(N_57_i));
    CascadeMux I__1589 (
            .O(N__7659),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_ ));
    InMux I__1588 (
            .O(N__7656),
            .I(N__7653));
    LocalMux I__1587 (
            .O(N__7653),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ));
    InMux I__1586 (
            .O(N__7650),
            .I(N__7647));
    LocalMux I__1585 (
            .O(N__7647),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ));
    InMux I__1584 (
            .O(N__7644),
            .I(N__7641));
    LocalMux I__1583 (
            .O(N__7641),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ));
    InMux I__1582 (
            .O(N__7638),
            .I(N__7635));
    LocalMux I__1581 (
            .O(N__7635),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ));
    IoInMux I__1580 (
            .O(N__7632),
            .I(N__7629));
    LocalMux I__1579 (
            .O(N__7629),
            .I(N__7626));
    Span4Mux_s3_h I__1578 (
            .O(N__7626),
            .I(N__7623));
    Span4Mux_v I__1577 (
            .O(N__7623),
            .I(N__7620));
    Sp12to4 I__1576 (
            .O(N__7620),
            .I(N__7617));
    Span12Mux_h I__1575 (
            .O(N__7617),
            .I(N__7614));
    Odrv12 I__1574 (
            .O(N__7614),
            .I(CMA_c_5));
    InMux I__1573 (
            .O(N__7611),
            .I(N__7608));
    LocalMux I__1572 (
            .O(N__7608),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ));
    InMux I__1571 (
            .O(N__7605),
            .I(N__7602));
    LocalMux I__1570 (
            .O(N__7602),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ));
    InMux I__1569 (
            .O(N__7599),
            .I(N__7596));
    LocalMux I__1568 (
            .O(N__7596),
            .I(N__7593));
    Span4Mux_v I__1567 (
            .O(N__7593),
            .I(N__7590));
    Sp12to4 I__1566 (
            .O(N__7590),
            .I(N__7587));
    Span12Mux_h I__1565 (
            .O(N__7587),
            .I(N__7584));
    Span12Mux_v I__1564 (
            .O(N__7584),
            .I(N__7581));
    Odrv12 I__1563 (
            .O(N__7581),
            .I(A_c_2));
    InMux I__1562 (
            .O(N__7578),
            .I(N__7575));
    LocalMux I__1561 (
            .O(N__7575),
            .I(N__7572));
    Span4Mux_v I__1560 (
            .O(N__7572),
            .I(N__7569));
    Sp12to4 I__1559 (
            .O(N__7569),
            .I(N__7566));
    Span12Mux_h I__1558 (
            .O(N__7566),
            .I(N__7563));
    Odrv12 I__1557 (
            .O(N__7563),
            .I(A_c_9));
    InMux I__1556 (
            .O(N__7560),
            .I(N__7557));
    LocalMux I__1555 (
            .O(N__7557),
            .I(N__7554));
    Span4Mux_v I__1554 (
            .O(N__7554),
            .I(N__7547));
    InMux I__1553 (
            .O(N__7553),
            .I(N__7544));
    CascadeMux I__1552 (
            .O(N__7552),
            .I(N__7541));
    InMux I__1551 (
            .O(N__7551),
            .I(N__7536));
    InMux I__1550 (
            .O(N__7550),
            .I(N__7536));
    Span4Mux_v I__1549 (
            .O(N__7547),
            .I(N__7531));
    LocalMux I__1548 (
            .O(N__7544),
            .I(N__7531));
    InMux I__1547 (
            .O(N__7541),
            .I(N__7528));
    LocalMux I__1546 (
            .O(N__7536),
            .I(N__7524));
    Span4Mux_v I__1545 (
            .O(N__7531),
            .I(N__7521));
    LocalMux I__1544 (
            .O(N__7528),
            .I(N__7518));
    InMux I__1543 (
            .O(N__7527),
            .I(N__7515));
    Span4Mux_v I__1542 (
            .O(N__7524),
            .I(N__7512));
    Span4Mux_h I__1541 (
            .O(N__7521),
            .I(N__7507));
    Span4Mux_v I__1540 (
            .O(N__7518),
            .I(N__7507));
    LocalMux I__1539 (
            .O(N__7515),
            .I(N__7504));
    Sp12to4 I__1538 (
            .O(N__7512),
            .I(N__7501));
    Span4Mux_v I__1537 (
            .O(N__7507),
            .I(N__7498));
    Span12Mux_v I__1536 (
            .O(N__7504),
            .I(N__7495));
    Span12Mux_h I__1535 (
            .O(N__7501),
            .I(N__7492));
    Sp12to4 I__1534 (
            .O(N__7498),
            .I(N__7489));
    Span12Mux_h I__1533 (
            .O(N__7495),
            .I(N__7486));
    Span12Mux_v I__1532 (
            .O(N__7492),
            .I(N__7481));
    Span12Mux_h I__1531 (
            .O(N__7489),
            .I(N__7481));
    Odrv12 I__1530 (
            .O(N__7486),
            .I(CASLn_c));
    Odrv12 I__1529 (
            .O(N__7481),
            .I(CASLn_c));
    InMux I__1528 (
            .O(N__7476),
            .I(N__7473));
    LocalMux I__1527 (
            .O(N__7473),
            .I(\U712_BYTE_ENABLE.N_342 ));
    CascadeMux I__1526 (
            .O(N__7470),
            .I(\U712_BYTE_ENABLE.N_341_cascade_ ));
    IoInMux I__1525 (
            .O(N__7467),
            .I(N__7464));
    LocalMux I__1524 (
            .O(N__7464),
            .I(N__7461));
    Span4Mux_s2_v I__1523 (
            .O(N__7461),
            .I(N__7458));
    Span4Mux_h I__1522 (
            .O(N__7458),
            .I(N__7455));
    Sp12to4 I__1521 (
            .O(N__7455),
            .I(N__7452));
    Span12Mux_v I__1520 (
            .O(N__7452),
            .I(N__7449));
    Odrv12 I__1519 (
            .O(N__7449),
            .I(N_55_i));
    InMux I__1518 (
            .O(N__7446),
            .I(N__7443));
    LocalMux I__1517 (
            .O(N__7443),
            .I(N__7440));
    Odrv12 I__1516 (
            .O(N__7440),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ));
    InMux I__1515 (
            .O(N__7437),
            .I(N__7434));
    LocalMux I__1514 (
            .O(N__7434),
            .I(N__7431));
    Span4Mux_v I__1513 (
            .O(N__7431),
            .I(N__7428));
    Sp12to4 I__1512 (
            .O(N__7428),
            .I(N__7425));
    Span12Mux_h I__1511 (
            .O(N__7425),
            .I(N__7422));
    Span12Mux_v I__1510 (
            .O(N__7422),
            .I(N__7419));
    Odrv12 I__1509 (
            .O(N__7419),
            .I(A_c_3));
    InMux I__1508 (
            .O(N__7416),
            .I(N__7413));
    LocalMux I__1507 (
            .O(N__7413),
            .I(N__7410));
    Span4Mux_v I__1506 (
            .O(N__7410),
            .I(N__7407));
    Sp12to4 I__1505 (
            .O(N__7407),
            .I(N__7404));
    Span12Mux_h I__1504 (
            .O(N__7404),
            .I(N__7401));
    Odrv12 I__1503 (
            .O(N__7401),
            .I(A_c_10));
    IoInMux I__1502 (
            .O(N__7398),
            .I(N__7395));
    LocalMux I__1501 (
            .O(N__7395),
            .I(N__7392));
    IoSpan4Mux I__1500 (
            .O(N__7392),
            .I(N__7389));
    IoSpan4Mux I__1499 (
            .O(N__7389),
            .I(N__7386));
    Span4Mux_s3_h I__1498 (
            .O(N__7386),
            .I(N__7383));
    Sp12to4 I__1497 (
            .O(N__7383),
            .I(N__7380));
    Odrv12 I__1496 (
            .O(N__7380),
            .I(N_180_i));
    InMux I__1495 (
            .O(N__7377),
            .I(N__7367));
    InMux I__1494 (
            .O(N__7376),
            .I(N__7367));
    InMux I__1493 (
            .O(N__7375),
            .I(N__7362));
    InMux I__1492 (
            .O(N__7374),
            .I(N__7362));
    InMux I__1491 (
            .O(N__7373),
            .I(N__7357));
    InMux I__1490 (
            .O(N__7372),
            .I(N__7357));
    LocalMux I__1489 (
            .O(N__7367),
            .I(N__7346));
    LocalMux I__1488 (
            .O(N__7362),
            .I(N__7346));
    LocalMux I__1487 (
            .O(N__7357),
            .I(N__7346));
    InMux I__1486 (
            .O(N__7356),
            .I(N__7343));
    InMux I__1485 (
            .O(N__7355),
            .I(N__7339));
    InMux I__1484 (
            .O(N__7354),
            .I(N__7336));
    InMux I__1483 (
            .O(N__7353),
            .I(N__7333));
    Span4Mux_h I__1482 (
            .O(N__7346),
            .I(N__7324));
    LocalMux I__1481 (
            .O(N__7343),
            .I(N__7324));
    InMux I__1480 (
            .O(N__7342),
            .I(N__7321));
    LocalMux I__1479 (
            .O(N__7339),
            .I(N__7318));
    LocalMux I__1478 (
            .O(N__7336),
            .I(N__7315));
    LocalMux I__1477 (
            .O(N__7333),
            .I(N__7312));
    InMux I__1476 (
            .O(N__7332),
            .I(N__7307));
    InMux I__1475 (
            .O(N__7331),
            .I(N__7307));
    InMux I__1474 (
            .O(N__7330),
            .I(N__7304));
    InMux I__1473 (
            .O(N__7329),
            .I(N__7301));
    Span4Mux_h I__1472 (
            .O(N__7324),
            .I(N__7296));
    LocalMux I__1471 (
            .O(N__7321),
            .I(N__7296));
    Span4Mux_v I__1470 (
            .O(N__7318),
            .I(N__7293));
    Span4Mux_v I__1469 (
            .O(N__7315),
            .I(N__7282));
    Span4Mux_v I__1468 (
            .O(N__7312),
            .I(N__7282));
    LocalMux I__1467 (
            .O(N__7307),
            .I(N__7282));
    LocalMux I__1466 (
            .O(N__7304),
            .I(N__7282));
    LocalMux I__1465 (
            .O(N__7301),
            .I(N__7282));
    Span4Mux_v I__1464 (
            .O(N__7296),
            .I(N__7278));
    Span4Mux_v I__1463 (
            .O(N__7293),
            .I(N__7273));
    Span4Mux_v I__1462 (
            .O(N__7282),
            .I(N__7273));
    InMux I__1461 (
            .O(N__7281),
            .I(N__7270));
    Sp12to4 I__1460 (
            .O(N__7278),
            .I(N__7263));
    Sp12to4 I__1459 (
            .O(N__7273),
            .I(N__7263));
    LocalMux I__1458 (
            .O(N__7270),
            .I(N__7263));
    Span12Mux_h I__1457 (
            .O(N__7263),
            .I(N__7260));
    Odrv12 I__1456 (
            .O(N__7260),
            .I(RESETn_c));
    IoInMux I__1455 (
            .O(N__7257),
            .I(N__7254));
    LocalMux I__1454 (
            .O(N__7254),
            .I(N__7251));
    Sp12to4 I__1453 (
            .O(N__7251),
            .I(N__7248));
    Odrv12 I__1452 (
            .O(N__7248),
            .I(RESETn_c_i));
    InMux I__1451 (
            .O(N__7245),
            .I(N__7242));
    LocalMux I__1450 (
            .O(N__7242),
            .I(N__7239));
    Odrv4 I__1449 (
            .O(N__7239),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    IoInMux I__1448 (
            .O(N__7236),
            .I(N__7233));
    LocalMux I__1447 (
            .O(N__7233),
            .I(N__7230));
    IoSpan4Mux I__1446 (
            .O(N__7230),
            .I(N__7227));
    Span4Mux_s1_h I__1445 (
            .O(N__7227),
            .I(N__7224));
    Sp12to4 I__1444 (
            .O(N__7224),
            .I(N__7221));
    Span12Mux_h I__1443 (
            .O(N__7221),
            .I(N__7218));
    Odrv12 I__1442 (
            .O(N__7218),
            .I(CMA_c_3));
    CascadeMux I__1441 (
            .O(N__7215),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1_cascade_ ));
    IoInMux I__1440 (
            .O(N__7212),
            .I(N__7209));
    LocalMux I__1439 (
            .O(N__7209),
            .I(N__7206));
    Span4Mux_s2_v I__1438 (
            .O(N__7206),
            .I(N__7203));
    Sp12to4 I__1437 (
            .O(N__7203),
            .I(N__7200));
    Span12Mux_h I__1436 (
            .O(N__7200),
            .I(N__7197));
    Odrv12 I__1435 (
            .O(N__7197),
            .I(CMA_c_1));
    SRMux I__1434 (
            .O(N__7194),
            .I(N__7191));
    LocalMux I__1433 (
            .O(N__7191),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    InMux I__1432 (
            .O(N__7188),
            .I(N__7184));
    InMux I__1431 (
            .O(N__7187),
            .I(N__7181));
    LocalMux I__1430 (
            .O(N__7184),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__1429 (
            .O(N__7181),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__1428 (
            .O(N__7176),
            .I(N__7172));
    InMux I__1427 (
            .O(N__7175),
            .I(N__7169));
    LocalMux I__1426 (
            .O(N__7172),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__1425 (
            .O(N__7169),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__1424 (
            .O(N__7164),
            .I(N__7160));
    InMux I__1423 (
            .O(N__7163),
            .I(N__7157));
    LocalMux I__1422 (
            .O(N__7160),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    LocalMux I__1421 (
            .O(N__7157),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    InMux I__1420 (
            .O(N__7152),
            .I(N__7149));
    LocalMux I__1419 (
            .O(N__7149),
            .I(N__7146));
    Odrv4 I__1418 (
            .O(N__7146),
            .I(\U712_CHIP_RAM.REFRESH5lt7 ));
    IoInMux I__1417 (
            .O(N__7143),
            .I(N__7140));
    LocalMux I__1416 (
            .O(N__7140),
            .I(N__7137));
    Span4Mux_s2_v I__1415 (
            .O(N__7137),
            .I(N__7133));
    InMux I__1414 (
            .O(N__7136),
            .I(N__7130));
    Span4Mux_v I__1413 (
            .O(N__7133),
            .I(N__7127));
    LocalMux I__1412 (
            .O(N__7130),
            .I(N__7124));
    Span4Mux_v I__1411 (
            .O(N__7127),
            .I(N__7121));
    Span4Mux_v I__1410 (
            .O(N__7124),
            .I(N__7118));
    Odrv4 I__1409 (
            .O(N__7121),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1408 (
            .O(N__7118),
            .I(CONSTANT_ONE_NET));
    InMux I__1407 (
            .O(N__7113),
            .I(N__7110));
    LocalMux I__1406 (
            .O(N__7110),
            .I(N__7107));
    Span12Mux_v I__1405 (
            .O(N__7107),
            .I(N__7104));
    Span12Mux_h I__1404 (
            .O(N__7104),
            .I(N__7101));
    Odrv12 I__1403 (
            .O(N__7101),
            .I(A_c_7));
    CascadeMux I__1402 (
            .O(N__7098),
            .I(\U712_CHIP_RAM.N_231_cascade_ ));
    CascadeMux I__1401 (
            .O(N__7095),
            .I(N__7092));
    InMux I__1400 (
            .O(N__7092),
            .I(N__7086));
    InMux I__1399 (
            .O(N__7091),
            .I(N__7086));
    LocalMux I__1398 (
            .O(N__7086),
            .I(N__7083));
    Span4Mux_v I__1397 (
            .O(N__7083),
            .I(N__7080));
    Span4Mux_v I__1396 (
            .O(N__7080),
            .I(N__7077));
    Sp12to4 I__1395 (
            .O(N__7077),
            .I(N__7074));
    Span12Mux_h I__1394 (
            .O(N__7074),
            .I(N__7071));
    Odrv12 I__1393 (
            .O(N__7071),
            .I(A_c_14));
    CascadeMux I__1392 (
            .O(N__7068),
            .I(N__7064));
    InMux I__1391 (
            .O(N__7067),
            .I(N__7059));
    InMux I__1390 (
            .O(N__7064),
            .I(N__7056));
    InMux I__1389 (
            .O(N__7063),
            .I(N__7051));
    InMux I__1388 (
            .O(N__7062),
            .I(N__7051));
    LocalMux I__1387 (
            .O(N__7059),
            .I(N__7044));
    LocalMux I__1386 (
            .O(N__7056),
            .I(N__7044));
    LocalMux I__1385 (
            .O(N__7051),
            .I(N__7044));
    Span4Mux_v I__1384 (
            .O(N__7044),
            .I(N__7041));
    Span4Mux_v I__1383 (
            .O(N__7041),
            .I(N__7038));
    Span4Mux_v I__1382 (
            .O(N__7038),
            .I(N__7035));
    IoSpan4Mux I__1381 (
            .O(N__7035),
            .I(N__7032));
    Odrv4 I__1380 (
            .O(N__7032),
            .I(CLK40_PLL_i));
    IoInMux I__1379 (
            .O(N__7029),
            .I(N__7026));
    LocalMux I__1378 (
            .O(N__7026),
            .I(N__7022));
    IoInMux I__1377 (
            .O(N__7025),
            .I(N__7019));
    IoSpan4Mux I__1376 (
            .O(N__7022),
            .I(N__7013));
    LocalMux I__1375 (
            .O(N__7019),
            .I(N__7013));
    IoInMux I__1374 (
            .O(N__7018),
            .I(N__7010));
    IoSpan4Mux I__1373 (
            .O(N__7013),
            .I(N__7007));
    LocalMux I__1372 (
            .O(N__7010),
            .I(N__7004));
    IoSpan4Mux I__1371 (
            .O(N__7007),
            .I(N__7001));
    Span4Mux_s3_h I__1370 (
            .O(N__7004),
            .I(N__6998));
    Sp12to4 I__1369 (
            .O(N__7001),
            .I(N__6995));
    Span4Mux_h I__1368 (
            .O(N__6998),
            .I(N__6992));
    Span12Mux_s6_v I__1367 (
            .O(N__6995),
            .I(N__6989));
    Span4Mux_h I__1366 (
            .O(N__6992),
            .I(N__6986));
    Span12Mux_v I__1365 (
            .O(N__6989),
            .I(N__6983));
    Span4Mux_h I__1364 (
            .O(N__6986),
            .I(N__6980));
    Odrv12 I__1363 (
            .O(N__6983),
            .I(CLK40_PLL_i_i));
    Odrv4 I__1362 (
            .O(N__6980),
            .I(CLK40_PLL_i_i));
    InMux I__1361 (
            .O(N__6975),
            .I(N__6968));
    InMux I__1360 (
            .O(N__6974),
            .I(N__6968));
    InMux I__1359 (
            .O(N__6973),
            .I(N__6965));
    LocalMux I__1358 (
            .O(N__6968),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__1357 (
            .O(N__6965),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    InMux I__1356 (
            .O(N__6960),
            .I(N__6956));
    InMux I__1355 (
            .O(N__6959),
            .I(N__6953));
    LocalMux I__1354 (
            .O(N__6956),
            .I(N__6950));
    LocalMux I__1353 (
            .O(N__6953),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    Odrv4 I__1352 (
            .O(N__6950),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    InMux I__1351 (
            .O(N__6945),
            .I(N__6942));
    LocalMux I__1350 (
            .O(N__6942),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ));
    InMux I__1349 (
            .O(N__6939),
            .I(N__6936));
    LocalMux I__1348 (
            .O(N__6936),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ));
    InMux I__1347 (
            .O(N__6933),
            .I(bfn_11_10_0_));
    InMux I__1346 (
            .O(N__6930),
            .I(N__6927));
    LocalMux I__1345 (
            .O(N__6927),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    InMux I__1344 (
            .O(N__6924),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__1343 (
            .O(N__6921),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__1342 (
            .O(N__6918),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    InMux I__1341 (
            .O(N__6915),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__1340 (
            .O(N__6912),
            .I(N__6908));
    InMux I__1339 (
            .O(N__6911),
            .I(N__6905));
    LocalMux I__1338 (
            .O(N__6908),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__1337 (
            .O(N__6905),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__1336 (
            .O(N__6900),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__1335 (
            .O(N__6897),
            .I(N__6893));
    InMux I__1334 (
            .O(N__6896),
            .I(N__6890));
    LocalMux I__1333 (
            .O(N__6893),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__1332 (
            .O(N__6890),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__1331 (
            .O(N__6885),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__1330 (
            .O(N__6882),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    CascadeMux I__1329 (
            .O(N__6879),
            .I(N__6876));
    InMux I__1328 (
            .O(N__6876),
            .I(N__6872));
    InMux I__1327 (
            .O(N__6875),
            .I(N__6869));
    LocalMux I__1326 (
            .O(N__6872),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    LocalMux I__1325 (
            .O(N__6869),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    ClkMux I__1324 (
            .O(N__6864),
            .I(N__6846));
    ClkMux I__1323 (
            .O(N__6863),
            .I(N__6846));
    ClkMux I__1322 (
            .O(N__6862),
            .I(N__6846));
    ClkMux I__1321 (
            .O(N__6861),
            .I(N__6846));
    ClkMux I__1320 (
            .O(N__6860),
            .I(N__6846));
    ClkMux I__1319 (
            .O(N__6859),
            .I(N__6846));
    GlobalMux I__1318 (
            .O(N__6846),
            .I(N__6843));
    gio2CtrlBuf I__1317 (
            .O(N__6843),
            .I(C1_c_g));
    CascadeMux I__1316 (
            .O(N__6840),
            .I(N__6836));
    InMux I__1315 (
            .O(N__6839),
            .I(N__6833));
    InMux I__1314 (
            .O(N__6836),
            .I(N__6830));
    LocalMux I__1313 (
            .O(N__6833),
            .I(N__6827));
    LocalMux I__1312 (
            .O(N__6830),
            .I(\U712_CHIP_RAM.N_314 ));
    Odrv4 I__1311 (
            .O(N__6827),
            .I(\U712_CHIP_RAM.N_314 ));
    CascadeMux I__1310 (
            .O(N__6822),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_cascade_ ));
    InMux I__1309 (
            .O(N__6819),
            .I(N__6816));
    LocalMux I__1308 (
            .O(N__6816),
            .I(\U712_CHIP_RAM.N_37 ));
    InMux I__1307 (
            .O(N__6813),
            .I(N__6809));
    InMux I__1306 (
            .O(N__6812),
            .I(N__6806));
    LocalMux I__1305 (
            .O(N__6809),
            .I(N__6803));
    LocalMux I__1304 (
            .O(N__6806),
            .I(CPU_TACKm));
    Odrv4 I__1303 (
            .O(N__6803),
            .I(CPU_TACKm));
    InMux I__1302 (
            .O(N__6798),
            .I(N__6794));
    InMux I__1301 (
            .O(N__6797),
            .I(N__6787));
    LocalMux I__1300 (
            .O(N__6794),
            .I(N__6781));
    InMux I__1299 (
            .O(N__6793),
            .I(N__6778));
    InMux I__1298 (
            .O(N__6792),
            .I(N__6775));
    InMux I__1297 (
            .O(N__6791),
            .I(N__6770));
    InMux I__1296 (
            .O(N__6790),
            .I(N__6770));
    LocalMux I__1295 (
            .O(N__6787),
            .I(N__6765));
    InMux I__1294 (
            .O(N__6786),
            .I(N__6762));
    InMux I__1293 (
            .O(N__6785),
            .I(N__6759));
    InMux I__1292 (
            .O(N__6784),
            .I(N__6756));
    Span4Mux_v I__1291 (
            .O(N__6781),
            .I(N__6747));
    LocalMux I__1290 (
            .O(N__6778),
            .I(N__6747));
    LocalMux I__1289 (
            .O(N__6775),
            .I(N__6747));
    LocalMux I__1288 (
            .O(N__6770),
            .I(N__6743));
    InMux I__1287 (
            .O(N__6769),
            .I(N__6737));
    InMux I__1286 (
            .O(N__6768),
            .I(N__6734));
    Span4Mux_h I__1285 (
            .O(N__6765),
            .I(N__6729));
    LocalMux I__1284 (
            .O(N__6762),
            .I(N__6729));
    LocalMux I__1283 (
            .O(N__6759),
            .I(N__6724));
    LocalMux I__1282 (
            .O(N__6756),
            .I(N__6724));
    InMux I__1281 (
            .O(N__6755),
            .I(N__6721));
    InMux I__1280 (
            .O(N__6754),
            .I(N__6718));
    Span4Mux_h I__1279 (
            .O(N__6747),
            .I(N__6715));
    InMux I__1278 (
            .O(N__6746),
            .I(N__6712));
    Span4Mux_h I__1277 (
            .O(N__6743),
            .I(N__6709));
    InMux I__1276 (
            .O(N__6742),
            .I(N__6702));
    InMux I__1275 (
            .O(N__6741),
            .I(N__6702));
    InMux I__1274 (
            .O(N__6740),
            .I(N__6702));
    LocalMux I__1273 (
            .O(N__6737),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1272 (
            .O(N__6734),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1271 (
            .O(N__6729),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1270 (
            .O(N__6724),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1269 (
            .O(N__6721),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1268 (
            .O(N__6718),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1267 (
            .O(N__6715),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1266 (
            .O(N__6712),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1265 (
            .O(N__6709),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1264 (
            .O(N__6702),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__1263 (
            .O(N__6681),
            .I(N__6675));
    InMux I__1262 (
            .O(N__6680),
            .I(N__6675));
    LocalMux I__1261 (
            .O(N__6675),
            .I(\U712_CHIP_RAM.N_396 ));
    InMux I__1260 (
            .O(N__6672),
            .I(N__6669));
    LocalMux I__1259 (
            .O(N__6669),
            .I(N__6666));
    Span4Mux_h I__1258 (
            .O(N__6666),
            .I(N__6661));
    InMux I__1257 (
            .O(N__6665),
            .I(N__6658));
    InMux I__1256 (
            .O(N__6664),
            .I(N__6655));
    Odrv4 I__1255 (
            .O(N__6661),
            .I(\U712_CHIP_RAM.N_400 ));
    LocalMux I__1254 (
            .O(N__6658),
            .I(\U712_CHIP_RAM.N_400 ));
    LocalMux I__1253 (
            .O(N__6655),
            .I(\U712_CHIP_RAM.N_400 ));
    InMux I__1252 (
            .O(N__6648),
            .I(N__6644));
    CascadeMux I__1251 (
            .O(N__6647),
            .I(N__6640));
    LocalMux I__1250 (
            .O(N__6644),
            .I(N__6637));
    InMux I__1249 (
            .O(N__6643),
            .I(N__6633));
    InMux I__1248 (
            .O(N__6640),
            .I(N__6630));
    Span4Mux_h I__1247 (
            .O(N__6637),
            .I(N__6627));
    InMux I__1246 (
            .O(N__6636),
            .I(N__6624));
    LocalMux I__1245 (
            .O(N__6633),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    LocalMux I__1244 (
            .O(N__6630),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    Odrv4 I__1243 (
            .O(N__6627),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    LocalMux I__1242 (
            .O(N__6624),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    CascadeMux I__1241 (
            .O(N__6615),
            .I(N__6611));
    InMux I__1240 (
            .O(N__6614),
            .I(N__6607));
    InMux I__1239 (
            .O(N__6611),
            .I(N__6604));
    CascadeMux I__1238 (
            .O(N__6610),
            .I(N__6601));
    LocalMux I__1237 (
            .O(N__6607),
            .I(N__6596));
    LocalMux I__1236 (
            .O(N__6604),
            .I(N__6596));
    InMux I__1235 (
            .O(N__6601),
            .I(N__6593));
    Span4Mux_h I__1234 (
            .O(N__6596),
            .I(N__6590));
    LocalMux I__1233 (
            .O(N__6593),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    Odrv4 I__1232 (
            .O(N__6590),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    InMux I__1231 (
            .O(N__6585),
            .I(N__6579));
    InMux I__1230 (
            .O(N__6584),
            .I(N__6572));
    InMux I__1229 (
            .O(N__6583),
            .I(N__6572));
    InMux I__1228 (
            .O(N__6582),
            .I(N__6572));
    LocalMux I__1227 (
            .O(N__6579),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__1226 (
            .O(N__6572),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    IoInMux I__1225 (
            .O(N__6567),
            .I(N__6564));
    LocalMux I__1224 (
            .O(N__6564),
            .I(N__6561));
    Span12Mux_s8_h I__1223 (
            .O(N__6561),
            .I(N__6558));
    Span12Mux_v I__1222 (
            .O(N__6558),
            .I(N__6554));
    InMux I__1221 (
            .O(N__6557),
            .I(N__6551));
    Odrv12 I__1220 (
            .O(N__6554),
            .I(TACK_OUTn));
    LocalMux I__1219 (
            .O(N__6551),
            .I(TACK_OUTn));
    CascadeMux I__1218 (
            .O(N__6546),
            .I(N__6543));
    InMux I__1217 (
            .O(N__6543),
            .I(N__6539));
    InMux I__1216 (
            .O(N__6542),
            .I(N__6536));
    LocalMux I__1215 (
            .O(N__6539),
            .I(N__6531));
    LocalMux I__1214 (
            .O(N__6536),
            .I(N__6531));
    Span4Mux_v I__1213 (
            .O(N__6531),
            .I(N__6527));
    InMux I__1212 (
            .O(N__6530),
            .I(N__6524));
    Odrv4 I__1211 (
            .O(N__6527),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__1210 (
            .O(N__6524),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    InMux I__1209 (
            .O(N__6519),
            .I(N__6516));
    LocalMux I__1208 (
            .O(N__6516),
            .I(N__6512));
    InMux I__1207 (
            .O(N__6515),
            .I(N__6509));
    Span4Mux_v I__1206 (
            .O(N__6512),
            .I(N__6506));
    LocalMux I__1205 (
            .O(N__6509),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    Odrv4 I__1204 (
            .O(N__6506),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    InMux I__1203 (
            .O(N__6501),
            .I(N__6493));
    InMux I__1202 (
            .O(N__6500),
            .I(N__6490));
    InMux I__1201 (
            .O(N__6499),
            .I(N__6487));
    InMux I__1200 (
            .O(N__6498),
            .I(N__6484));
    InMux I__1199 (
            .O(N__6497),
            .I(N__6479));
    InMux I__1198 (
            .O(N__6496),
            .I(N__6479));
    LocalMux I__1197 (
            .O(N__6493),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__1196 (
            .O(N__6490),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__1195 (
            .O(N__6487),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__1194 (
            .O(N__6484),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__1193 (
            .O(N__6479),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    InMux I__1192 (
            .O(N__6468),
            .I(N__6464));
    InMux I__1191 (
            .O(N__6467),
            .I(N__6461));
    LocalMux I__1190 (
            .O(N__6464),
            .I(\U712_REG_SM.N_216 ));
    LocalMux I__1189 (
            .O(N__6461),
            .I(\U712_REG_SM.N_216 ));
    InMux I__1188 (
            .O(N__6456),
            .I(N__6448));
    InMux I__1187 (
            .O(N__6455),
            .I(N__6445));
    InMux I__1186 (
            .O(N__6454),
            .I(N__6442));
    InMux I__1185 (
            .O(N__6453),
            .I(N__6435));
    InMux I__1184 (
            .O(N__6452),
            .I(N__6435));
    InMux I__1183 (
            .O(N__6451),
            .I(N__6435));
    LocalMux I__1182 (
            .O(N__6448),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__1181 (
            .O(N__6445),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__1180 (
            .O(N__6442),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__1179 (
            .O(N__6435),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    InMux I__1178 (
            .O(N__6426),
            .I(N__6422));
    InMux I__1177 (
            .O(N__6425),
            .I(N__6419));
    LocalMux I__1176 (
            .O(N__6422),
            .I(\U712_REG_SM.N_239 ));
    LocalMux I__1175 (
            .O(N__6419),
            .I(\U712_REG_SM.N_239 ));
    CascadeMux I__1174 (
            .O(N__6414),
            .I(N__6411));
    InMux I__1173 (
            .O(N__6411),
            .I(N__6406));
    InMux I__1172 (
            .O(N__6410),
            .I(N__6400));
    InMux I__1171 (
            .O(N__6409),
            .I(N__6400));
    LocalMux I__1170 (
            .O(N__6406),
            .I(N__6394));
    InMux I__1169 (
            .O(N__6405),
            .I(N__6387));
    LocalMux I__1168 (
            .O(N__6400),
            .I(N__6384));
    CascadeMux I__1167 (
            .O(N__6399),
            .I(N__6381));
    InMux I__1166 (
            .O(N__6398),
            .I(N__6376));
    InMux I__1165 (
            .O(N__6397),
            .I(N__6376));
    Span4Mux_h I__1164 (
            .O(N__6394),
            .I(N__6373));
    InMux I__1163 (
            .O(N__6393),
            .I(N__6368));
    InMux I__1162 (
            .O(N__6392),
            .I(N__6368));
    InMux I__1161 (
            .O(N__6391),
            .I(N__6363));
    InMux I__1160 (
            .O(N__6390),
            .I(N__6363));
    LocalMux I__1159 (
            .O(N__6387),
            .I(N__6358));
    Span4Mux_h I__1158 (
            .O(N__6384),
            .I(N__6358));
    InMux I__1157 (
            .O(N__6381),
            .I(N__6355));
    LocalMux I__1156 (
            .O(N__6376),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__1155 (
            .O(N__6373),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1154 (
            .O(N__6368),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1153 (
            .O(N__6363),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__1152 (
            .O(N__6358),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1151 (
            .O(N__6355),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    IoInMux I__1150 (
            .O(N__6342),
            .I(N__6339));
    LocalMux I__1149 (
            .O(N__6339),
            .I(N__6335));
    IoInMux I__1148 (
            .O(N__6338),
            .I(N__6332));
    Span4Mux_s2_v I__1147 (
            .O(N__6335),
            .I(N__6329));
    LocalMux I__1146 (
            .O(N__6332),
            .I(N__6326));
    Span4Mux_h I__1145 (
            .O(N__6329),
            .I(N__6323));
    Span4Mux_s2_v I__1144 (
            .O(N__6326),
            .I(N__6320));
    Sp12to4 I__1143 (
            .O(N__6323),
            .I(N__6317));
    Sp12to4 I__1142 (
            .O(N__6320),
            .I(N__6314));
    Span12Mux_h I__1141 (
            .O(N__6317),
            .I(N__6309));
    Span12Mux_h I__1140 (
            .O(N__6314),
            .I(N__6309));
    Odrv12 I__1139 (
            .O(N__6309),
            .I(ASn_c));
    CEMux I__1138 (
            .O(N__6306),
            .I(N__6303));
    LocalMux I__1137 (
            .O(N__6303),
            .I(\U712_REG_SM.N_239_0_0 ));
    InMux I__1136 (
            .O(N__6300),
            .I(N__6295));
    InMux I__1135 (
            .O(N__6299),
            .I(N__6292));
    InMux I__1134 (
            .O(N__6298),
            .I(N__6289));
    LocalMux I__1133 (
            .O(N__6295),
            .I(N__6284));
    LocalMux I__1132 (
            .O(N__6292),
            .I(N__6284));
    LocalMux I__1131 (
            .O(N__6289),
            .I(N__6280));
    Span4Mux_v I__1130 (
            .O(N__6284),
            .I(N__6277));
    InMux I__1129 (
            .O(N__6283),
            .I(N__6274));
    Span4Mux_v I__1128 (
            .O(N__6280),
            .I(N__6271));
    Span4Mux_v I__1127 (
            .O(N__6277),
            .I(N__6266));
    LocalMux I__1126 (
            .O(N__6274),
            .I(N__6266));
    Sp12to4 I__1125 (
            .O(N__6271),
            .I(N__6263));
    Span4Mux_v I__1124 (
            .O(N__6266),
            .I(N__6260));
    Span12Mux_h I__1123 (
            .O(N__6263),
            .I(N__6257));
    Sp12to4 I__1122 (
            .O(N__6260),
            .I(N__6254));
    Span12Mux_v I__1121 (
            .O(N__6257),
            .I(N__6249));
    Span12Mux_h I__1120 (
            .O(N__6254),
            .I(N__6249));
    Odrv12 I__1119 (
            .O(N__6249),
            .I(RnW_c));
    InMux I__1118 (
            .O(N__6246),
            .I(N__6243));
    LocalMux I__1117 (
            .O(N__6243),
            .I(N__6239));
    InMux I__1116 (
            .O(N__6242),
            .I(N__6232));
    Span4Mux_v I__1115 (
            .O(N__6239),
            .I(N__6229));
    InMux I__1114 (
            .O(N__6238),
            .I(N__6226));
    InMux I__1113 (
            .O(N__6237),
            .I(N__6223));
    InMux I__1112 (
            .O(N__6236),
            .I(N__6218));
    InMux I__1111 (
            .O(N__6235),
            .I(N__6218));
    LocalMux I__1110 (
            .O(N__6232),
            .I(N__6214));
    Span4Mux_v I__1109 (
            .O(N__6229),
            .I(N__6209));
    LocalMux I__1108 (
            .O(N__6226),
            .I(N__6209));
    LocalMux I__1107 (
            .O(N__6223),
            .I(N__6206));
    LocalMux I__1106 (
            .O(N__6218),
            .I(N__6203));
    InMux I__1105 (
            .O(N__6217),
            .I(N__6200));
    Span12Mux_s11_v I__1104 (
            .O(N__6214),
            .I(N__6197));
    Span4Mux_v I__1103 (
            .O(N__6209),
            .I(N__6188));
    Span4Mux_v I__1102 (
            .O(N__6206),
            .I(N__6188));
    Span4Mux_h I__1101 (
            .O(N__6203),
            .I(N__6188));
    LocalMux I__1100 (
            .O(N__6200),
            .I(N__6188));
    Odrv12 I__1099 (
            .O(N__6197),
            .I(WRITE_CYCLEm));
    Odrv4 I__1098 (
            .O(N__6188),
            .I(WRITE_CYCLEm));
    IoInMux I__1097 (
            .O(N__6183),
            .I(N__6180));
    LocalMux I__1096 (
            .O(N__6180),
            .I(N__6177));
    IoSpan4Mux I__1095 (
            .O(N__6177),
            .I(N__6174));
    Span4Mux_s3_h I__1094 (
            .O(N__6174),
            .I(N__6171));
    Span4Mux_h I__1093 (
            .O(N__6171),
            .I(N__6168));
    Span4Mux_v I__1092 (
            .O(N__6168),
            .I(N__6165));
    Sp12to4 I__1091 (
            .O(N__6165),
            .I(N__6162));
    Odrv12 I__1090 (
            .O(N__6162),
            .I(N_259));
    InMux I__1089 (
            .O(N__6159),
            .I(N__6151));
    InMux I__1088 (
            .O(N__6158),
            .I(N__6148));
    InMux I__1087 (
            .O(N__6157),
            .I(N__6144));
    InMux I__1086 (
            .O(N__6156),
            .I(N__6141));
    InMux I__1085 (
            .O(N__6155),
            .I(N__6136));
    InMux I__1084 (
            .O(N__6154),
            .I(N__6136));
    LocalMux I__1083 (
            .O(N__6151),
            .I(N__6131));
    LocalMux I__1082 (
            .O(N__6148),
            .I(N__6131));
    InMux I__1081 (
            .O(N__6147),
            .I(N__6128));
    LocalMux I__1080 (
            .O(N__6144),
            .I(N__6123));
    LocalMux I__1079 (
            .O(N__6141),
            .I(N__6123));
    LocalMux I__1078 (
            .O(N__6136),
            .I(\U712_CHIP_RAM.N_360 ));
    Odrv4 I__1077 (
            .O(N__6131),
            .I(\U712_CHIP_RAM.N_360 ));
    LocalMux I__1076 (
            .O(N__6128),
            .I(\U712_CHIP_RAM.N_360 ));
    Odrv4 I__1075 (
            .O(N__6123),
            .I(\U712_CHIP_RAM.N_360 ));
    CEMux I__1074 (
            .O(N__6114),
            .I(N__6111));
    LocalMux I__1073 (
            .O(N__6111),
            .I(N__6108));
    Span4Mux_h I__1072 (
            .O(N__6108),
            .I(N__6105));
    Odrv4 I__1071 (
            .O(N__6105),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0_0 ));
    CascadeMux I__1070 (
            .O(N__6102),
            .I(N__6099));
    InMux I__1069 (
            .O(N__6099),
            .I(N__6096));
    LocalMux I__1068 (
            .O(N__6096),
            .I(\U712_CHIP_RAM.CLK_EN_5_0 ));
    IoInMux I__1067 (
            .O(N__6093),
            .I(N__6090));
    LocalMux I__1066 (
            .O(N__6090),
            .I(N__6087));
    Span4Mux_s3_h I__1065 (
            .O(N__6087),
            .I(N__6084));
    Span4Mux_v I__1064 (
            .O(N__6084),
            .I(N__6081));
    Sp12to4 I__1063 (
            .O(N__6081),
            .I(N__6078));
    Span12Mux_h I__1062 (
            .O(N__6078),
            .I(N__6074));
    InMux I__1061 (
            .O(N__6077),
            .I(N__6071));
    Odrv12 I__1060 (
            .O(N__6074),
            .I(CLK_EN_c));
    LocalMux I__1059 (
            .O(N__6071),
            .I(CLK_EN_c));
    InMux I__1058 (
            .O(N__6066),
            .I(N__6062));
    InMux I__1057 (
            .O(N__6065),
            .I(N__6059));
    LocalMux I__1056 (
            .O(N__6062),
            .I(\U712_CHIP_RAM.N_404 ));
    LocalMux I__1055 (
            .O(N__6059),
            .I(\U712_CHIP_RAM.N_404 ));
    InMux I__1054 (
            .O(N__6054),
            .I(N__6048));
    InMux I__1053 (
            .O(N__6053),
            .I(N__6048));
    LocalMux I__1052 (
            .O(N__6048),
            .I(\U712_CHIP_RAM.N_313_2 ));
    CascadeMux I__1051 (
            .O(N__6045),
            .I(\U712_CHIP_RAM.N_312_cascade_ ));
    CascadeMux I__1050 (
            .O(N__6042),
            .I(N__6037));
    InMux I__1049 (
            .O(N__6041),
            .I(N__6026));
    InMux I__1048 (
            .O(N__6040),
            .I(N__6026));
    InMux I__1047 (
            .O(N__6037),
            .I(N__6023));
    InMux I__1046 (
            .O(N__6036),
            .I(N__6018));
    InMux I__1045 (
            .O(N__6035),
            .I(N__6015));
    CascadeMux I__1044 (
            .O(N__6034),
            .I(N__6008));
    CascadeMux I__1043 (
            .O(N__6033),
            .I(N__6002));
    InMux I__1042 (
            .O(N__6032),
            .I(N__5996));
    InMux I__1041 (
            .O(N__6031),
            .I(N__5996));
    LocalMux I__1040 (
            .O(N__6026),
            .I(N__5992));
    LocalMux I__1039 (
            .O(N__6023),
            .I(N__5989));
    InMux I__1038 (
            .O(N__6022),
            .I(N__5986));
    InMux I__1037 (
            .O(N__6021),
            .I(N__5983));
    LocalMux I__1036 (
            .O(N__6018),
            .I(N__5978));
    LocalMux I__1035 (
            .O(N__6015),
            .I(N__5978));
    InMux I__1034 (
            .O(N__6014),
            .I(N__5975));
    InMux I__1033 (
            .O(N__6013),
            .I(N__5968));
    InMux I__1032 (
            .O(N__6012),
            .I(N__5968));
    InMux I__1031 (
            .O(N__6011),
            .I(N__5968));
    InMux I__1030 (
            .O(N__6008),
            .I(N__5961));
    InMux I__1029 (
            .O(N__6007),
            .I(N__5961));
    InMux I__1028 (
            .O(N__6006),
            .I(N__5961));
    InMux I__1027 (
            .O(N__6005),
            .I(N__5954));
    InMux I__1026 (
            .O(N__6002),
            .I(N__5954));
    InMux I__1025 (
            .O(N__6001),
            .I(N__5954));
    LocalMux I__1024 (
            .O(N__5996),
            .I(N__5951));
    InMux I__1023 (
            .O(N__5995),
            .I(N__5948));
    Odrv4 I__1022 (
            .O(N__5992),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1021 (
            .O(N__5989),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1020 (
            .O(N__5986),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1019 (
            .O(N__5983),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv12 I__1018 (
            .O(N__5978),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1017 (
            .O(N__5975),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1016 (
            .O(N__5968),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1015 (
            .O(N__5961),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1014 (
            .O(N__5954),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1013 (
            .O(N__5951),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1012 (
            .O(N__5948),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    InMux I__1011 (
            .O(N__5925),
            .I(N__5918));
    InMux I__1010 (
            .O(N__5924),
            .I(N__5911));
    InMux I__1009 (
            .O(N__5923),
            .I(N__5911));
    InMux I__1008 (
            .O(N__5922),
            .I(N__5911));
    InMux I__1007 (
            .O(N__5921),
            .I(N__5904));
    LocalMux I__1006 (
            .O(N__5918),
            .I(N__5899));
    LocalMux I__1005 (
            .O(N__5911),
            .I(N__5899));
    InMux I__1004 (
            .O(N__5910),
            .I(N__5896));
    InMux I__1003 (
            .O(N__5909),
            .I(N__5891));
    InMux I__1002 (
            .O(N__5908),
            .I(N__5891));
    InMux I__1001 (
            .O(N__5907),
            .I(N__5888));
    LocalMux I__1000 (
            .O(N__5904),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__999 (
            .O(N__5899),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__998 (
            .O(N__5896),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__997 (
            .O(N__5891),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__996 (
            .O(N__5888),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    InMux I__995 (
            .O(N__5877),
            .I(N__5867));
    InMux I__994 (
            .O(N__5876),
            .I(N__5867));
    InMux I__993 (
            .O(N__5875),
            .I(N__5864));
    InMux I__992 (
            .O(N__5874),
            .I(N__5857));
    InMux I__991 (
            .O(N__5873),
            .I(N__5851));
    InMux I__990 (
            .O(N__5872),
            .I(N__5851));
    LocalMux I__989 (
            .O(N__5867),
            .I(N__5848));
    LocalMux I__988 (
            .O(N__5864),
            .I(N__5845));
    InMux I__987 (
            .O(N__5863),
            .I(N__5840));
    InMux I__986 (
            .O(N__5862),
            .I(N__5840));
    InMux I__985 (
            .O(N__5861),
            .I(N__5835));
    InMux I__984 (
            .O(N__5860),
            .I(N__5835));
    LocalMux I__983 (
            .O(N__5857),
            .I(N__5831));
    InMux I__982 (
            .O(N__5856),
            .I(N__5828));
    LocalMux I__981 (
            .O(N__5851),
            .I(N__5819));
    Span4Mux_h I__980 (
            .O(N__5848),
            .I(N__5819));
    Span4Mux_v I__979 (
            .O(N__5845),
            .I(N__5819));
    LocalMux I__978 (
            .O(N__5840),
            .I(N__5819));
    LocalMux I__977 (
            .O(N__5835),
            .I(N__5816));
    InMux I__976 (
            .O(N__5834),
            .I(N__5813));
    Span4Mux_h I__975 (
            .O(N__5831),
            .I(N__5810));
    LocalMux I__974 (
            .O(N__5828),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__973 (
            .O(N__5819),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__972 (
            .O(N__5816),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__971 (
            .O(N__5813),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__970 (
            .O(N__5810),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    InMux I__969 (
            .O(N__5799),
            .I(N__5794));
    InMux I__968 (
            .O(N__5798),
            .I(N__5790));
    InMux I__967 (
            .O(N__5797),
            .I(N__5786));
    LocalMux I__966 (
            .O(N__5794),
            .I(N__5779));
    CascadeMux I__965 (
            .O(N__5793),
            .I(N__5776));
    LocalMux I__964 (
            .O(N__5790),
            .I(N__5772));
    InMux I__963 (
            .O(N__5789),
            .I(N__5769));
    LocalMux I__962 (
            .O(N__5786),
            .I(N__5766));
    CascadeMux I__961 (
            .O(N__5785),
            .I(N__5763));
    CascadeMux I__960 (
            .O(N__5784),
            .I(N__5757));
    InMux I__959 (
            .O(N__5783),
            .I(N__5752));
    InMux I__958 (
            .O(N__5782),
            .I(N__5752));
    Span4Mux_h I__957 (
            .O(N__5779),
            .I(N__5747));
    InMux I__956 (
            .O(N__5776),
            .I(N__5744));
    InMux I__955 (
            .O(N__5775),
            .I(N__5741));
    Span4Mux_h I__954 (
            .O(N__5772),
            .I(N__5734));
    LocalMux I__953 (
            .O(N__5769),
            .I(N__5734));
    Span4Mux_h I__952 (
            .O(N__5766),
            .I(N__5734));
    InMux I__951 (
            .O(N__5763),
            .I(N__5729));
    InMux I__950 (
            .O(N__5762),
            .I(N__5729));
    InMux I__949 (
            .O(N__5761),
            .I(N__5722));
    InMux I__948 (
            .O(N__5760),
            .I(N__5722));
    InMux I__947 (
            .O(N__5757),
            .I(N__5722));
    LocalMux I__946 (
            .O(N__5752),
            .I(N__5719));
    InMux I__945 (
            .O(N__5751),
            .I(N__5714));
    InMux I__944 (
            .O(N__5750),
            .I(N__5714));
    Odrv4 I__943 (
            .O(N__5747),
            .I(\U712_CHIP_RAM.N_352 ));
    LocalMux I__942 (
            .O(N__5744),
            .I(\U712_CHIP_RAM.N_352 ));
    LocalMux I__941 (
            .O(N__5741),
            .I(\U712_CHIP_RAM.N_352 ));
    Odrv4 I__940 (
            .O(N__5734),
            .I(\U712_CHIP_RAM.N_352 ));
    LocalMux I__939 (
            .O(N__5729),
            .I(\U712_CHIP_RAM.N_352 ));
    LocalMux I__938 (
            .O(N__5722),
            .I(\U712_CHIP_RAM.N_352 ));
    Odrv4 I__937 (
            .O(N__5719),
            .I(\U712_CHIP_RAM.N_352 ));
    LocalMux I__936 (
            .O(N__5714),
            .I(\U712_CHIP_RAM.N_352 ));
    CascadeMux I__935 (
            .O(N__5697),
            .I(N__5693));
    InMux I__934 (
            .O(N__5696),
            .I(N__5688));
    InMux I__933 (
            .O(N__5693),
            .I(N__5685));
    InMux I__932 (
            .O(N__5692),
            .I(N__5680));
    InMux I__931 (
            .O(N__5691),
            .I(N__5677));
    LocalMux I__930 (
            .O(N__5688),
            .I(N__5672));
    LocalMux I__929 (
            .O(N__5685),
            .I(N__5672));
    CascadeMux I__928 (
            .O(N__5684),
            .I(N__5667));
    InMux I__927 (
            .O(N__5683),
            .I(N__5660));
    LocalMux I__926 (
            .O(N__5680),
            .I(N__5657));
    LocalMux I__925 (
            .O(N__5677),
            .I(N__5652));
    Span4Mux_v I__924 (
            .O(N__5672),
            .I(N__5652));
    InMux I__923 (
            .O(N__5671),
            .I(N__5643));
    InMux I__922 (
            .O(N__5670),
            .I(N__5643));
    InMux I__921 (
            .O(N__5667),
            .I(N__5643));
    InMux I__920 (
            .O(N__5666),
            .I(N__5643));
    InMux I__919 (
            .O(N__5665),
            .I(N__5638));
    InMux I__918 (
            .O(N__5664),
            .I(N__5638));
    InMux I__917 (
            .O(N__5663),
            .I(N__5635));
    LocalMux I__916 (
            .O(N__5660),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__915 (
            .O(N__5657),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__914 (
            .O(N__5652),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__913 (
            .O(N__5643),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__912 (
            .O(N__5638),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__911 (
            .O(N__5635),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__910 (
            .O(N__5622),
            .I(N__5619));
    LocalMux I__909 (
            .O(N__5619),
            .I(N__5615));
    InMux I__908 (
            .O(N__5618),
            .I(N__5612));
    Odrv4 I__907 (
            .O(N__5615),
            .I(\U712_REG_SM.N_232 ));
    LocalMux I__906 (
            .O(N__5612),
            .I(\U712_REG_SM.N_232 ));
    CascadeMux I__905 (
            .O(N__5607),
            .I(N__5604));
    InMux I__904 (
            .O(N__5604),
            .I(N__5600));
    InMux I__903 (
            .O(N__5603),
            .I(N__5597));
    LocalMux I__902 (
            .O(N__5600),
            .I(REG_TACK));
    LocalMux I__901 (
            .O(N__5597),
            .I(REG_TACK));
    InMux I__900 (
            .O(N__5592),
            .I(N__5589));
    LocalMux I__899 (
            .O(N__5589),
            .I(\U712_REG_SM.N_289 ));
    InMux I__898 (
            .O(N__5586),
            .I(N__5583));
    LocalMux I__897 (
            .O(N__5583),
            .I(N__5578));
    InMux I__896 (
            .O(N__5582),
            .I(N__5567));
    InMux I__895 (
            .O(N__5581),
            .I(N__5567));
    Span4Mux_h I__894 (
            .O(N__5578),
            .I(N__5564));
    InMux I__893 (
            .O(N__5577),
            .I(N__5561));
    InMux I__892 (
            .O(N__5576),
            .I(N__5558));
    InMux I__891 (
            .O(N__5575),
            .I(N__5555));
    InMux I__890 (
            .O(N__5574),
            .I(N__5552));
    InMux I__889 (
            .O(N__5573),
            .I(N__5547));
    InMux I__888 (
            .O(N__5572),
            .I(N__5547));
    LocalMux I__887 (
            .O(N__5567),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__886 (
            .O(N__5564),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__885 (
            .O(N__5561),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__884 (
            .O(N__5558),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__883 (
            .O(N__5555),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__882 (
            .O(N__5552),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__881 (
            .O(N__5547),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    InMux I__880 (
            .O(N__5532),
            .I(N__5529));
    LocalMux I__879 (
            .O(N__5529),
            .I(N__5526));
    Odrv4 I__878 (
            .O(N__5526),
            .I(\U712_REG_SM.N_254 ));
    CascadeMux I__877 (
            .O(N__5523),
            .I(\U712_REG_SM.N_254_cascade_ ));
    InMux I__876 (
            .O(N__5520),
            .I(N__5517));
    LocalMux I__875 (
            .O(N__5517),
            .I(\U712_REG_SM.N_26 ));
    InMux I__874 (
            .O(N__5514),
            .I(N__5511));
    LocalMux I__873 (
            .O(N__5511),
            .I(N__5507));
    IoInMux I__872 (
            .O(N__5510),
            .I(N__5504));
    Span4Mux_v I__871 (
            .O(N__5507),
            .I(N__5501));
    LocalMux I__870 (
            .O(N__5504),
            .I(N__5498));
    Sp12to4 I__869 (
            .O(N__5501),
            .I(N__5495));
    IoSpan4Mux I__868 (
            .O(N__5498),
            .I(N__5492));
    Span12Mux_h I__867 (
            .O(N__5495),
            .I(N__5489));
    IoSpan4Mux I__866 (
            .O(N__5492),
            .I(N__5486));
    Span12Mux_v I__865 (
            .O(N__5489),
            .I(N__5483));
    IoSpan4Mux I__864 (
            .O(N__5486),
            .I(N__5480));
    Odrv12 I__863 (
            .O(N__5483),
            .I(C1_c));
    Odrv4 I__862 (
            .O(N__5480),
            .I(C1_c));
    InMux I__861 (
            .O(N__5475),
            .I(N__5472));
    LocalMux I__860 (
            .O(N__5472),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    InMux I__859 (
            .O(N__5469),
            .I(N__5466));
    LocalMux I__858 (
            .O(N__5466),
            .I(N__5463));
    Span4Mux_h I__857 (
            .O(N__5463),
            .I(N__5460));
    Odrv4 I__856 (
            .O(N__5460),
            .I(\U712_CHIP_RAM.un3_DMA_CYCLE_START ));
    InMux I__855 (
            .O(N__5457),
            .I(N__5454));
    LocalMux I__854 (
            .O(N__5454),
            .I(\U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_0 ));
    InMux I__853 (
            .O(N__5451),
            .I(N__5448));
    LocalMux I__852 (
            .O(N__5448),
            .I(N__5444));
    InMux I__851 (
            .O(N__5447),
            .I(N__5439));
    Span4Mux_h I__850 (
            .O(N__5444),
            .I(N__5436));
    InMux I__849 (
            .O(N__5443),
            .I(N__5433));
    InMux I__848 (
            .O(N__5442),
            .I(N__5430));
    LocalMux I__847 (
            .O(N__5439),
            .I(\U712_CHIP_RAM.N_207 ));
    Odrv4 I__846 (
            .O(N__5436),
            .I(\U712_CHIP_RAM.N_207 ));
    LocalMux I__845 (
            .O(N__5433),
            .I(\U712_CHIP_RAM.N_207 ));
    LocalMux I__844 (
            .O(N__5430),
            .I(\U712_CHIP_RAM.N_207 ));
    InMux I__843 (
            .O(N__5421),
            .I(N__5418));
    LocalMux I__842 (
            .O(N__5418),
            .I(N__5415));
    Odrv4 I__841 (
            .O(N__5415),
            .I(\U712_CHIP_RAM.CLK_EN_5_0_a2_1_a2_0 ));
    InMux I__840 (
            .O(N__5412),
            .I(N__5409));
    LocalMux I__839 (
            .O(N__5409),
            .I(N__5406));
    Span4Mux_h I__838 (
            .O(N__5406),
            .I(N__5403));
    Odrv4 I__837 (
            .O(N__5403),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0_1 ));
    InMux I__836 (
            .O(N__5400),
            .I(N__5393));
    CascadeMux I__835 (
            .O(N__5399),
            .I(N__5388));
    InMux I__834 (
            .O(N__5398),
            .I(N__5385));
    InMux I__833 (
            .O(N__5397),
            .I(N__5379));
    InMux I__832 (
            .O(N__5396),
            .I(N__5379));
    LocalMux I__831 (
            .O(N__5393),
            .I(N__5376));
    InMux I__830 (
            .O(N__5392),
            .I(N__5370));
    InMux I__829 (
            .O(N__5391),
            .I(N__5370));
    InMux I__828 (
            .O(N__5388),
            .I(N__5367));
    LocalMux I__827 (
            .O(N__5385),
            .I(N__5364));
    InMux I__826 (
            .O(N__5384),
            .I(N__5361));
    LocalMux I__825 (
            .O(N__5379),
            .I(N__5358));
    Span4Mux_h I__824 (
            .O(N__5376),
            .I(N__5355));
    InMux I__823 (
            .O(N__5375),
            .I(N__5352));
    LocalMux I__822 (
            .O(N__5370),
            .I(N__5349));
    LocalMux I__821 (
            .O(N__5367),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__820 (
            .O(N__5364),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__819 (
            .O(N__5361),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__818 (
            .O(N__5358),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__817 (
            .O(N__5355),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__816 (
            .O(N__5352),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__815 (
            .O(N__5349),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    CascadeMux I__814 (
            .O(N__5334),
            .I(N__5328));
    CascadeMux I__813 (
            .O(N__5333),
            .I(N__5324));
    CascadeMux I__812 (
            .O(N__5332),
            .I(N__5321));
    CascadeMux I__811 (
            .O(N__5331),
            .I(N__5318));
    InMux I__810 (
            .O(N__5328),
            .I(N__5315));
    InMux I__809 (
            .O(N__5327),
            .I(N__5312));
    InMux I__808 (
            .O(N__5324),
            .I(N__5307));
    InMux I__807 (
            .O(N__5321),
            .I(N__5307));
    InMux I__806 (
            .O(N__5318),
            .I(N__5304));
    LocalMux I__805 (
            .O(N__5315),
            .I(N__5297));
    LocalMux I__804 (
            .O(N__5312),
            .I(N__5297));
    LocalMux I__803 (
            .O(N__5307),
            .I(N__5297));
    LocalMux I__802 (
            .O(N__5304),
            .I(N__5294));
    Span4Mux_h I__801 (
            .O(N__5297),
            .I(N__5291));
    Odrv4 I__800 (
            .O(N__5294),
            .I(\U712_CHIP_RAM.N_370 ));
    Odrv4 I__799 (
            .O(N__5291),
            .I(\U712_CHIP_RAM.N_370 ));
    InMux I__798 (
            .O(N__5286),
            .I(N__5283));
    LocalMux I__797 (
            .O(N__5283),
            .I(\U712_CHIP_RAM.N_307 ));
    InMux I__796 (
            .O(N__5280),
            .I(N__5277));
    LocalMux I__795 (
            .O(N__5277),
            .I(N__5273));
    InMux I__794 (
            .O(N__5276),
            .I(N__5270));
    Span4Mux_h I__793 (
            .O(N__5273),
            .I(N__5267));
    LocalMux I__792 (
            .O(N__5270),
            .I(\U712_CHIP_RAM.N_411 ));
    Odrv4 I__791 (
            .O(N__5267),
            .I(\U712_CHIP_RAM.N_411 ));
    InMux I__790 (
            .O(N__5262),
            .I(N__5257));
    InMux I__789 (
            .O(N__5261),
            .I(N__5254));
    InMux I__788 (
            .O(N__5260),
            .I(N__5251));
    LocalMux I__787 (
            .O(N__5257),
            .I(N__5248));
    LocalMux I__786 (
            .O(N__5254),
            .I(N__5245));
    LocalMux I__785 (
            .O(N__5251),
            .I(\U712_CHIP_RAM.N_403 ));
    Odrv4 I__784 (
            .O(N__5248),
            .I(\U712_CHIP_RAM.N_403 ));
    Odrv4 I__783 (
            .O(N__5245),
            .I(\U712_CHIP_RAM.N_403 ));
    CascadeMux I__782 (
            .O(N__5238),
            .I(\U712_CHIP_RAM.N_411_cascade_ ));
    InMux I__781 (
            .O(N__5235),
            .I(N__5232));
    LocalMux I__780 (
            .O(N__5232),
            .I(\U712_CHIP_RAM.N_308 ));
    InMux I__779 (
            .O(N__5229),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    InMux I__778 (
            .O(N__5226),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__777 (
            .O(N__5223),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__776 (
            .O(N__5220),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    InMux I__775 (
            .O(N__5217),
            .I(N__5208));
    InMux I__774 (
            .O(N__5216),
            .I(N__5201));
    InMux I__773 (
            .O(N__5215),
            .I(N__5201));
    InMux I__772 (
            .O(N__5214),
            .I(N__5201));
    InMux I__771 (
            .O(N__5213),
            .I(N__5194));
    InMux I__770 (
            .O(N__5212),
            .I(N__5194));
    InMux I__769 (
            .O(N__5211),
            .I(N__5194));
    LocalMux I__768 (
            .O(N__5208),
            .I(\U712_CHIP_RAM.N_49 ));
    LocalMux I__767 (
            .O(N__5201),
            .I(\U712_CHIP_RAM.N_49 ));
    LocalMux I__766 (
            .O(N__5194),
            .I(\U712_CHIP_RAM.N_49 ));
    InMux I__765 (
            .O(N__5187),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    CEMux I__764 (
            .O(N__5184),
            .I(N__5181));
    LocalMux I__763 (
            .O(N__5181),
            .I(N__5177));
    CEMux I__762 (
            .O(N__5180),
            .I(N__5173));
    Span4Mux_h I__761 (
            .O(N__5177),
            .I(N__5170));
    CEMux I__760 (
            .O(N__5176),
            .I(N__5167));
    LocalMux I__759 (
            .O(N__5173),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    Odrv4 I__758 (
            .O(N__5170),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    LocalMux I__757 (
            .O(N__5167),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    InMux I__756 (
            .O(N__5160),
            .I(N__5156));
    InMux I__755 (
            .O(N__5159),
            .I(N__5153));
    LocalMux I__754 (
            .O(N__5156),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__753 (
            .O(N__5153),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__752 (
            .O(N__5148),
            .I(N__5144));
    InMux I__751 (
            .O(N__5147),
            .I(N__5141));
    LocalMux I__750 (
            .O(N__5144),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__749 (
            .O(N__5141),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    CascadeMux I__748 (
            .O(N__5136),
            .I(N__5133));
    InMux I__747 (
            .O(N__5133),
            .I(N__5129));
    InMux I__746 (
            .O(N__5132),
            .I(N__5126));
    LocalMux I__745 (
            .O(N__5129),
            .I(N__5123));
    LocalMux I__744 (
            .O(N__5126),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    Odrv4 I__743 (
            .O(N__5123),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    InMux I__742 (
            .O(N__5118),
            .I(N__5114));
    InMux I__741 (
            .O(N__5117),
            .I(N__5111));
    LocalMux I__740 (
            .O(N__5114),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__739 (
            .O(N__5111),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    CascadeMux I__738 (
            .O(N__5106),
            .I(\U712_CHIP_RAM.N_352_cascade_ ));
    CascadeMux I__737 (
            .O(N__5103),
            .I(\U712_CHIP_RAM.N_328_cascade_ ));
    InMux I__736 (
            .O(N__5100),
            .I(N__5097));
    LocalMux I__735 (
            .O(N__5097),
            .I(\U712_CHIP_RAM.N_323 ));
    InMux I__734 (
            .O(N__5094),
            .I(N__5091));
    LocalMux I__733 (
            .O(N__5091),
            .I(\U712_CHIP_RAM.N_63 ));
    IoInMux I__732 (
            .O(N__5088),
            .I(N__5085));
    LocalMux I__731 (
            .O(N__5085),
            .I(N__5082));
    IoSpan4Mux I__730 (
            .O(N__5082),
            .I(N__5079));
    Span4Mux_s3_v I__729 (
            .O(N__5079),
            .I(N__5076));
    Sp12to4 I__728 (
            .O(N__5076),
            .I(N__5073));
    Span12Mux_s10_v I__727 (
            .O(N__5073),
            .I(N__5070));
    Span12Mux_v I__726 (
            .O(N__5070),
            .I(N__5066));
    InMux I__725 (
            .O(N__5069),
            .I(N__5063));
    Odrv12 I__724 (
            .O(N__5066),
            .I(LATCH_CLK_c));
    LocalMux I__723 (
            .O(N__5063),
            .I(LATCH_CLK_c));
    InMux I__722 (
            .O(N__5058),
            .I(N__5052));
    InMux I__721 (
            .O(N__5057),
            .I(N__5049));
    InMux I__720 (
            .O(N__5056),
            .I(N__5046));
    InMux I__719 (
            .O(N__5055),
            .I(N__5043));
    LocalMux I__718 (
            .O(N__5052),
            .I(N__5040));
    LocalMux I__717 (
            .O(N__5049),
            .I(N__5033));
    LocalMux I__716 (
            .O(N__5046),
            .I(N__5033));
    LocalMux I__715 (
            .O(N__5043),
            .I(N__5033));
    Span4Mux_h I__714 (
            .O(N__5040),
            .I(N__5026));
    Span4Mux_v I__713 (
            .O(N__5033),
            .I(N__5026));
    InMux I__712 (
            .O(N__5032),
            .I(N__5021));
    InMux I__711 (
            .O(N__5031),
            .I(N__5021));
    Odrv4 I__710 (
            .O(N__5026),
            .I(\U712_CHIP_RAM.N_363 ));
    LocalMux I__709 (
            .O(N__5021),
            .I(\U712_CHIP_RAM.N_363 ));
    CascadeMux I__708 (
            .O(N__5016),
            .I(\U712_CHIP_RAM.N_363_cascade_ ));
    InMux I__707 (
            .O(N__5013),
            .I(N__5010));
    LocalMux I__706 (
            .O(N__5010),
            .I(\U712_CHIP_RAM.N_369 ));
    InMux I__705 (
            .O(N__5007),
            .I(N__5001));
    InMux I__704 (
            .O(N__5006),
            .I(N__4996));
    InMux I__703 (
            .O(N__5005),
            .I(N__4996));
    InMux I__702 (
            .O(N__5004),
            .I(N__4993));
    LocalMux I__701 (
            .O(N__5001),
            .I(\U712_CHIP_RAM.N_397 ));
    LocalMux I__700 (
            .O(N__4996),
            .I(\U712_CHIP_RAM.N_397 ));
    LocalMux I__699 (
            .O(N__4993),
            .I(\U712_CHIP_RAM.N_397 ));
    InMux I__698 (
            .O(N__4986),
            .I(N__4983));
    LocalMux I__697 (
            .O(N__4983),
            .I(N__4979));
    InMux I__696 (
            .O(N__4982),
            .I(N__4976));
    Odrv4 I__695 (
            .O(N__4979),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0 ));
    LocalMux I__694 (
            .O(N__4976),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0 ));
    InMux I__693 (
            .O(N__4971),
            .I(N__4968));
    LocalMux I__692 (
            .O(N__4968),
            .I(N__4965));
    Odrv4 I__691 (
            .O(N__4965),
            .I(\U712_CHIP_RAM.N_306 ));
    InMux I__690 (
            .O(N__4962),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__689 (
            .O(N__4959),
            .I(N__4956));
    LocalMux I__688 (
            .O(N__4956),
            .I(N__4953));
    Odrv4 I__687 (
            .O(N__4953),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    InMux I__686 (
            .O(N__4950),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    CascadeMux I__685 (
            .O(N__4947),
            .I(N__4944));
    InMux I__684 (
            .O(N__4944),
            .I(N__4940));
    InMux I__683 (
            .O(N__4943),
            .I(N__4937));
    LocalMux I__682 (
            .O(N__4940),
            .I(\U712_REG_SM.N_255 ));
    LocalMux I__681 (
            .O(N__4937),
            .I(\U712_REG_SM.N_255 ));
    IoInMux I__680 (
            .O(N__4932),
            .I(N__4929));
    LocalMux I__679 (
            .O(N__4929),
            .I(N__4926));
    IoSpan4Mux I__678 (
            .O(N__4926),
            .I(N__4923));
    Span4Mux_s3_h I__677 (
            .O(N__4923),
            .I(N__4920));
    Span4Mux_h I__676 (
            .O(N__4920),
            .I(N__4917));
    Sp12to4 I__675 (
            .O(N__4917),
            .I(N__4913));
    InMux I__674 (
            .O(N__4916),
            .I(N__4910));
    Span12Mux_h I__673 (
            .O(N__4913),
            .I(N__4905));
    LocalMux I__672 (
            .O(N__4910),
            .I(N__4905));
    Span12Mux_h I__671 (
            .O(N__4905),
            .I(N__4902));
    Span12Mux_v I__670 (
            .O(N__4902),
            .I(N__4899));
    Odrv12 I__669 (
            .O(N__4899),
            .I(C3_c));
    InMux I__668 (
            .O(N__4896),
            .I(N__4893));
    LocalMux I__667 (
            .O(N__4893),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    CascadeMux I__666 (
            .O(N__4890),
            .I(N__4887));
    InMux I__665 (
            .O(N__4887),
            .I(N__4884));
    LocalMux I__664 (
            .O(N__4884),
            .I(\U712_REG_SM.STATE_COUNT_srsts_i_0_a2_0_0_0 ));
    InMux I__663 (
            .O(N__4881),
            .I(N__4877));
    InMux I__662 (
            .O(N__4880),
            .I(N__4872));
    LocalMux I__661 (
            .O(N__4877),
            .I(N__4869));
    InMux I__660 (
            .O(N__4876),
            .I(N__4864));
    InMux I__659 (
            .O(N__4875),
            .I(N__4864));
    LocalMux I__658 (
            .O(N__4872),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    Odrv4 I__657 (
            .O(N__4869),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__656 (
            .O(N__4864),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    InMux I__655 (
            .O(N__4857),
            .I(N__4854));
    LocalMux I__654 (
            .O(N__4854),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    InMux I__653 (
            .O(N__4851),
            .I(N__4846));
    InMux I__652 (
            .O(N__4850),
            .I(N__4841));
    InMux I__651 (
            .O(N__4849),
            .I(N__4841));
    LocalMux I__650 (
            .O(N__4846),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__649 (
            .O(N__4841),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    InMux I__648 (
            .O(N__4836),
            .I(N__4833));
    LocalMux I__647 (
            .O(N__4833),
            .I(\U712_REG_SM.N_264 ));
    InMux I__646 (
            .O(N__4830),
            .I(N__4827));
    LocalMux I__645 (
            .O(N__4827),
            .I(\U712_REG_SM.N_24 ));
    CascadeMux I__644 (
            .O(N__4824),
            .I(N__4821));
    InMux I__643 (
            .O(N__4821),
            .I(N__4817));
    CascadeMux I__642 (
            .O(N__4820),
            .I(N__4814));
    LocalMux I__641 (
            .O(N__4817),
            .I(N__4808));
    InMux I__640 (
            .O(N__4814),
            .I(N__4805));
    InMux I__639 (
            .O(N__4813),
            .I(N__4802));
    InMux I__638 (
            .O(N__4812),
            .I(N__4799));
    InMux I__637 (
            .O(N__4811),
            .I(N__4796));
    Odrv4 I__636 (
            .O(N__4808),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__635 (
            .O(N__4805),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__634 (
            .O(N__4802),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__633 (
            .O(N__4799),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__632 (
            .O(N__4796),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    InMux I__631 (
            .O(N__4785),
            .I(N__4782));
    LocalMux I__630 (
            .O(N__4782),
            .I(\U712_CHIP_RAM.N_262 ));
    CascadeMux I__629 (
            .O(N__4779),
            .I(\U712_CHIP_RAM.N_354_cascade_ ));
    InMux I__628 (
            .O(N__4776),
            .I(N__4773));
    LocalMux I__627 (
            .O(N__4773),
            .I(\U712_CHIP_RAM.N_408 ));
    CascadeMux I__626 (
            .O(N__4770),
            .I(\U712_CHIP_RAM.N_408_cascade_ ));
    InMux I__625 (
            .O(N__4767),
            .I(N__4764));
    LocalMux I__624 (
            .O(N__4764),
            .I(N__4759));
    InMux I__623 (
            .O(N__4763),
            .I(N__4756));
    InMux I__622 (
            .O(N__4762),
            .I(N__4753));
    Odrv12 I__621 (
            .O(N__4759),
            .I(\U712_CHIP_RAM.N_359 ));
    LocalMux I__620 (
            .O(N__4756),
            .I(\U712_CHIP_RAM.N_359 ));
    LocalMux I__619 (
            .O(N__4753),
            .I(\U712_CHIP_RAM.N_359 ));
    InMux I__618 (
            .O(N__4746),
            .I(N__4740));
    InMux I__617 (
            .O(N__4745),
            .I(N__4740));
    LocalMux I__616 (
            .O(N__4740),
            .I(\U712_CHIP_RAM.N_305 ));
    CascadeMux I__615 (
            .O(N__4737),
            .I(\U712_CYCLE_TERM.N_236_i_0_en_cascade_ ));
    CEMux I__614 (
            .O(N__4734),
            .I(N__4731));
    LocalMux I__613 (
            .O(N__4731),
            .I(\U712_CYCLE_TERM.N_236_i_0_en_0 ));
    InMux I__612 (
            .O(N__4728),
            .I(N__4725));
    LocalMux I__611 (
            .O(N__4725),
            .I(\U712_REG_SM.STATE_COUNTc_1_0 ));
    CascadeMux I__610 (
            .O(N__4722),
            .I(N__4719));
    InMux I__609 (
            .O(N__4719),
            .I(N__4714));
    InMux I__608 (
            .O(N__4718),
            .I(N__4711));
    InMux I__607 (
            .O(N__4717),
            .I(N__4708));
    LocalMux I__606 (
            .O(N__4714),
            .I(N__4705));
    LocalMux I__605 (
            .O(N__4711),
            .I(N__4702));
    LocalMux I__604 (
            .O(N__4708),
            .I(N__4699));
    Span4Mux_v I__603 (
            .O(N__4705),
            .I(N__4694));
    Span4Mux_h I__602 (
            .O(N__4702),
            .I(N__4689));
    Span4Mux_h I__601 (
            .O(N__4699),
            .I(N__4689));
    InMux I__600 (
            .O(N__4698),
            .I(N__4684));
    InMux I__599 (
            .O(N__4697),
            .I(N__4684));
    Odrv4 I__598 (
            .O(N__4694),
            .I(DBR_SYNCZ0Z_1));
    Odrv4 I__597 (
            .O(N__4689),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__596 (
            .O(N__4684),
            .I(DBR_SYNCZ0Z_1));
    InMux I__595 (
            .O(N__4677),
            .I(N__4674));
    LocalMux I__594 (
            .O(N__4674),
            .I(N__4671));
    Span4Mux_v I__593 (
            .O(N__4671),
            .I(N__4668));
    Span4Mux_v I__592 (
            .O(N__4668),
            .I(N__4665));
    Sp12to4 I__591 (
            .O(N__4665),
            .I(N__4662));
    Odrv12 I__590 (
            .O(N__4662),
            .I(A_c_15));
    InMux I__589 (
            .O(N__4659),
            .I(N__4656));
    LocalMux I__588 (
            .O(N__4656),
            .I(N__4653));
    Span4Mux_v I__587 (
            .O(N__4653),
            .I(N__4650));
    Span4Mux_h I__586 (
            .O(N__4650),
            .I(N__4647));
    Sp12to4 I__585 (
            .O(N__4647),
            .I(N__4644));
    Odrv12 I__584 (
            .O(N__4644),
            .I(A_c_8));
    InMux I__583 (
            .O(N__4641),
            .I(N__4638));
    LocalMux I__582 (
            .O(N__4638),
            .I(N__4635));
    Odrv4 I__581 (
            .O(N__4635),
            .I(\U712_CHIP_RAM.N_217 ));
    InMux I__580 (
            .O(N__4632),
            .I(N__4629));
    LocalMux I__579 (
            .O(N__4629),
            .I(\U712_CHIP_RAM.N_361 ));
    CascadeMux I__578 (
            .O(N__4626),
            .I(\U712_CHIP_RAM.N_217_cascade_ ));
    CascadeMux I__577 (
            .O(N__4623),
            .I(N__4619));
    InMux I__576 (
            .O(N__4622),
            .I(N__4616));
    InMux I__575 (
            .O(N__4619),
            .I(N__4613));
    LocalMux I__574 (
            .O(N__4616),
            .I(\U712_CHIP_RAM.N_222 ));
    LocalMux I__573 (
            .O(N__4613),
            .I(\U712_CHIP_RAM.N_222 ));
    CascadeMux I__572 (
            .O(N__4608),
            .I(N__4602));
    InMux I__571 (
            .O(N__4607),
            .I(N__4599));
    InMux I__570 (
            .O(N__4606),
            .I(N__4592));
    InMux I__569 (
            .O(N__4605),
            .I(N__4592));
    InMux I__568 (
            .O(N__4602),
            .I(N__4592));
    LocalMux I__567 (
            .O(N__4599),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    LocalMux I__566 (
            .O(N__4592),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    CascadeMux I__565 (
            .O(N__4587),
            .I(\U712_CHIP_RAM.N_359_cascade_ ));
    InMux I__564 (
            .O(N__4584),
            .I(N__4580));
    CascadeMux I__563 (
            .O(N__4583),
            .I(N__4577));
    LocalMux I__562 (
            .O(N__4580),
            .I(N__4574));
    InMux I__561 (
            .O(N__4577),
            .I(N__4569));
    Span4Mux_h I__560 (
            .O(N__4574),
            .I(N__4566));
    InMux I__559 (
            .O(N__4573),
            .I(N__4561));
    InMux I__558 (
            .O(N__4572),
            .I(N__4561));
    LocalMux I__557 (
            .O(N__4569),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    Odrv4 I__556 (
            .O(N__4566),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__555 (
            .O(N__4561),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    CascadeMux I__554 (
            .O(N__4554),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15_cascade_ ));
    CascadeMux I__553 (
            .O(N__4551),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_ ));
    InMux I__552 (
            .O(N__4548),
            .I(N__4545));
    LocalMux I__551 (
            .O(N__4545),
            .I(N__4542));
    Sp12to4 I__550 (
            .O(N__4542),
            .I(N__4539));
    Span12Mux_v I__549 (
            .O(N__4539),
            .I(N__4536));
    Span12Mux_h I__548 (
            .O(N__4536),
            .I(N__4533));
    Odrv12 I__547 (
            .O(N__4533),
            .I(A_c_20));
    CascadeMux I__546 (
            .O(N__4530),
            .I(N__4527));
    InMux I__545 (
            .O(N__4527),
            .I(N__4523));
    InMux I__544 (
            .O(N__4526),
            .I(N__4519));
    LocalMux I__543 (
            .O(N__4523),
            .I(N__4516));
    InMux I__542 (
            .O(N__4522),
            .I(N__4511));
    LocalMux I__541 (
            .O(N__4519),
            .I(N__4506));
    Span4Mux_v I__540 (
            .O(N__4516),
            .I(N__4506));
    InMux I__539 (
            .O(N__4515),
            .I(N__4503));
    InMux I__538 (
            .O(N__4514),
            .I(N__4500));
    LocalMux I__537 (
            .O(N__4511),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    Odrv4 I__536 (
            .O(N__4506),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    LocalMux I__535 (
            .O(N__4503),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    LocalMux I__534 (
            .O(N__4500),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    CascadeMux I__533 (
            .O(N__4491),
            .I(\U712_CHIP_RAM.N_330_cascade_ ));
    InMux I__532 (
            .O(N__4488),
            .I(N__4485));
    LocalMux I__531 (
            .O(N__4485),
            .I(N__4482));
    Odrv4 I__530 (
            .O(N__4482),
            .I(\U712_CHIP_RAM.N_331 ));
    CascadeMux I__529 (
            .O(N__4479),
            .I(\U712_CHIP_RAM.BANK0_9_cascade_ ));
    CascadeMux I__528 (
            .O(N__4476),
            .I(N__4472));
    InMux I__527 (
            .O(N__4475),
            .I(N__4469));
    InMux I__526 (
            .O(N__4472),
            .I(N__4466));
    LocalMux I__525 (
            .O(N__4469),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ));
    LocalMux I__524 (
            .O(N__4466),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ));
    IoInMux I__523 (
            .O(N__4461),
            .I(N__4458));
    LocalMux I__522 (
            .O(N__4458),
            .I(N__4455));
    Span4Mux_s3_v I__521 (
            .O(N__4455),
            .I(N__4452));
    Span4Mux_v I__520 (
            .O(N__4452),
            .I(N__4449));
    Span4Mux_v I__519 (
            .O(N__4449),
            .I(N__4445));
    InMux I__518 (
            .O(N__4448),
            .I(N__4442));
    Odrv4 I__517 (
            .O(N__4445),
            .I(BANK0_c));
    LocalMux I__516 (
            .O(N__4442),
            .I(BANK0_c));
    InMux I__515 (
            .O(N__4437),
            .I(N__4434));
    LocalMux I__514 (
            .O(N__4434),
            .I(N__4431));
    Odrv4 I__513 (
            .O(N__4431),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_0 ));
    InMux I__512 (
            .O(N__4428),
            .I(N__4425));
    LocalMux I__511 (
            .O(N__4425),
            .I(\U712_CHIP_RAM.N_16 ));
    CascadeMux I__510 (
            .O(N__4422),
            .I(\U712_CHIP_RAM.N_49_cascade_ ));
    InMux I__509 (
            .O(N__4419),
            .I(N__4416));
    LocalMux I__508 (
            .O(N__4416),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_55_i_a2_0_a2_0_0 ));
    InMux I__507 (
            .O(N__4413),
            .I(N__4410));
    LocalMux I__506 (
            .O(N__4410),
            .I(N__4406));
    InMux I__505 (
            .O(N__4409),
            .I(N__4403));
    Span4Mux_v I__504 (
            .O(N__4406),
            .I(N__4398));
    LocalMux I__503 (
            .O(N__4403),
            .I(N__4395));
    InMux I__502 (
            .O(N__4402),
            .I(N__4392));
    InMux I__501 (
            .O(N__4401),
            .I(N__4389));
    Odrv4 I__500 (
            .O(N__4398),
            .I(REG_CYCLEm));
    Odrv4 I__499 (
            .O(N__4395),
            .I(REG_CYCLEm));
    LocalMux I__498 (
            .O(N__4392),
            .I(REG_CYCLEm));
    LocalMux I__497 (
            .O(N__4389),
            .I(REG_CYCLEm));
    IoInMux I__496 (
            .O(N__4380),
            .I(N__4376));
    IoInMux I__495 (
            .O(N__4379),
            .I(N__4373));
    LocalMux I__494 (
            .O(N__4376),
            .I(N__4370));
    LocalMux I__493 (
            .O(N__4373),
            .I(N__4367));
    Sp12to4 I__492 (
            .O(N__4370),
            .I(N__4364));
    IoSpan4Mux I__491 (
            .O(N__4367),
            .I(N__4361));
    Span12Mux_v I__490 (
            .O(N__4364),
            .I(N__4358));
    Sp12to4 I__489 (
            .O(N__4361),
            .I(N__4355));
    Span12Mux_h I__488 (
            .O(N__4358),
            .I(N__4350));
    Span12Mux_v I__487 (
            .O(N__4355),
            .I(N__4350));
    Odrv12 I__486 (
            .O(N__4350),
            .I(DRDENn_c));
    CascadeMux I__485 (
            .O(N__4347),
            .I(\U712_CHIP_RAM.LATCH_CLK_8_i_0_0_cascade_ ));
    CascadeMux I__484 (
            .O(N__4344),
            .I(\U712_CHIP_RAM.N_368_cascade_ ));
    CascadeMux I__483 (
            .O(N__4341),
            .I(\U712_CHIP_RAM.N_323_cascade_ ));
    CascadeMux I__482 (
            .O(N__4338),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0_cascade_ ));
    InMux I__481 (
            .O(N__4335),
            .I(N__4332));
    LocalMux I__480 (
            .O(N__4332),
            .I(N__4329));
    Span4Mux_v I__479 (
            .O(N__4329),
            .I(N__4326));
    Sp12to4 I__478 (
            .O(N__4326),
            .I(N__4323));
    Span12Mux_h I__477 (
            .O(N__4323),
            .I(N__4320));
    Odrv12 I__476 (
            .O(N__4320),
            .I(A_c_12));
    InMux I__475 (
            .O(N__4317),
            .I(N__4314));
    LocalMux I__474 (
            .O(N__4314),
            .I(N__4311));
    Span12Mux_v I__473 (
            .O(N__4311),
            .I(N__4308));
    Odrv12 I__472 (
            .O(N__4308),
            .I(A_c_5));
    InMux I__471 (
            .O(N__4305),
            .I(N__4302));
    LocalMux I__470 (
            .O(N__4302),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    InMux I__469 (
            .O(N__4299),
            .I(N__4295));
    InMux I__468 (
            .O(N__4298),
            .I(N__4292));
    LocalMux I__467 (
            .O(N__4295),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    LocalMux I__466 (
            .O(N__4292),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    InMux I__465 (
            .O(N__4287),
            .I(N__4284));
    LocalMux I__464 (
            .O(N__4284),
            .I(TACK_EN_i_ess));
    CascadeMux I__463 (
            .O(N__4281),
            .I(\U712_REG_SM.N_294_cascade_ ));
    InMux I__462 (
            .O(N__4278),
            .I(N__4275));
    LocalMux I__461 (
            .O(N__4275),
            .I(N__4271));
    InMux I__460 (
            .O(N__4274),
            .I(N__4268));
    Span4Mux_v I__459 (
            .O(N__4271),
            .I(N__4265));
    LocalMux I__458 (
            .O(N__4268),
            .I(N__4262));
    Sp12to4 I__457 (
            .O(N__4265),
            .I(N__4259));
    Span12Mux_h I__456 (
            .O(N__4262),
            .I(N__4256));
    Span12Mux_h I__455 (
            .O(N__4259),
            .I(N__4253));
    Span12Mux_v I__454 (
            .O(N__4256),
            .I(N__4250));
    Span12Mux_v I__453 (
            .O(N__4253),
            .I(N__4247));
    Odrv12 I__452 (
            .O(N__4250),
            .I(TSn_c));
    Odrv12 I__451 (
            .O(N__4247),
            .I(TSn_c));
    CascadeMux I__450 (
            .O(N__4242),
            .I(N__4239));
    InMux I__449 (
            .O(N__4239),
            .I(N__4236));
    LocalMux I__448 (
            .O(N__4236),
            .I(N__4233));
    Span4Mux_v I__447 (
            .O(N__4233),
            .I(N__4230));
    Sp12to4 I__446 (
            .O(N__4230),
            .I(N__4227));
    Span12Mux_h I__445 (
            .O(N__4227),
            .I(N__4224));
    Span12Mux_v I__444 (
            .O(N__4224),
            .I(N__4221));
    Odrv12 I__443 (
            .O(N__4221),
            .I(REGSPACEn_c));
    InMux I__442 (
            .O(N__4218),
            .I(N__4214));
    InMux I__441 (
            .O(N__4217),
            .I(N__4211));
    LocalMux I__440 (
            .O(N__4214),
            .I(N__4206));
    LocalMux I__439 (
            .O(N__4211),
            .I(N__4206));
    Span12Mux_h I__438 (
            .O(N__4206),
            .I(N__4203));
    Span12Mux_v I__437 (
            .O(N__4203),
            .I(N__4200));
    Odrv12 I__436 (
            .O(N__4200),
            .I(AWEn_c));
    InMux I__435 (
            .O(N__4197),
            .I(N__4192));
    InMux I__434 (
            .O(N__4196),
            .I(N__4187));
    InMux I__433 (
            .O(N__4195),
            .I(N__4187));
    LocalMux I__432 (
            .O(N__4192),
            .I(\U712_CHIP_RAM.N_371 ));
    LocalMux I__431 (
            .O(N__4187),
            .I(\U712_CHIP_RAM.N_371 ));
    IoInMux I__430 (
            .O(N__4182),
            .I(N__4179));
    LocalMux I__429 (
            .O(N__4179),
            .I(N__4176));
    IoSpan4Mux I__428 (
            .O(N__4176),
            .I(N__4173));
    Span4Mux_s2_v I__427 (
            .O(N__4173),
            .I(N__4169));
    CascadeMux I__426 (
            .O(N__4172),
            .I(N__4166));
    Sp12to4 I__425 (
            .O(N__4169),
            .I(N__4163));
    InMux I__424 (
            .O(N__4166),
            .I(N__4160));
    Odrv12 I__423 (
            .O(N__4163),
            .I(DBDIR_c));
    LocalMux I__422 (
            .O(N__4160),
            .I(DBDIR_c));
    CascadeMux I__421 (
            .O(N__4155),
            .I(\U712_CHIP_RAM.N_285_cascade_ ));
    CascadeMux I__420 (
            .O(N__4152),
            .I(\U712_CHIP_RAM.N_309_cascade_ ));
    InMux I__419 (
            .O(N__4149),
            .I(N__4146));
    LocalMux I__418 (
            .O(N__4146),
            .I(\U712_CHIP_RAM.N_311 ));
    CascadeMux I__417 (
            .O(N__4143),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_55_i_a2_0_0_cascade_ ));
    InMux I__416 (
            .O(N__4140),
            .I(N__4134));
    InMux I__415 (
            .O(N__4139),
            .I(N__4127));
    InMux I__414 (
            .O(N__4138),
            .I(N__4127));
    InMux I__413 (
            .O(N__4137),
            .I(N__4127));
    LocalMux I__412 (
            .O(N__4134),
            .I(N__4124));
    LocalMux I__411 (
            .O(N__4127),
            .I(\U712_CHIP_RAM.N_212 ));
    Odrv4 I__410 (
            .O(N__4124),
            .I(\U712_CHIP_RAM.N_212 ));
    CascadeMux I__409 (
            .O(N__4119),
            .I(\U712_CHIP_RAM.N_326_cascade_ ));
    CascadeMux I__408 (
            .O(N__4116),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_cascade_ ));
    CEMux I__407 (
            .O(N__4113),
            .I(N__4110));
    LocalMux I__406 (
            .O(N__4110),
            .I(N__4107));
    Odrv4 I__405 (
            .O(N__4107),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_0 ));
    CascadeMux I__404 (
            .O(N__4104),
            .I(\U712_CHIP_RAM.N_371_cascade_ ));
    CascadeMux I__403 (
            .O(N__4101),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_cascade_ ));
    CEMux I__402 (
            .O(N__4098),
            .I(N__4095));
    LocalMux I__401 (
            .O(N__4095),
            .I(N__4092));
    Span4Mux_v I__400 (
            .O(N__4092),
            .I(N__4089));
    Odrv4 I__399 (
            .O(N__4089),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0 ));
    InMux I__398 (
            .O(N__4086),
            .I(N__4083));
    LocalMux I__397 (
            .O(N__4083),
            .I(\U712_CHIP_RAM.N_321 ));
    InMux I__396 (
            .O(N__4080),
            .I(N__4077));
    LocalMux I__395 (
            .O(N__4077),
            .I(N__4074));
    Span4Mux_v I__394 (
            .O(N__4074),
            .I(N__4071));
    Span4Mux_v I__393 (
            .O(N__4071),
            .I(N__4068));
    Sp12to4 I__392 (
            .O(N__4068),
            .I(N__4065));
    Odrv12 I__391 (
            .O(N__4065),
            .I(A_c_18));
    InMux I__390 (
            .O(N__4062),
            .I(N__4059));
    LocalMux I__389 (
            .O(N__4059),
            .I(N__4056));
    Span4Mux_v I__388 (
            .O(N__4056),
            .I(N__4053));
    Span4Mux_v I__387 (
            .O(N__4053),
            .I(N__4050));
    Sp12to4 I__386 (
            .O(N__4050),
            .I(N__4047));
    Odrv12 I__385 (
            .O(N__4047),
            .I(A_c_16));
    IoInMux I__384 (
            .O(N__4044),
            .I(N__4041));
    LocalMux I__383 (
            .O(N__4041),
            .I(N__4038));
    Span4Mux_s0_h I__382 (
            .O(N__4038),
            .I(N__4035));
    Sp12to4 I__381 (
            .O(N__4035),
            .I(N__4032));
    Span12Mux_v I__380 (
            .O(N__4032),
            .I(N__4029));
    Odrv12 I__379 (
            .O(N__4029),
            .I(N_848_i));
    IoInMux I__378 (
            .O(N__4026),
            .I(N__4023));
    LocalMux I__377 (
            .O(N__4023),
            .I(N__4020));
    Span12Mux_s8_v I__376 (
            .O(N__4020),
            .I(N__4017));
    Odrv12 I__375 (
            .O(N__4017),
            .I(N_336));
    IoInMux I__374 (
            .O(N__4014),
            .I(N__4011));
    LocalMux I__373 (
            .O(N__4011),
            .I(N__4008));
    Span12Mux_s3_v I__372 (
            .O(N__4008),
            .I(N__4005));
    Odrv12 I__371 (
            .O(N__4005),
            .I(VBENn_c));
    CascadeMux I__370 (
            .O(N__4002),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER18_cascade_ ));
    IoInMux I__369 (
            .O(N__3999),
            .I(N__3996));
    LocalMux I__368 (
            .O(N__3996),
            .I(N__3993));
    Span4Mux_s2_v I__367 (
            .O(N__3993),
            .I(N__3990));
    Span4Mux_v I__366 (
            .O(N__3990),
            .I(N__3987));
    Odrv4 I__365 (
            .O(N__3987),
            .I(CLK80_PLL_i_i));
    IoInMux I__364 (
            .O(N__3984),
            .I(N__3981));
    LocalMux I__363 (
            .O(N__3981),
            .I(N__3978));
    IoSpan4Mux I__362 (
            .O(N__3978),
            .I(N__3975));
    Span4Mux_s3_h I__361 (
            .O(N__3975),
            .I(N__3972));
    Odrv4 I__360 (
            .O(N__3972),
            .I(DBRn_c_i_0));
    InMux I__359 (
            .O(N__3969),
            .I(N__3966));
    LocalMux I__358 (
            .O(N__3966),
            .I(N__3963));
    Span4Mux_v I__357 (
            .O(N__3963),
            .I(N__3959));
    InMux I__356 (
            .O(N__3962),
            .I(N__3956));
    Sp12to4 I__355 (
            .O(N__3959),
            .I(N__3951));
    LocalMux I__354 (
            .O(N__3956),
            .I(N__3951));
    Span12Mux_h I__353 (
            .O(N__3951),
            .I(N__3948));
    Span12Mux_v I__352 (
            .O(N__3948),
            .I(N__3945));
    Odrv12 I__351 (
            .O(N__3945),
            .I(DBRn_c));
    InMux I__350 (
            .O(N__3942),
            .I(N__3939));
    LocalMux I__349 (
            .O(N__3939),
            .I(DBR_SYNCZ0Z_0));
    InMux I__348 (
            .O(N__3936),
            .I(N__3933));
    LocalMux I__347 (
            .O(N__3933),
            .I(N__3930));
    Span12Mux_v I__346 (
            .O(N__3930),
            .I(N__3927));
    Span12Mux_v I__345 (
            .O(N__3927),
            .I(N__3924));
    Odrv12 I__344 (
            .O(N__3924),
            .I(RAMSPACEn_c));
    IoInMux I__343 (
            .O(N__3921),
            .I(N__3918));
    LocalMux I__342 (
            .O(N__3918),
            .I(N__3915));
    Span4Mux_s0_v I__341 (
            .O(N__3915),
            .I(N__3912));
    Span4Mux_v I__340 (
            .O(N__3912),
            .I(N__3909));
    Sp12to4 I__339 (
            .O(N__3909),
            .I(N__3906));
    Span12Mux_h I__338 (
            .O(N__3906),
            .I(N__3903));
    Span12Mux_v I__337 (
            .O(N__3903),
            .I(N__3900));
    Odrv12 I__336 (
            .O(N__3900),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .I(N__6864));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .I(N__6862));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .I(N__6863));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .I(N__6861));
    INV \INVU712_CHIP_RAM.DMA_A20C  (
            .O(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .I(N__6860));
    defparam IN_MUX_bfv_10_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_6_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_10_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__7257),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__5510),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB DBRn_c_i_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__3984),
            .GLOBALBUFFEROUTPUT(DBRn_c_i_0_g));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__4932),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_3_1_6.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_3_1_6.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_3_1_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLKRAM_obuf_RNO_LC_3_1_6 (
            .in0(N__8970),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_3_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_3_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_3_10_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_3_10_2  (
            .in0(N__10479),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8648),
            .lcout(DBRn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBRn_ibuf_RNIBAB_LC_5_9_6.C_ON=1'b0;
    defparam DBRn_ibuf_RNIBAB_LC_5_9_6.SEQ_MODE=4'b0000;
    defparam DBRn_ibuf_RNIBAB_LC_5_9_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 DBRn_ibuf_RNIBAB_LC_5_9_6 (
            .in0(N__3962),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DBRn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBR_SYNC_1_LC_6_7_4.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_6_7_4.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_6_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_6_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3942),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8955),
            .ce(),
            .sr(N__10442));
    defparam DBR_SYNC_0_LC_6_8_7.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_6_8_7.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_6_8_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 DBR_SYNC_0_LC_6_8_7 (
            .in0(N__3969),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8956),
            .ce(),
            .sr(N__10434));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_7_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_7_5_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_7_5_0 .LUT_INIT=16'b0101000001110011;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_7_5_0  (
            .in0(N__9378),
            .in1(N__4274),
            .in2(N__4583),
            .in3(N__3936),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8943),
            .ce(),
            .sr(N__10451));
    defparam \U712_CHIP_RAM.DBENn_LC_7_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_7_5_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_7_5_1 .LUT_INIT=16'b0101111111001100;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_7_5_1  (
            .in0(N__10176),
            .in1(N__7693),
            .in2(N__4530),
            .in3(N__4986),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8943),
            .ce(),
            .sr(N__10451));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_7_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_7_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_7_6_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_LC_7_6_0  (
            .in0(N__4698),
            .in1(N__4573),
            .in2(N__5334),
            .in3(N__4526),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8948),
            .ce(N__4113),
            .sr(N__10443));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_7_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_7_6_2 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_7_6_2  (
            .in0(N__4697),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4572),
            .lcout(\U712_CHIP_RAM.N_212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_7_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_7_6_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_7_6_3  (
            .in0(N__9209),
            .in1(N__4080),
            .in2(_gnd_net_),
            .in3(N__4062),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_7_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_7_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_7_7_0 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_7_7_0  (
            .in0(N__4217),
            .in1(N__6298),
            .in2(_gnd_net_),
            .in3(N__5398),
            .lcout(WRITE_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8952),
            .ce(N__4098),
            .sr(N__10435));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_7_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_7_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_7_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4299),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8957),
            .ce(),
            .sr(N__10420));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_7_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_7_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_7_10_2 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_7_10_2  (
            .in0(N__7560),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7836),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8961),
            .ce(),
            .sr(N__10413));
    defparam TACKn_obuft_RNO_LC_7_11_6.C_ON=1'b0;
    defparam TACKn_obuft_RNO_LC_7_11_6.SEQ_MODE=4'b0000;
    defparam TACKn_obuft_RNO_LC_7_11_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 TACKn_obuft_RNO_LC_7_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4287),
            .lcout(N_848_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DMA_LATCH_EN_i_i_a2_LC_7_18_7 .C_ON=1'b0;
    defparam \U712_BUFFERS.DMA_LATCH_EN_i_i_a2_LC_7_18_7 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DMA_LATCH_EN_i_i_a2_LC_7_18_7 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \U712_BUFFERS.DMA_LATCH_EN_i_i_a2_LC_7_18_7  (
            .in0(N__7553),
            .in1(N__7827),
            .in2(_gnd_net_),
            .in3(N__6242),
            .lcout(N_336),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_4_6 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_4_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a2_LC_8_4_6  (
            .in0(N__4413),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9423),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_5_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_5_4  (
            .in0(N__5058),
            .in1(N__6769),
            .in2(N__6042),
            .in3(N__5799),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_5_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_5_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4002),
            .in3(N__5856),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8934),
            .ce(),
            .sr(N__10444));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4HBB7_2_LC_8_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4HBB7_2_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4HBB7_2_LC_8_5_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4HBB7_2_LC_8_5_7  (
            .in0(_gnd_net_),
            .in1(N__4514),
            .in2(_gnd_net_),
            .in3(N__6147),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_8_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_8_6_0 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_8_6_0  (
            .in0(N__4137),
            .in1(N__4195),
            .in2(N__5332),
            .in3(N__4086),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_8_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_8_6_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_8_6_1  (
            .in0(N__10477),
            .in1(_gnd_net_),
            .in2(N__4116),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIGGM16_LC_8_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIGGM16_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIGGM16_LC_8_6_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIGGM16_LC_8_6_2  (
            .in0(N__4139),
            .in1(N__7353),
            .in2(N__5333),
            .in3(N__4196),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_2_LC_8_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_2_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_2_LC_8_6_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_2_LC_8_6_3  (
            .in0(_gnd_net_),
            .in1(N__6755),
            .in2(_gnd_net_),
            .in3(N__6156),
            .lcout(\U712_CHIP_RAM.N_371 ),
            .ltout(\U712_CHIP_RAM.N_371_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIQ6QH5_LC_8_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIQ6QH5_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIQ6QH5_LC_8_6_4 .LUT_INIT=16'b1111000000010000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIQ6QH5_LC_8_6_4  (
            .in0(N__4138),
            .in1(N__6542),
            .in2(N__4104),
            .in3(N__5400),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_8_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_8_6_5 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_8_6_5  (
            .in0(N__10478),
            .in1(_gnd_net_),
            .in2(N__4101),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_8_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_8_6_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_8_6_6  (
            .in0(N__5442),
            .in1(N__5004),
            .in2(_gnd_net_),
            .in3(N__6014),
            .lcout(\U712_CHIP_RAM.N_321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_6_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_6_7  (
            .in0(N__4959),
            .in1(N__7354),
            .in2(N__4476),
            .in3(N__5217),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8944),
            .ce(N__5176),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_8_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_8_7_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_8_7_2  (
            .in0(N__7376),
            .in1(N__5396),
            .in2(N__6546),
            .in3(N__6155),
            .lcout(\U712_CHIP_RAM.N_311 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBDIR_LC_8_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_8_7_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_8_7_4 .LUT_INIT=16'b0111010011110000;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_8_7_4  (
            .in0(N__4218),
            .in1(N__5397),
            .in2(N__4172),
            .in3(N__4197),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8949),
            .ce(),
            .sr(N__10425));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_8_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_8_7_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_8_7_6  (
            .in0(_gnd_net_),
            .in1(N__6768),
            .in2(_gnd_net_),
            .in3(N__6154),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_285_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_7_7 .LUT_INIT=16'b1111101111110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_7_7  (
            .in0(N__4622),
            .in1(N__7377),
            .in2(N__4155),
            .in3(N__5057),
            .lcout(\U712_CHIP_RAM.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_8_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__4776),
            .in2(_gnd_net_),
            .in3(N__5280),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_309_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_8_1 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_8_1  (
            .in0(N__5873),
            .in1(N__5798),
            .in2(N__4152),
            .in3(N__4419),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_55_i_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_8_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_8_8_2 .LUT_INIT=16'b1010101000000011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_8_8_2  (
            .in0(N__9198),
            .in1(N__4149),
            .in2(N__4143),
            .in3(N__4607),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8953),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIHOOI5_LC_8_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIHOOI5_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIHOOI5_LC_8_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIHOOI5_LC_8_8_3  (
            .in0(N__6159),
            .in1(N__7331),
            .in2(N__5331),
            .in3(N__4140),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_326_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI77IM9_LC_8_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI77IM9_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI77IM9_LC_8_8_4 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI77IM9_LC_8_8_4  (
            .in0(N__5412),
            .in1(N__5872),
            .in2(N__4119),
            .in3(N__5797),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI12QHH_2_LC_8_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI12QHH_2_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI12QHH_2_LC_8_8_5 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI12QHH_2_LC_8_8_5  (
            .in0(N__6798),
            .in1(N__4785),
            .in2(N__4338),
            .in3(N__7332),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_8_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_8_8_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_8_8_7  (
            .in0(N__4335),
            .in1(N__4317),
            .in2(_gnd_net_),
            .in3(N__9197),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_8_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_8_9_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__4305),
            .in2(_gnd_net_),
            .in3(N__4298),
            .lcout(\U712_CHIP_RAM.un3_DMA_CYCLE_START ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_10_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_10_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_10_0 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_10_0  (
            .in0(N__7330),
            .in1(N__6614),
            .in2(_gnd_net_),
            .in3(N__6648),
            .lcout(TACK_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8958),
            .ce(N__4734),
            .sr(N__10409));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_8_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_8_11_1 .LUT_INIT=16'b0000111000001111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_8_11_1  (
            .in0(N__6409),
            .in1(N__5577),
            .in2(N__4820),
            .in3(N__4881),
            .lcout(\U712_REG_SM.STATE_COUNTc_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_8_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_8_11_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_0_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(N__4943),
            .in2(_gnd_net_),
            .in3(N__6410),
            .lcout(),
            .ltout(\U712_REG_SM.N_294_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_8_11_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_8_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_8_11_5 .LUT_INIT=16'b1110110011100100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_8_11_5  (
            .in0(N__7281),
            .in1(N__4402),
            .in2(N__4281),
            .in3(N__5532),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8962),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_8_12_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_8_12_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_8_12_1 .LUT_INIT=16'b0011000000110001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_8_12_1  (
            .in0(N__6500),
            .in1(N__5618),
            .in2(N__4890),
            .in3(N__6467),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8963),
            .ce(),
            .sr(N__10401));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_8_12_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_8_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_8_12_4 .LUT_INIT=16'b0101011100000011;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_8_12_4  (
            .in0(N__4401),
            .in1(N__4278),
            .in2(N__4242),
            .in3(N__4851),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8963),
            .ce(),
            .sr(N__10401));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_8_13_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_8_13_7 .LUT_INIT=16'b1010100011111100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_8_13_7  (
            .in0(N__4880),
            .in1(N__5586),
            .in2(N__6414),
            .in3(N__4836),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8966),
            .ce(),
            .sr(N__10400));
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_LC_8_14_1 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_LC_8_14_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_BUFFERS.un1_DRDENn_0_a2_LC_8_14_1  (
            .in0(N__7527),
            .in1(N__7823),
            .in2(_gnd_net_),
            .in3(N__4409),
            .lcout(DRDENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_9_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_9_5_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_0_LC_9_5_0  (
            .in0(_gnd_net_),
            .in1(N__4641),
            .in2(_gnd_net_),
            .in3(N__5006),
            .lcout(\U712_CHIP_RAM.N_331 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_9_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_9_5_1 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_9_5_1  (
            .in0(N__7898),
            .in1(N__5392),
            .in2(_gnd_net_),
            .in3(N__4515),
            .lcout(),
            .ltout(\U712_CHIP_RAM.LATCH_CLK_8_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_9_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_9_5_2 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_9_5_2  (
            .in0(N__5032),
            .in1(N__5789),
            .in2(N__4347),
            .in3(N__6036),
            .lcout(\U712_CHIP_RAM.N_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3FV43_LC_9_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3FV43_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3FV43_LC_9_5_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3FV43_LC_9_5_3  (
            .in0(N__5860),
            .in1(N__5782),
            .in2(_gnd_net_),
            .in3(N__5031),
            .lcout(\U712_CHIP_RAM.N_397 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI7MCB2_LC_9_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI7MCB2_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI7MCB2_LC_9_5_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNI7MCB2_LC_9_5_4  (
            .in0(N__5391),
            .in1(N__6754),
            .in2(_gnd_net_),
            .in3(N__4763),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_368_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIGK316_LC_9_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIGK316_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIGK316_LC_9_5_5 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIGK316_LC_9_5_5  (
            .in0(N__5861),
            .in1(N__5783),
            .in2(N__4344),
            .in3(N__5013),
            .lcout(\U712_CHIP_RAM.N_323 ),
            .ltout(\U712_CHIP_RAM.N_323_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIHBKDA_LC_9_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIHBKDA_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIHBKDA_LC_9_5_6 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIHBKDA_LC_9_5_6  (
            .in0(N__5262),
            .in1(N__6237),
            .in2(N__4341),
            .in3(N__5005),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_9_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_9_6_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_9_6_0  (
            .in0(N__5907),
            .in1(N__5995),
            .in2(_gnd_net_),
            .in3(N__5663),
            .lcout(\U712_CHIP_RAM.N_359 ),
            .ltout(\U712_CHIP_RAM.N_359_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_9_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_9_6_1 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_9_6_1  (
            .in0(N__5751),
            .in1(_gnd_net_),
            .in2(N__4587),
            .in3(N__6746),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER15 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIVLD65_LC_9_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIVLD65_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIVLD65_LC_9_6_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIVLD65_LC_9_6_2  (
            .in0(N__5327),
            .in1(N__4584),
            .in2(N__4554),
            .in3(N__4718),
            .lcout(),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_2_LC_9_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_2_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_2_LC_9_6_3 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_2_LC_9_6_3  (
            .in0(N__10710),
            .in1(_gnd_net_),
            .in2(N__4551),
            .in3(N__4548),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_330_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_9_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_9_6_4 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_1_LC_9_6_4  (
            .in0(N__4522),
            .in1(N__5384),
            .in2(N__4491),
            .in3(N__8628),
            .lcout(),
            .ltout(\U712_CHIP_RAM.BANK0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_LC_9_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.BANK0_LC_9_6_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \U712_CHIP_RAM.BANK0_LC_9_6_5  (
            .in0(N__4488),
            .in1(N__4448),
            .in2(N__4479),
            .in3(N__4475),
            .lcout(BANK0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8935),
            .ce(),
            .sr(N__10426));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI05TJ3_LC_9_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI05TJ3_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI05TJ3_LC_9_6_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI05TJ3_LC_9_6_6  (
            .in0(N__5834),
            .in1(N__4762),
            .in2(_gnd_net_),
            .in3(N__5750),
            .lcout(\U712_CHIP_RAM.N_360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5OHEF_LC_9_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5OHEF_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5OHEF_LC_9_7_0 .LUT_INIT=16'b1111101110111011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5OHEF_LC_9_7_0  (
            .in0(N__4437),
            .in1(N__7375),
            .in2(N__4623),
            .in3(N__5056),
            .lcout(\U712_CHIP_RAM.N_49 ),
            .ltout(\U712_CHIP_RAM.N_49_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_7_1 .LUT_INIT=16'b0101001101011100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_7_1  (
            .in0(N__4428),
            .in1(N__7136),
            .in2(N__4422),
            .in3(N__6005),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8945),
            .ce(N__5180),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_9_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_9_7_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_9_7_2  (
            .in0(N__6742),
            .in1(N__5683),
            .in2(N__6033),
            .in3(N__7374),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_55_i_a2_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_2_LC_9_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_2_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_2_LC_9_7_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_2_LC_9_7_3  (
            .in0(_gnd_net_),
            .in1(N__6740),
            .in2(_gnd_net_),
            .in3(N__6001),
            .lcout(\U712_CHIP_RAM.N_403 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1IJO_LC_9_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1IJO_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1IJO_LC_9_7_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1IJO_LC_9_7_6  (
            .in0(N__6741),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6217),
            .lcout(\U712_CHIP_RAM.N_207 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_8_0 .LUT_INIT=16'b1100000011010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_8_0  (
            .in0(N__5286),
            .in1(N__4605),
            .in2(N__8101),
            .in3(N__5235),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8950),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_8_1 .LUT_INIT=16'b1111000100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_8_1  (
            .in0(N__4746),
            .in1(N__6672),
            .in2(N__4608),
            .in3(N__8346),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8950),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI1DV43_LC_9_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI1DV43_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI1DV43_LC_9_8_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI1DV43_LC_9_8_2  (
            .in0(N__5862),
            .in1(N__6006),
            .in2(N__5784),
            .in3(N__6792),
            .lcout(\U712_CHIP_RAM.N_361 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_8_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_8_3  (
            .in0(N__4677),
            .in1(N__4659),
            .in2(_gnd_net_),
            .in3(N__9199),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI71B91_LC_9_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI71B91_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI71B91_LC_9_8_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNI71B91_LC_9_8_4  (
            .in0(N__7897),
            .in1(N__6007),
            .in2(_gnd_net_),
            .in3(N__5443),
            .lcout(\U712_CHIP_RAM.N_217 ),
            .ltout(\U712_CHIP_RAM.N_217_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIDDEL6_LC_9_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIDDEL6_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIDDEL6_LC_9_8_5 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIDDEL6_LC_9_8_5  (
            .in0(N__4632),
            .in1(N__5760),
            .in2(N__4626),
            .in3(N__5863),
            .lcout(\U712_CHIP_RAM.N_222 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_8_6 .LUT_INIT=16'b1100000011010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_8_6  (
            .in0(N__4971),
            .in1(N__4606),
            .in2(N__8433),
            .in3(N__4745),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8950),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5PDS6_0_LC_9_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5PDS6_0_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5PDS6_0_LC_9_8_7 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI5PDS6_0_LC_9_8_7  (
            .in0(N__5055),
            .in1(N__5761),
            .in2(N__6034),
            .in3(N__6158),
            .lcout(\U712_CHIP_RAM.N_262 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_9_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_9_9_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_9_9_5  (
            .in0(N__6784),
            .in1(N__5925),
            .in2(N__5697),
            .in3(N__6035),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_354_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIFJSJ3_LC_9_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIFJSJ3_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIFJSJ3_LC_9_9_6 .LUT_INIT=16'b0000000011111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIFJSJ3_LC_9_9_6  (
            .in0(N__5696),
            .in1(N__5261),
            .in2(N__4779),
            .in3(N__5875),
            .lcout(\U712_CHIP_RAM.N_408 ),
            .ltout(\U712_CHIP_RAM.N_408_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI997R7_2_LC_9_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI997R7_2_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI997R7_2_LC_9_9_7 .LUT_INIT=16'b1010001010100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI997R7_2_LC_9_9_7  (
            .in0(N__5276),
            .in1(N__6785),
            .in2(N__4770),
            .in3(N__4767),
            .lcout(\U712_CHIP_RAM.N_305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_10_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_10_1 .LUT_INIT=16'b1010101011101010;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_10_1  (
            .in0(N__6519),
            .in1(N__7329),
            .in2(N__6615),
            .in3(N__6636),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_236_i_0_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_10_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_10_2 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_10_2  (
            .in0(N__10474),
            .in1(_gnd_net_),
            .in2(N__4737),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.N_236_i_0_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNITI8N_2_LC_9_10_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNITI8N_2_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNITI8N_2_LC_9_10_4 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNITI8N_2_LC_9_10_4  (
            .in0(N__4812),
            .in1(N__5575),
            .in2(_gnd_net_),
            .in3(N__4717),
            .lcout(\U712_REG_SM.N_255 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_1_LC_9_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_9_11_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_9_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4896),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8959),
            .ce(),
            .sr(N__10402));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_9_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_9_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_9_11_2 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_9_11_2  (
            .in0(N__5581),
            .in1(N__4728),
            .in2(N__4722),
            .in3(N__6398),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8959),
            .ce(),
            .sr(N__10402));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_9_11_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_9_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_9_11_5 .LUT_INIT=16'b1011101100001011;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_9_11_5  (
            .in0(N__6397),
            .in1(N__5582),
            .in2(N__4947),
            .in3(N__6501),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8959),
            .ce(),
            .sr(N__10402));
    defparam \U712_REG_SM.C3_SYNC_0_LC_9_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_9_11_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_9_11_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_9_11_6  (
            .in0(N__4916),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8959),
            .ce(),
            .sr(N__10402));
    defparam \U712_REG_SM.STATE_COUNT_RNIVCF31_1_LC_9_12_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIVCF31_1_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIVCF31_1_LC_9_12_0 .LUT_INIT=16'b1101110011011111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIVCF31_1_LC_9_12_0  (
            .in0(N__6451),
            .in1(N__5572),
            .in2(N__6399),
            .in3(N__4875),
            .lcout(\U712_REG_SM.N_239 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_9_12_1 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_9_12_1 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_0_LC_9_12_1  (
            .in0(N__6299),
            .in1(N__4813),
            .in2(_gnd_net_),
            .in3(N__6453),
            .lcout(\U712_REG_SM.N_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_9_12_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_9_12_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_9_12_2  (
            .in0(N__4850),
            .in1(N__6455),
            .in2(_gnd_net_),
            .in3(N__6498),
            .lcout(\U712_REG_SM.STATE_COUNT_srsts_i_0_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_9_12_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_9_12_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(N__4811),
            .in2(_gnd_net_),
            .in3(N__4876),
            .lcout(\U712_REG_SM.N_232 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_9_12_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_9_12_5 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_9_12_5  (
            .in0(N__6393),
            .in1(N__4857),
            .in2(_gnd_net_),
            .in3(N__4849),
            .lcout(\U712_REG_SM.N_264 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_9_12_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_9_12_6 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_9_12_6  (
            .in0(N__6452),
            .in1(N__5573),
            .in2(_gnd_net_),
            .in3(N__6392),
            .lcout(\U712_REG_SM.N_216 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_LC_9_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DS_EN_LC_9_13_3 .LUT_INIT=16'b0101110101010001;
    LogicCell40 \U712_REG_SM.DS_EN_LC_9_13_3  (
            .in0(N__4830),
            .in1(N__6426),
            .in2(N__4824),
            .in3(N__9863),
            .lcout(DS_ENm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8964),
            .ce(),
            .sr(N__10398));
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_10_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_10_4_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_10_4_5 .LUT_INIT=16'b0000010011111110;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_LC_10_4_5  (
            .in0(N__5100),
            .in1(N__5069),
            .in2(N__6840),
            .in3(N__5094),
            .lcout(LATCH_CLK_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8925),
            .ce(),
            .sr(N__10436));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_10_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_10_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_10_5_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_10_5_1  (
            .in0(_gnd_net_),
            .in1(N__5908),
            .in2(_gnd_net_),
            .in3(N__5664),
            .lcout(\U712_CHIP_RAM.N_363 ),
            .ltout(\U712_CHIP_RAM.N_363_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI4VIE1_LC_10_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI4VIE1_LC_10_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI4VIE1_LC_10_5_2 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNI4VIE1_LC_10_5_2  (
            .in0(_gnd_net_),
            .in1(N__7864),
            .in2(N__5016),
            .in3(N__6031),
            .lcout(\U712_CHIP_RAM.N_369 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_5_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_5_3  (
            .in0(N__9424),
            .in1(N__5909),
            .in2(_gnd_net_),
            .in3(N__5665),
            .lcout(\U712_CHIP_RAM.CLK_EN_5_0_a2_1_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1NGC4_0_LC_10_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1NGC4_0_LC_10_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1NGC4_0_LC_10_5_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI1NGC4_0_LC_10_5_4  (
            .in0(N__5451),
            .in1(N__5007),
            .in2(_gnd_net_),
            .in3(N__6032),
            .lcout(\U712_CHIP_RAM.N_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_5_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_5_6  (
            .in0(_gnd_net_),
            .in1(N__10476),
            .in2(_gnd_net_),
            .in3(N__4982),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_6_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_6_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_6_0  (
            .in0(_gnd_net_),
            .in1(N__6021),
            .in2(_gnd_net_),
            .in3(N__6665),
            .lcout(\U712_CHIP_RAM.N_306 ),
            .ltout(),
            .carryin(bfn_10_6_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_6_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_6_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_6_1  (
            .in0(N__5214),
            .in1(N__5691),
            .in2(_gnd_net_),
            .in3(N__4962),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(N__8929),
            .ce(N__5184),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_6_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_6_2  (
            .in0(_gnd_net_),
            .in1(N__6786),
            .in2(_gnd_net_),
            .in3(N__4950),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_6_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_6_3  (
            .in0(N__5215),
            .in1(N__5921),
            .in2(_gnd_net_),
            .in3(N__5229),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__8929),
            .ce(N__5184),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_6_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_6_4  (
            .in0(N__5211),
            .in1(N__5148),
            .in2(_gnd_net_),
            .in3(N__5226),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__8929),
            .ce(N__5184),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_6_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_6_5  (
            .in0(N__5216),
            .in1(N__5132),
            .in2(_gnd_net_),
            .in3(N__5223),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__8929),
            .ce(N__5184),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_6_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_6_6  (
            .in0(N__5212),
            .in1(N__5160),
            .in2(_gnd_net_),
            .in3(N__5220),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__8929),
            .ce(N__5184),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_6_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_6_7  (
            .in0(N__5118),
            .in1(N__5213),
            .in2(_gnd_net_),
            .in3(N__5187),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8929),
            .ce(N__5184),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_7_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_7_0  (
            .in0(N__5159),
            .in1(N__5147),
            .in2(N__5136),
            .in3(N__5117),
            .lcout(\U712_CHIP_RAM.N_352 ),
            .ltout(\U712_CHIP_RAM.N_352_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3M1M2_LC_10_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3M1M2_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3M1M2_LC_10_7_1 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3M1M2_LC_10_7_1  (
            .in0(N__5666),
            .in1(_gnd_net_),
            .in2(N__5106),
            .in3(N__5874),
            .lcout(\U712_CHIP_RAM.N_396 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_10_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_10_7_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_10_7_2  (
            .in0(N__6065),
            .in1(N__5457),
            .in2(N__9512),
            .in3(N__5775),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_328_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_7_3 .LUT_INIT=16'b1111000111110000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_7_3  (
            .in0(N__5671),
            .in1(N__6236),
            .in2(N__5103),
            .in3(N__9483),
            .lcout(\U712_CHIP_RAM.N_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_7_4 .LUT_INIT=16'b1011100011111000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_7_4  (
            .in0(N__5469),
            .in1(N__7372),
            .in2(N__5399),
            .in3(N__7876),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8936),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_10_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_10_7_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_10_7_5  (
            .in0(N__5670),
            .in1(N__6235),
            .in2(_gnd_net_),
            .in3(N__6012),
            .lcout(\U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_7_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_7_6  (
            .in0(N__6013),
            .in1(N__5447),
            .in2(N__5793),
            .in3(N__5421),
            .lcout(\U712_CHIP_RAM.CLK_EN_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHFLS1_3_LC_10_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHFLS1_3_LC_10_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHFLS1_3_LC_10_7_7 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIHFLS1_3_LC_10_7_7  (
            .in0(N__7373),
            .in1(N__5910),
            .in2(N__5684),
            .in3(N__6011),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIRILU_LC_10_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIRILU_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIRILU_LC_10_8_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIRILU_LC_10_8_0  (
            .in0(_gnd_net_),
            .in1(N__6530),
            .in2(_gnd_net_),
            .in3(N__5375),
            .lcout(\U712_CHIP_RAM.N_370 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_8_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_8_2  (
            .in0(N__6238),
            .in1(N__6664),
            .in2(_gnd_net_),
            .in3(N__6022),
            .lcout(\U712_CHIP_RAM.N_307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_10_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_10_8_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_10_8_3  (
            .in0(N__7342),
            .in1(N__5762),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_411 ),
            .ltout(\U712_CHIP_RAM.N_411_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_8_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_8_4  (
            .in0(N__5924),
            .in1(N__5260),
            .in2(N__5238),
            .in3(N__5877),
            .lcout(\U712_CHIP_RAM.N_308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_10_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_10_8_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_10_8_5  (
            .in0(_gnd_net_),
            .in1(N__6793),
            .in2(_gnd_net_),
            .in3(N__5922),
            .lcout(\U712_CHIP_RAM.N_404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_3_LC_10_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_3_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_3_LC_10_8_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_3_LC_10_8_6  (
            .in0(N__5923),
            .in1(N__5876),
            .in2(N__5785),
            .in3(N__5692),
            .lcout(\U712_CHIP_RAM.N_313_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_9_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_9_5  (
            .in0(N__8337),
            .in1(N__8404),
            .in2(N__8076),
            .in3(N__9235),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_10_9_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_10_9_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN6_LC_10_9_7  (
            .in0(N__6813),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5603),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_LC_10_10_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_10_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_10_10_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_10_10_3  (
            .in0(N__5622),
            .in1(N__5520),
            .in2(N__5607),
            .in3(N__5592),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8954),
            .ce(),
            .sr(N__10403));
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_10_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_10_11_1 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_1_LC_10_11_1  (
            .in0(N__6391),
            .in1(N__5576),
            .in2(_gnd_net_),
            .in3(N__6497),
            .lcout(\U712_REG_SM.N_289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_11_6 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_11_6  (
            .in0(N__6454),
            .in1(N__5574),
            .in2(_gnd_net_),
            .in3(N__6390),
            .lcout(\U712_REG_SM.N_254 ),
            .ltout(\U712_REG_SM.N_254_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_11_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_11_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_10_11_7  (
            .in0(_gnd_net_),
            .in1(N__6300),
            .in2(N__5523),
            .in3(N__6496),
            .lcout(\U712_REG_SM.N_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_1_LC_10_12_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_10_12_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_10_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5475),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8960),
            .ce(),
            .sr(N__10399));
    defparam \U712_REG_SM.C1_SYNC_0_LC_10_12_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_10_12_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_10_12_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_10_12_3  (
            .in0(N__5514),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8960),
            .ce(),
            .sr(N__10399));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_10_12_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_10_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_10_12_4 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_10_12_4  (
            .in0(N__6499),
            .in1(N__6468),
            .in2(_gnd_net_),
            .in3(N__6456),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8960),
            .ce(),
            .sr(N__10399));
    defparam \U712_REG_SM.ASn_ess_RNO_LC_10_13_2 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_10_13_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \U712_REG_SM.ASn_ess_RNO_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(N__10473),
            .in2(_gnd_net_),
            .in3(N__6425),
            .lcout(\U712_REG_SM.N_239_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_ess_LC_10_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_LC_10_14_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_ess_LC_10_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.ASn_ess_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6405),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8965),
            .ce(N__6306),
            .sr(N__10394));
    defparam \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_10_18_6 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_10_18_6 .LUT_INIT=16'b0100000001111111;
    LogicCell40 \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_10_18_6  (
            .in0(N__6283),
            .in1(N__7793),
            .in2(N__7552),
            .in3(N__6246),
            .lcout(N_259),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_11_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_11_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_11_6_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_LC_11_6_0  (
            .in0(_gnd_net_),
            .in1(N__6797),
            .in2(_gnd_net_),
            .in3(N__6157),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8926),
            .ce(N__6114),
            .sr(N__10414));
    defparam \U712_CHIP_RAM.CLK_EN_LC_11_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_11_7_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_11_7_1 .LUT_INIT=16'b0111111100001000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_11_7_1  (
            .in0(N__6054),
            .in1(N__6041),
            .in2(N__6102),
            .in3(N__6077),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8930),
            .ce(),
            .sr(N__10410));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_11_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_11_7_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_11_7_2  (
            .in0(N__6681),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6066),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_312_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_7_3 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_7_3  (
            .in0(N__6053),
            .in1(N__6791),
            .in2(N__6045),
            .in3(N__6040),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_11_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_11_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_11_7_4 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_11_7_4  (
            .in0(N__6812),
            .in1(N__6839),
            .in2(N__6822),
            .in3(N__6819),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8930),
            .ce(),
            .sr(N__10410));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIONRK3_2_LC_11_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIONRK3_2_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIONRK3_2_LC_11_7_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIONRK3_2_LC_11_7_7  (
            .in0(N__7356),
            .in1(N__6790),
            .in2(_gnd_net_),
            .in3(N__6680),
            .lcout(\U712_CHIP_RAM.N_400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_11_8_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_11_8_4 .LUT_INIT=16'b1100100011111000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_11_8_4  (
            .in0(N__7062),
            .in1(N__6584),
            .in2(N__6610),
            .in3(N__6643),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8937),
            .ce(),
            .sr(N__10405));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_11_8_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_11_8_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_11_8_5  (
            .in0(N__6583),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7063),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8937),
            .ce(),
            .sr(N__10405));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_11_8_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_11_8_6 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_11_8_6 .LUT_INIT=16'b0011001100100000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_11_8_6  (
            .in0(N__6945),
            .in1(N__6582),
            .in2(N__6647),
            .in3(N__6515),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8937),
            .ce(),
            .sr(N__10405));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_11_8_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_11_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_11_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6959),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8937),
            .ce(),
            .sr(N__10405));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_11_9_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_11_9_2 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_11_9_2 .LUT_INIT=16'b1111111110100010;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_11_9_2  (
            .in0(N__6557),
            .in1(N__6585),
            .in2(N__7068),
            .in3(N__6974),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8946),
            .ce(),
            .sr(N__10404));
    defparam \U712_CHIP_RAM.REFRESH_LC_11_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_11_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_11_9_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_11_9_4  (
            .in0(N__6896),
            .in1(N__6911),
            .in2(N__6879),
            .in3(N__7152),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8946),
            .ce(),
            .sr(N__10404));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_11_9_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_11_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_11_9_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_11_9_5  (
            .in0(N__6975),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8946),
            .ce(),
            .sr(N__10404));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_10_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_10_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__6939),
            .in2(_gnd_net_),
            .in3(N__6933),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__6859),
            .ce(),
            .sr(N__7194));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_10_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_10_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__6930),
            .in2(_gnd_net_),
            .in3(N__6924),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__6859),
            .ce(),
            .sr(N__7194));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_10_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_10_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(N__7164),
            .in2(_gnd_net_),
            .in3(N__6921),
            .lcout(\U712_CHIP_RAM.REFRESH5lto2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__6859),
            .ce(),
            .sr(N__7194));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_10_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_10_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__7176),
            .in2(_gnd_net_),
            .in3(N__6918),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__6859),
            .ce(),
            .sr(N__7194));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_10_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_10_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(N__7188),
            .in2(_gnd_net_),
            .in3(N__6915),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__6859),
            .ce(),
            .sr(N__7194));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_10_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_10_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(N__6912),
            .in2(_gnd_net_),
            .in3(N__6900),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__6859),
            .ce(),
            .sr(N__7194));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_10_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_10_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__6897),
            .in2(_gnd_net_),
            .in3(N__6885),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__6859),
            .ce(),
            .sr(N__7194));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_10_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_10_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(N__6875),
            .in2(_gnd_net_),
            .in3(N__6882),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6859),
            .ce(),
            .sr(N__7194));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_11_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_11_1  (
            .in0(N__7187),
            .in1(N__7175),
            .in2(_gnd_net_),
            .in3(N__7163),
            .lcout(\U712_CHIP_RAM.REFRESH5lt7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_5_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_5_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_5_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIHMEA_1_LC_12_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIHMEA_1_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIHMEA_1_LC_12_6_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIHMEA_1_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(N__9396),
            .in2(_gnd_net_),
            .in3(N__9273),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_RNIHMEAZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_6_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_6_5  (
            .in0(N__7113),
            .in1(N__9422),
            .in2(_gnd_net_),
            .in3(N__10161),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_231_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_6_6 .LUT_INIT=16'b0011000011111100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_6_6  (
            .in0(_gnd_net_),
            .in1(N__9073),
            .in2(N__7098),
            .in3(N__9274),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_7_0 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_7_0  (
            .in0(N__8137),
            .in1(N__7091),
            .in2(N__9513),
            .in3(N__9950),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_7_7 .LUT_INIT=16'b1111001110111011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_7_7  (
            .in0(N__9951),
            .in1(N__8138),
            .in2(N__7095),
            .in3(N__9487),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pll_RNI8MQ3_LC_12_8_1.C_ON=1'b0;
    defparam pll_RNI8MQ3_LC_12_8_1.SEQ_MODE=4'b0000;
    defparam pll_RNI8MQ3_LC_12_8_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 pll_RNI8MQ3_LC_12_8_1 (
            .in0(N__7067),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK40_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_12_8_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_12_8_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_12_8_2  (
            .in0(_gnd_net_),
            .in1(N__6973),
            .in2(_gnd_net_),
            .in3(N__6960),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_8_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_8_3  (
            .in0(N__9475),
            .in1(N__7446),
            .in2(N__9272),
            .in3(N__10293),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_12_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_12_8_6 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_12_8_6  (
            .in0(N__9250),
            .in1(N__8423),
            .in2(_gnd_net_),
            .in3(N__8089),
            .lcout(\U712_CHIP_RAM.CMA_5_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_12_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_12_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_12_8_7  (
            .in0(N__7437),
            .in1(N__7416),
            .in2(_gnd_net_),
            .in3(N__9251),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_180_i_LC_12_9_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_180_i_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_180_i_LC_12_9_5 .LUT_INIT=16'b0101000101010101;
    LogicCell40 \U712_BYTE_ENABLE.N_180_i_LC_12_9_5  (
            .in0(N__8265),
            .in1(N__7724),
            .in2(N__7832),
            .in3(N__7899),
            .lcout(N_180_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_17_1.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_17_1.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_17_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7355),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_6_5 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_13_6_5  (
            .in0(N__9075),
            .in1(N__9621),
            .in2(N__9031),
            .in3(N__7245),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8927),
            .ce(N__8836),
            .sr(N__10415));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_7_1 .LUT_INIT=16'b0011001100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_7_1  (
            .in0(N__8760),
            .in1(N__9279),
            .in2(N__9516),
            .in3(N__9074),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_13_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_13_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_13_7_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_13_7_2  (
            .in0(_gnd_net_),
            .in1(N__7656),
            .in2(N__7215),
            .in3(N__7605),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8931),
            .ce(N__8815),
            .sr(N__10411));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_13_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_13_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_13_7_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_13_7_3  (
            .in0(_gnd_net_),
            .in1(N__8437),
            .in2(_gnd_net_),
            .in3(N__8097),
            .lcout(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ),
            .ltout(\U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_7_4 .LUT_INIT=16'b0101111101011101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_7_4  (
            .in0(N__9278),
            .in1(N__8759),
            .in2(N__7659),
            .in3(N__9494),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_13_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_13_7_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_13_7_7  (
            .in0(N__7650),
            .in1(N__7644),
            .in2(_gnd_net_),
            .in3(N__7638),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8931),
            .ce(N__8815),
            .sr(N__10411));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_13_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_13_8_0 .LUT_INIT=16'b0001001000010011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_13_8_0  (
            .in0(N__8422),
            .in1(N__8347),
            .in2(N__9244),
            .in3(N__8093),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_8_2 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_8_2  (
            .in0(N__9214),
            .in1(N__7611),
            .in2(N__9511),
            .in3(N__9549),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_8_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_8_3  (
            .in0(N__7599),
            .in1(N__7578),
            .in2(_gnd_net_),
            .in3(N__9213),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_13_9_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_13_9_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_LC_13_9_3  (
            .in0(N__7725),
            .in1(N__7550),
            .in2(_gnd_net_),
            .in3(N__7900),
            .lcout(\U712_BYTE_ENABLE.N_342 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_LC_13_9_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_LC_13_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_LC_13_9_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_LC_13_9_7  (
            .in0(N__7726),
            .in1(N__7551),
            .in2(_gnd_net_),
            .in3(N__7901),
            .lcout(\U712_BYTE_ENABLE.N_320 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_LC_13_10_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_LC_13_10_4 .LUT_INIT=16'b1000101000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_LC_13_10_4  (
            .in0(N__8594),
            .in1(N__9851),
            .in2(N__9759),
            .in3(N__9503),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_341_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_55_i_LC_13_10_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_55_i_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_55_i_LC_13_10_5 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \U712_BYTE_ENABLE.N_55_i_LC_13_10_5  (
            .in0(N__9502),
            .in1(N__7476),
            .in2(N__7470),
            .in3(N__8285),
            .lcout(N_55_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_13_10_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_13_10_6 .LUT_INIT=16'b0000110100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_13_10_6  (
            .in0(N__9758),
            .in1(N__9852),
            .in2(N__8598),
            .in3(N__9504),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_318_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_105_i_LC_13_10_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_105_i_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_105_i_LC_13_10_7 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \U712_BYTE_ENABLE.N_105_i_LC_13_10_7  (
            .in0(N__9501),
            .in1(N__8010),
            .in2(N__8004),
            .in3(N__8284),
            .lcout(N_105_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_x2_LC_13_18_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_x2_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_x2_LC_13_18_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_x2_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(N__9743),
            .in2(_gnd_net_),
            .in3(N__8516),
            .lcout(\U712_BYTE_ENABLE.N_206_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_14_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_14_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_14_6_3 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_14_6_3  (
            .in0(N__9084),
            .in1(N__9633),
            .in2(N__9042),
            .in3(N__7917),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8932),
            .ce(N__8835),
            .sr(N__10421));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_14_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_14_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_14_7_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_14_7_6  (
            .in0(N__10475),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7959),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_14_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_14_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_14_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_14_8_4  (
            .in0(N__7953),
            .in1(N__7938),
            .in2(_gnd_net_),
            .in3(N__9280),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_14_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_14_8_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_14_8_5  (
            .in0(N__9281),
            .in1(N__9476),
            .in2(N__7920),
            .in3(N__10254),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_14_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_14_8_7 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_14_8_7  (
            .in0(N__9282),
            .in1(N__7908),
            .in2(N__9517),
            .in3(N__9912),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_57_i_LC_14_9_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_57_i_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_57_i_LC_14_9_0 .LUT_INIT=16'b0011001100110001;
    LogicCell40 \U712_BYTE_ENABLE.N_57_i_LC_14_9_0  (
            .in0(N__7902),
            .in1(N__8301),
            .in2(N__7831),
            .in3(N__7733),
            .lcout(N_57_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_14_10_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_14_10_0 .LUT_INIT=16'b0100000011110000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_14_10_0  (
            .in0(N__9849),
            .in1(N__8592),
            .in2(N__9518),
            .in3(N__8294),
            .lcout(\U712_BYTE_ENABLE.N_339 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_14_10_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_14_10_4 .LUT_INIT=16'b0001000011110000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_14_10_4  (
            .in0(N__9850),
            .in1(N__8593),
            .in2(N__9519),
            .in3(N__8295),
            .lcout(\U712_BYTE_ENABLE.N_316 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_277_i_LC_14_20_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_277_i_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_277_i_LC_14_20_3 .LUT_INIT=16'b0101010010101000;
    LogicCell40 \U712_BYTE_ENABLE.N_277_i_LC_14_20_3  (
            .in0(N__9733),
            .in1(N__9833),
            .in2(N__8581),
            .in3(N__8495),
            .lcout(N_277_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LLBE_i_o2_i_LC_14_20_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LLBE_i_o2_i_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LLBE_i_o2_i_LC_14_20_4 .LUT_INIT=16'b0000011100110000;
    LogicCell40 \U712_BYTE_ENABLE.LLBE_i_o2_i_LC_14_20_4  (
            .in0(N__9832),
            .in1(N__8570),
            .in2(N__8505),
            .in3(N__9732),
            .lcout(LLBE_i_o2_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WEn_LC_15_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_15_4_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_15_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_15_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8103),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8928),
            .ce(),
            .sr(N__10445));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_15_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_15_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_15_6_6 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_15_6_6  (
            .in0(N__8147),
            .in1(N__8205),
            .in2(N__9515),
            .in3(N__9642),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8938),
            .ce(N__8837),
            .sr(N__10427));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_15_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_15_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_15_6_7 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_15_6_7  (
            .in0(N__8166),
            .in1(N__8769),
            .in2(N__9514),
            .in3(N__8148),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8938),
            .ce(N__8837),
            .sr(N__10427));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_15_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_15_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_15_7_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_15_7_5  (
            .in0(N__8444),
            .in1(N__9294),
            .in2(N__8361),
            .in3(N__8102),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8947),
            .ce(N__8831),
            .sr(N__10422));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_15_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_15_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_15_7_6 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_15_7_6  (
            .in0(N__9085),
            .in1(N__9918),
            .in2(N__9043),
            .in3(N__8733),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8947),
            .ce(N__8831),
            .sr(N__10422));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_15_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_15_8_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_15_8_3  (
            .in0(N__9473),
            .in1(N__8706),
            .in2(N__9295),
            .in3(N__10098),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_15_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_15_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_15_8_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_15_8_5  (
            .in0(N__8694),
            .in1(N__8676),
            .in2(_gnd_net_),
            .in3(N__9283),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_15_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_15_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_15_8_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_15_8_6  (
            .in0(N__9284),
            .in1(N__9474),
            .in2(N__8655),
            .in3(N__10146),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_A20_LC_15_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A20_LC_15_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A20_LC_15_9_1 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_A20_LC_15_9_1  (
            .in0(N__8652),
            .in1(N__10680),
            .in2(N__10766),
            .in3(N__8624),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .ce(),
            .sr(N__10412));
    defparam \U712_BYTE_ENABLE.UMBE_0_LC_15_19_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UMBE_0_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UMBE_0_LC_15_19_2 .LUT_INIT=16'b0000101110100000;
    LogicCell40 \U712_BYTE_ENABLE.UMBE_0_LC_15_19_2  (
            .in0(N__8544),
            .in1(N__9834),
            .in2(N__8520),
            .in3(N__9749),
            .lcout(UMBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_276_i_LC_15_20_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_276_i_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_276_i_LC_15_20_4 .LUT_INIT=16'b0101000110100010;
    LogicCell40 \U712_BYTE_ENABLE.N_276_i_LC_15_20_4  (
            .in0(N__9747),
            .in1(N__8574),
            .in2(N__9848),
            .in3(N__8515),
            .lcout(N_276_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RASn_LC_16_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_16_4_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_16_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_16_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8445),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8933),
            .ce(),
            .sr(N__10452));
    defparam \U712_CHIP_RAM.CRCSn_LC_16_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_16_4_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_16_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_16_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8357),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8933),
            .ce(),
            .sr(N__10452));
    defparam \U712_CHIP_RAM.CASn_LC_16_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_16_5_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_16_5_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_16_5_1  (
            .in0(N__9299),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8939),
            .ce(),
            .sr(N__10446));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_16_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_16_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_16_6_6 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_16_6_6  (
            .in0(N__9472),
            .in1(N__9312),
            .in2(N__9300),
            .in3(N__10521),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_16_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_16_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_16_7_2 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_16_7_2  (
            .in0(N__9094),
            .in1(N__10038),
            .in2(N__9044),
            .in3(N__9141),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8951),
            .ce(N__8841),
            .sr(N__10428));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_16_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_16_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_16_7_6 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_16_7_6  (
            .in0(N__9095),
            .in1(N__9609),
            .in2(N__9045),
            .in3(N__9120),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8951),
            .ce(N__8841),
            .sr(N__10428));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_16_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_16_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_16_7_7 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_16_7_7  (
            .in0(N__9096),
            .in1(N__9041),
            .in2(N__8742),
            .in3(N__8994),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8951),
            .ce(N__8841),
            .sr(N__10428));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_16_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_16_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_16_8_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_16_8_0  (
            .in0(N__10767),
            .in1(N__10660),
            .in2(_gnd_net_),
            .in3(N__8781),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9934),
            .ce(N__10503),
            .sr(N__10423));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_16_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_16_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_16_8_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_16_8_1  (
            .in0(N__10245),
            .in1(_gnd_net_),
            .in2(N__10693),
            .in3(N__9603),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9934),
            .ce(N__10503),
            .sr(N__10423));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_16_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_16_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_16_8_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_16_8_3  (
            .in0(N__10026),
            .in1(_gnd_net_),
            .in2(N__10694),
            .in3(N__10133),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9934),
            .ce(N__10503),
            .sr(N__10423));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_16_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_16_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_16_8_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_16_8_4  (
            .in0(N__10200),
            .in1(N__10653),
            .in2(_gnd_net_),
            .in3(N__10244),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9934),
            .ce(N__10503),
            .sr(N__10423));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_16_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_16_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_16_9_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_16_9_3  (
            .in0(N__9597),
            .in1(N__10679),
            .in2(_gnd_net_),
            .in3(N__10235),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__10502),
            .sr(N__10416));
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_16_19_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_16_19_3 .LUT_INIT=16'b0100010011111111;
    LogicCell40 \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_16_19_3  (
            .in0(N__9830),
            .in1(N__9712),
            .in2(_gnd_net_),
            .in3(N__9881),
            .lcout(un1_LDSn_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_16_20_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_16_20_2 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_16_20_2  (
            .in0(N__9882),
            .in1(N__9831),
            .in2(_gnd_net_),
            .in3(N__9748),
            .lcout(N_87),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_17_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_17_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_17_6_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_17_6_0  (
            .in0(N__10554),
            .in1(N__10703),
            .in2(_gnd_net_),
            .in3(N__10753),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9936),
            .ce(N__10509),
            .sr(N__10447));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_17_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_17_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_17_7_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_17_7_2  (
            .in0(N__9599),
            .in1(N__10688),
            .in2(_gnd_net_),
            .in3(N__10283),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9935),
            .ce(N__10507),
            .sr(N__10437));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_17_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_17_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_17_7_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_17_7_3  (
            .in0(N__10284),
            .in1(_gnd_net_),
            .in2(N__10708),
            .in3(N__10084),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9935),
            .ce(N__10507),
            .sr(N__10437));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_7_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_7_7  (
            .in0(N__10692),
            .in1(N__10553),
            .in2(_gnd_net_),
            .in3(N__10134),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9935),
            .ce(N__10507),
            .sr(N__10437));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_17_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_17_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_17_8_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_17_8_2  (
            .in0(N__10276),
            .in1(N__10697),
            .in2(_gnd_net_),
            .in3(N__9598),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__10505),
            .sr(N__10429));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_17_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_17_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_17_8_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_17_8_3  (
            .in0(N__10086),
            .in1(_gnd_net_),
            .in2(N__10709),
            .in3(N__9984),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__10505),
            .sr(N__10429));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_17_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_17_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_17_8_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_17_8_4  (
            .in0(N__10277),
            .in1(N__10698),
            .in2(_gnd_net_),
            .in3(N__10085),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__10505),
            .sr(N__10429));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_17_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_17_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_17_8_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_17_8_5  (
            .in0(N__10696),
            .in1(N__10234),
            .in2(_gnd_net_),
            .in3(N__10199),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__10505),
            .sr(N__10429));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_17_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_17_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_17_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_17_8_6  (
            .in0(N__10132),
            .in1(N__10022),
            .in2(_gnd_net_),
            .in3(N__10702),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__10505),
            .sr(N__10429));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_17_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_17_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_17_9_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_17_9_0  (
            .in0(N__10020),
            .in1(N__10661),
            .in2(_gnd_net_),
            .in3(N__9980),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__10504),
            .sr(N__10424));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_17_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_17_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_17_9_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_17_9_3  (
            .in0(N__10546),
            .in1(_gnd_net_),
            .in2(N__10695),
            .in3(N__10131),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__10504),
            .sr(N__10424));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_18_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_18_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_18_8_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_18_8_1  (
            .in0(N__9978),
            .in1(N__10684),
            .in2(_gnd_net_),
            .in3(N__10075),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9933),
            .ce(N__10508),
            .sr(N__10438));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_18_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_18_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_18_8_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_18_8_2  (
            .in0(N__10021),
            .in1(_gnd_net_),
            .in2(N__10707),
            .in3(N__9979),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9933),
            .ce(N__10508),
            .sr(N__10438));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_18_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_18_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_18_9_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_18_9_0  (
            .in0(N__10744),
            .in1(N__10621),
            .in2(_gnd_net_),
            .in3(N__10537),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .ce(N__10506),
            .sr(N__10430));
endmodule // U712_TOP

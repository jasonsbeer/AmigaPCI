----------------------------------------------------------------------------------
--This work is shared under the Attribution-NonCommercial-ShareAlike 4.0 International (CC BY-NC-SA 4.0) License
--https://creativecommons.org/licenses/by-nc-sa/4.0/legalcode
	
--You are free to:
--Share - copy and redistribute the material in any medium or format
--Adapt - remix, transform, and build upon the material

--Under the following terms:

--Attribution - You must give appropriate credit, provide a link to the license, and indicate if changes were made. 
--You may do so in any reasonable manner, but not in any way that suggests the licensor endorses you or your use.

--NonCommercial - You may not use the material for commercial purposes.

--ShareAlike - If you remix, transform, or build upon the material, you must distribute your contributions under the 
--same license as the original.

--No additional restrictions - You may not apply legal terms or technological measures that legally restrict others 
--from doing anything the license permits.
--------------------------------------------------------------------------------------------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity C4Clock is
    Port ( 
      
		VCDAC : IN  STD_LOGIC;
      VC3 : IN  STD_LOGIC;
		
      C4 : OUT  STD_LOGIC
		
    );
	 
end C4Clock;

architecture Behavioral of C4Clock is

begin

   --------------
   -- C4 CLOCK --
	--------------
	
	--C4 IS A CLOCK GENERATED BY GARY IN THE A2000 AND SIMPLE FF IN THE A3000.
	--IT IS CONSUMED BY VIDEO DEVICES ON THE VIDEO SLOT.
	
	PROCESS (VCDAC) BEGIN
	
		IF RISING_EDGE (VCDAC) THEN
		
			C4 <= VC3;
			
		END IF;
		
	END PROCESS;


end Behavioral;


// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Sep 14 2025 10:30:51

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    SIZ,
    DRA,
    CMA,
    DA,
    A,
    TBIn,
    RAMSPACEn,
    DBRn,
    RAMENn,
    TSn,
    LMBEn,
    DMA_LATCH_EN,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    UUBEn,
    LDSn,
    LATCH_CLK,
    CASUn,
    RAS1n,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    UMBEn,
    RAS0n,
    PRnW,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    BLSn,
    TCIn,
    WEn,
    REGENn,
    LLBEn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    input [1:0] SIZ;
    input [9:0] DRA;
    output [10:0] CMA;
    output [2:0] DA;
    input [20:0] A;
    output TBIn;
    input RAMSPACEn;
    input DBRn;
    output RAMENn;
    input TSn;
    output LMBEn;
    output DMA_LATCH_EN;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output UUBEn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    input RAS1n;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    output UMBEn;
    input RAS0n;
    output PRnW;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    output BLSn;
    output TCIn;
    output WEn;
    output REGENn;
    output LLBEn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__13161;
    wire N__13160;
    wire N__13159;
    wire N__13152;
    wire N__13151;
    wire N__13150;
    wire N__13143;
    wire N__13142;
    wire N__13141;
    wire N__13134;
    wire N__13133;
    wire N__13132;
    wire N__13125;
    wire N__13124;
    wire N__13123;
    wire N__13116;
    wire N__13115;
    wire N__13114;
    wire N__13107;
    wire N__13106;
    wire N__13105;
    wire N__13098;
    wire N__13097;
    wire N__13096;
    wire N__13089;
    wire N__13088;
    wire N__13087;
    wire N__13080;
    wire N__13079;
    wire N__13078;
    wire N__13071;
    wire N__13070;
    wire N__13069;
    wire N__13062;
    wire N__13061;
    wire N__13060;
    wire N__13053;
    wire N__13052;
    wire N__13051;
    wire N__13044;
    wire N__13043;
    wire N__13042;
    wire N__13035;
    wire N__13034;
    wire N__13033;
    wire N__13026;
    wire N__13025;
    wire N__13024;
    wire N__13017;
    wire N__13016;
    wire N__13015;
    wire N__13008;
    wire N__13007;
    wire N__13006;
    wire N__12999;
    wire N__12998;
    wire N__12997;
    wire N__12990;
    wire N__12989;
    wire N__12988;
    wire N__12981;
    wire N__12980;
    wire N__12979;
    wire N__12972;
    wire N__12971;
    wire N__12970;
    wire N__12963;
    wire N__12962;
    wire N__12961;
    wire N__12954;
    wire N__12953;
    wire N__12952;
    wire N__12945;
    wire N__12944;
    wire N__12943;
    wire N__12936;
    wire N__12935;
    wire N__12934;
    wire N__12927;
    wire N__12926;
    wire N__12925;
    wire N__12918;
    wire N__12917;
    wire N__12916;
    wire N__12909;
    wire N__12908;
    wire N__12907;
    wire N__12900;
    wire N__12899;
    wire N__12898;
    wire N__12891;
    wire N__12890;
    wire N__12889;
    wire N__12882;
    wire N__12881;
    wire N__12880;
    wire N__12873;
    wire N__12872;
    wire N__12871;
    wire N__12864;
    wire N__12863;
    wire N__12862;
    wire N__12855;
    wire N__12854;
    wire N__12853;
    wire N__12846;
    wire N__12845;
    wire N__12844;
    wire N__12837;
    wire N__12836;
    wire N__12835;
    wire N__12828;
    wire N__12827;
    wire N__12826;
    wire N__12819;
    wire N__12818;
    wire N__12817;
    wire N__12810;
    wire N__12809;
    wire N__12808;
    wire N__12801;
    wire N__12800;
    wire N__12799;
    wire N__12792;
    wire N__12791;
    wire N__12790;
    wire N__12783;
    wire N__12782;
    wire N__12781;
    wire N__12774;
    wire N__12773;
    wire N__12772;
    wire N__12765;
    wire N__12764;
    wire N__12763;
    wire N__12756;
    wire N__12755;
    wire N__12754;
    wire N__12747;
    wire N__12746;
    wire N__12745;
    wire N__12738;
    wire N__12737;
    wire N__12736;
    wire N__12729;
    wire N__12728;
    wire N__12727;
    wire N__12720;
    wire N__12719;
    wire N__12718;
    wire N__12711;
    wire N__12710;
    wire N__12709;
    wire N__12702;
    wire N__12701;
    wire N__12700;
    wire N__12693;
    wire N__12692;
    wire N__12691;
    wire N__12684;
    wire N__12683;
    wire N__12682;
    wire N__12675;
    wire N__12674;
    wire N__12673;
    wire N__12666;
    wire N__12665;
    wire N__12664;
    wire N__12657;
    wire N__12656;
    wire N__12655;
    wire N__12648;
    wire N__12647;
    wire N__12646;
    wire N__12639;
    wire N__12638;
    wire N__12637;
    wire N__12630;
    wire N__12629;
    wire N__12628;
    wire N__12621;
    wire N__12620;
    wire N__12619;
    wire N__12612;
    wire N__12611;
    wire N__12610;
    wire N__12603;
    wire N__12602;
    wire N__12601;
    wire N__12594;
    wire N__12593;
    wire N__12592;
    wire N__12585;
    wire N__12584;
    wire N__12583;
    wire N__12576;
    wire N__12575;
    wire N__12574;
    wire N__12567;
    wire N__12566;
    wire N__12565;
    wire N__12558;
    wire N__12557;
    wire N__12556;
    wire N__12549;
    wire N__12548;
    wire N__12547;
    wire N__12540;
    wire N__12539;
    wire N__12538;
    wire N__12531;
    wire N__12530;
    wire N__12529;
    wire N__12522;
    wire N__12521;
    wire N__12520;
    wire N__12513;
    wire N__12512;
    wire N__12511;
    wire N__12504;
    wire N__12503;
    wire N__12502;
    wire N__12495;
    wire N__12494;
    wire N__12493;
    wire N__12486;
    wire N__12485;
    wire N__12484;
    wire N__12477;
    wire N__12476;
    wire N__12475;
    wire N__12468;
    wire N__12467;
    wire N__12466;
    wire N__12459;
    wire N__12458;
    wire N__12457;
    wire N__12450;
    wire N__12449;
    wire N__12448;
    wire N__12441;
    wire N__12440;
    wire N__12439;
    wire N__12432;
    wire N__12431;
    wire N__12430;
    wire N__12423;
    wire N__12422;
    wire N__12421;
    wire N__12414;
    wire N__12413;
    wire N__12412;
    wire N__12405;
    wire N__12404;
    wire N__12403;
    wire N__12396;
    wire N__12395;
    wire N__12394;
    wire N__12387;
    wire N__12386;
    wire N__12385;
    wire N__12378;
    wire N__12377;
    wire N__12376;
    wire N__12369;
    wire N__12368;
    wire N__12367;
    wire N__12360;
    wire N__12359;
    wire N__12358;
    wire N__12351;
    wire N__12350;
    wire N__12349;
    wire N__12342;
    wire N__12341;
    wire N__12340;
    wire N__12333;
    wire N__12332;
    wire N__12331;
    wire N__12324;
    wire N__12323;
    wire N__12322;
    wire N__12315;
    wire N__12314;
    wire N__12313;
    wire N__12306;
    wire N__12305;
    wire N__12304;
    wire N__12297;
    wire N__12296;
    wire N__12295;
    wire N__12288;
    wire N__12287;
    wire N__12286;
    wire N__12269;
    wire N__12266;
    wire N__12263;
    wire N__12260;
    wire N__12257;
    wire N__12254;
    wire N__12251;
    wire N__12248;
    wire N__12247;
    wire N__12244;
    wire N__12243;
    wire N__12242;
    wire N__12241;
    wire N__12240;
    wire N__12237;
    wire N__12234;
    wire N__12231;
    wire N__12230;
    wire N__12229;
    wire N__12228;
    wire N__12227;
    wire N__12226;
    wire N__12225;
    wire N__12224;
    wire N__12221;
    wire N__12218;
    wire N__12215;
    wire N__12214;
    wire N__12209;
    wire N__12206;
    wire N__12203;
    wire N__12200;
    wire N__12199;
    wire N__12196;
    wire N__12193;
    wire N__12190;
    wire N__12187;
    wire N__12186;
    wire N__12185;
    wire N__12184;
    wire N__12183;
    wire N__12182;
    wire N__12181;
    wire N__12178;
    wire N__12171;
    wire N__12168;
    wire N__12165;
    wire N__12164;
    wire N__12163;
    wire N__12160;
    wire N__12157;
    wire N__12154;
    wire N__12153;
    wire N__12152;
    wire N__12151;
    wire N__12150;
    wire N__12149;
    wire N__12148;
    wire N__12141;
    wire N__12134;
    wire N__12127;
    wire N__12124;
    wire N__12123;
    wire N__12122;
    wire N__12121;
    wire N__12120;
    wire N__12119;
    wire N__12118;
    wire N__12115;
    wire N__12112;
    wire N__12107;
    wire N__12104;
    wire N__12099;
    wire N__12092;
    wire N__12085;
    wire N__12080;
    wire N__12077;
    wire N__12070;
    wire N__12063;
    wire N__12056;
    wire N__12051;
    wire N__12026;
    wire N__12023;
    wire N__12020;
    wire N__12017;
    wire N__12014;
    wire N__12013;
    wire N__12010;
    wire N__12007;
    wire N__12006;
    wire N__12003;
    wire N__12000;
    wire N__11997;
    wire N__11996;
    wire N__11991;
    wire N__11988;
    wire N__11985;
    wire N__11984;
    wire N__11979;
    wire N__11976;
    wire N__11973;
    wire N__11970;
    wire N__11967;
    wire N__11960;
    wire N__11957;
    wire N__11954;
    wire N__11951;
    wire N__11948;
    wire N__11945;
    wire N__11942;
    wire N__11939;
    wire N__11938;
    wire N__11937;
    wire N__11936;
    wire N__11933;
    wire N__11930;
    wire N__11927;
    wire N__11924;
    wire N__11921;
    wire N__11918;
    wire N__11913;
    wire N__11908;
    wire N__11905;
    wire N__11902;
    wire N__11899;
    wire N__11894;
    wire N__11893;
    wire N__11890;
    wire N__11887;
    wire N__11886;
    wire N__11885;
    wire N__11880;
    wire N__11877;
    wire N__11874;
    wire N__11867;
    wire N__11864;
    wire N__11861;
    wire N__11858;
    wire N__11855;
    wire N__11852;
    wire N__11849;
    wire N__11846;
    wire N__11845;
    wire N__11842;
    wire N__11841;
    wire N__11838;
    wire N__11835;
    wire N__11832;
    wire N__11829;
    wire N__11828;
    wire N__11825;
    wire N__11822;
    wire N__11819;
    wire N__11816;
    wire N__11811;
    wire N__11806;
    wire N__11803;
    wire N__11798;
    wire N__11795;
    wire N__11792;
    wire N__11789;
    wire N__11786;
    wire N__11783;
    wire N__11782;
    wire N__11781;
    wire N__11780;
    wire N__11779;
    wire N__11778;
    wire N__11777;
    wire N__11776;
    wire N__11775;
    wire N__11772;
    wire N__11769;
    wire N__11766;
    wire N__11761;
    wire N__11756;
    wire N__11753;
    wire N__11752;
    wire N__11751;
    wire N__11750;
    wire N__11749;
    wire N__11748;
    wire N__11747;
    wire N__11746;
    wire N__11743;
    wire N__11740;
    wire N__11737;
    wire N__11728;
    wire N__11723;
    wire N__11720;
    wire N__11717;
    wire N__11714;
    wire N__11711;
    wire N__11710;
    wire N__11707;
    wire N__11706;
    wire N__11705;
    wire N__11702;
    wire N__11701;
    wire N__11700;
    wire N__11695;
    wire N__11682;
    wire N__11679;
    wire N__11676;
    wire N__11671;
    wire N__11668;
    wire N__11665;
    wire N__11662;
    wire N__11657;
    wire N__11654;
    wire N__11651;
    wire N__11642;
    wire N__11637;
    wire N__11634;
    wire N__11631;
    wire N__11628;
    wire N__11623;
    wire N__11620;
    wire N__11615;
    wire N__11612;
    wire N__11609;
    wire N__11606;
    wire N__11603;
    wire N__11602;
    wire N__11601;
    wire N__11600;
    wire N__11599;
    wire N__11598;
    wire N__11597;
    wire N__11596;
    wire N__11579;
    wire N__11576;
    wire N__11573;
    wire N__11572;
    wire N__11571;
    wire N__11570;
    wire N__11569;
    wire N__11568;
    wire N__11567;
    wire N__11566;
    wire N__11565;
    wire N__11564;
    wire N__11563;
    wire N__11562;
    wire N__11561;
    wire N__11560;
    wire N__11559;
    wire N__11528;
    wire N__11525;
    wire N__11522;
    wire N__11521;
    wire N__11518;
    wire N__11515;
    wire N__11512;
    wire N__11509;
    wire N__11504;
    wire N__11501;
    wire N__11498;
    wire N__11495;
    wire N__11492;
    wire N__11489;
    wire N__11486;
    wire N__11483;
    wire N__11480;
    wire N__11477;
    wire N__11474;
    wire N__11471;
    wire N__11470;
    wire N__11469;
    wire N__11468;
    wire N__11467;
    wire N__11466;
    wire N__11465;
    wire N__11464;
    wire N__11463;
    wire N__11462;
    wire N__11461;
    wire N__11460;
    wire N__11459;
    wire N__11458;
    wire N__11457;
    wire N__11456;
    wire N__11455;
    wire N__11454;
    wire N__11453;
    wire N__11452;
    wire N__11451;
    wire N__11450;
    wire N__11449;
    wire N__11448;
    wire N__11447;
    wire N__11446;
    wire N__11445;
    wire N__11444;
    wire N__11443;
    wire N__11442;
    wire N__11441;
    wire N__11440;
    wire N__11439;
    wire N__11438;
    wire N__11437;
    wire N__11436;
    wire N__11435;
    wire N__11432;
    wire N__11431;
    wire N__11430;
    wire N__11429;
    wire N__11428;
    wire N__11427;
    wire N__11426;
    wire N__11425;
    wire N__11424;
    wire N__11423;
    wire N__11330;
    wire N__11327;
    wire N__11326;
    wire N__11325;
    wire N__11324;
    wire N__11323;
    wire N__11320;
    wire N__11317;
    wire N__11314;
    wire N__11311;
    wire N__11308;
    wire N__11307;
    wire N__11306;
    wire N__11303;
    wire N__11302;
    wire N__11301;
    wire N__11300;
    wire N__11299;
    wire N__11298;
    wire N__11297;
    wire N__11296;
    wire N__11295;
    wire N__11294;
    wire N__11293;
    wire N__11292;
    wire N__11291;
    wire N__11290;
    wire N__11289;
    wire N__11288;
    wire N__11287;
    wire N__11286;
    wire N__11285;
    wire N__11284;
    wire N__11283;
    wire N__11282;
    wire N__11281;
    wire N__11280;
    wire N__11279;
    wire N__11278;
    wire N__11277;
    wire N__11276;
    wire N__11275;
    wire N__11272;
    wire N__11269;
    wire N__11268;
    wire N__11267;
    wire N__11266;
    wire N__11265;
    wire N__11264;
    wire N__11263;
    wire N__11262;
    wire N__11261;
    wire N__11260;
    wire N__11259;
    wire N__11258;
    wire N__11257;
    wire N__11256;
    wire N__11255;
    wire N__11254;
    wire N__11251;
    wire N__11250;
    wire N__11247;
    wire N__11246;
    wire N__11245;
    wire N__11244;
    wire N__11135;
    wire N__11132;
    wire N__11129;
    wire N__11126;
    wire N__11123;
    wire N__11122;
    wire N__11119;
    wire N__11116;
    wire N__11113;
    wire N__11110;
    wire N__11109;
    wire N__11108;
    wire N__11105;
    wire N__11102;
    wire N__11099;
    wire N__11096;
    wire N__11087;
    wire N__11084;
    wire N__11081;
    wire N__11080;
    wire N__11077;
    wire N__11076;
    wire N__11073;
    wire N__11072;
    wire N__11071;
    wire N__11070;
    wire N__11067;
    wire N__11066;
    wire N__11065;
    wire N__11064;
    wire N__11063;
    wire N__11062;
    wire N__11061;
    wire N__11060;
    wire N__11057;
    wire N__11052;
    wire N__11047;
    wire N__11046;
    wire N__11045;
    wire N__11044;
    wire N__11043;
    wire N__11040;
    wire N__11031;
    wire N__11030;
    wire N__11029;
    wire N__11026;
    wire N__11023;
    wire N__11022;
    wire N__11019;
    wire N__11016;
    wire N__11013;
    wire N__11010;
    wire N__11005;
    wire N__11004;
    wire N__11001;
    wire N__11000;
    wire N__10999;
    wire N__10998;
    wire N__10995;
    wire N__10994;
    wire N__10993;
    wire N__10992;
    wire N__10987;
    wire N__10984;
    wire N__10981;
    wire N__10976;
    wire N__10973;
    wire N__10970;
    wire N__10961;
    wire N__10958;
    wire N__10955;
    wire N__10948;
    wire N__10945;
    wire N__10940;
    wire N__10939;
    wire N__10938;
    wire N__10937;
    wire N__10934;
    wire N__10929;
    wire N__10916;
    wire N__10915;
    wire N__10908;
    wire N__10905;
    wire N__10898;
    wire N__10895;
    wire N__10890;
    wire N__10887;
    wire N__10880;
    wire N__10871;
    wire N__10868;
    wire N__10865;
    wire N__10862;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10852;
    wire N__10849;
    wire N__10846;
    wire N__10845;
    wire N__10840;
    wire N__10837;
    wire N__10836;
    wire N__10831;
    wire N__10830;
    wire N__10827;
    wire N__10824;
    wire N__10819;
    wire N__10816;
    wire N__10813;
    wire N__10810;
    wire N__10807;
    wire N__10802;
    wire N__10801;
    wire N__10798;
    wire N__10795;
    wire N__10794;
    wire N__10793;
    wire N__10792;
    wire N__10789;
    wire N__10786;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10772;
    wire N__10769;
    wire N__10766;
    wire N__10763;
    wire N__10758;
    wire N__10755;
    wire N__10748;
    wire N__10745;
    wire N__10742;
    wire N__10739;
    wire N__10736;
    wire N__10735;
    wire N__10732;
    wire N__10729;
    wire N__10724;
    wire N__10723;
    wire N__10720;
    wire N__10717;
    wire N__10712;
    wire N__10709;
    wire N__10708;
    wire N__10707;
    wire N__10704;
    wire N__10701;
    wire N__10698;
    wire N__10693;
    wire N__10690;
    wire N__10685;
    wire N__10684;
    wire N__10683;
    wire N__10680;
    wire N__10675;
    wire N__10670;
    wire N__10667;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10655;
    wire N__10652;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10642;
    wire N__10639;
    wire N__10636;
    wire N__10631;
    wire N__10630;
    wire N__10629;
    wire N__10626;
    wire N__10623;
    wire N__10620;
    wire N__10617;
    wire N__10612;
    wire N__10607;
    wire N__10604;
    wire N__10601;
    wire N__10598;
    wire N__10595;
    wire N__10592;
    wire N__10589;
    wire N__10586;
    wire N__10583;
    wire N__10580;
    wire N__10579;
    wire N__10576;
    wire N__10573;
    wire N__10572;
    wire N__10571;
    wire N__10566;
    wire N__10563;
    wire N__10560;
    wire N__10557;
    wire N__10552;
    wire N__10549;
    wire N__10544;
    wire N__10541;
    wire N__10538;
    wire N__10535;
    wire N__10532;
    wire N__10529;
    wire N__10528;
    wire N__10527;
    wire N__10524;
    wire N__10521;
    wire N__10518;
    wire N__10517;
    wire N__10510;
    wire N__10507;
    wire N__10504;
    wire N__10501;
    wire N__10498;
    wire N__10495;
    wire N__10492;
    wire N__10489;
    wire N__10486;
    wire N__10483;
    wire N__10478;
    wire N__10475;
    wire N__10472;
    wire N__10469;
    wire N__10466;
    wire N__10463;
    wire N__10460;
    wire N__10457;
    wire N__10454;
    wire N__10451;
    wire N__10450;
    wire N__10447;
    wire N__10444;
    wire N__10441;
    wire N__10438;
    wire N__10435;
    wire N__10432;
    wire N__10429;
    wire N__10426;
    wire N__10423;
    wire N__10418;
    wire N__10417;
    wire N__10414;
    wire N__10413;
    wire N__10410;
    wire N__10409;
    wire N__10406;
    wire N__10403;
    wire N__10400;
    wire N__10397;
    wire N__10390;
    wire N__10387;
    wire N__10384;
    wire N__10381;
    wire N__10378;
    wire N__10375;
    wire N__10372;
    wire N__10369;
    wire N__10364;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10351;
    wire N__10350;
    wire N__10347;
    wire N__10344;
    wire N__10341;
    wire N__10338;
    wire N__10337;
    wire N__10332;
    wire N__10331;
    wire N__10330;
    wire N__10327;
    wire N__10324;
    wire N__10321;
    wire N__10318;
    wire N__10315;
    wire N__10312;
    wire N__10309;
    wire N__10298;
    wire N__10297;
    wire N__10292;
    wire N__10289;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10274;
    wire N__10271;
    wire N__10268;
    wire N__10265;
    wire N__10264;
    wire N__10263;
    wire N__10262;
    wire N__10259;
    wire N__10256;
    wire N__10253;
    wire N__10252;
    wire N__10249;
    wire N__10246;
    wire N__10243;
    wire N__10236;
    wire N__10235;
    wire N__10232;
    wire N__10227;
    wire N__10224;
    wire N__10217;
    wire N__10214;
    wire N__10211;
    wire N__10208;
    wire N__10205;
    wire N__10202;
    wire N__10199;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10187;
    wire N__10186;
    wire N__10183;
    wire N__10180;
    wire N__10177;
    wire N__10174;
    wire N__10169;
    wire N__10168;
    wire N__10167;
    wire N__10164;
    wire N__10161;
    wire N__10156;
    wire N__10155;
    wire N__10152;
    wire N__10149;
    wire N__10146;
    wire N__10143;
    wire N__10140;
    wire N__10137;
    wire N__10134;
    wire N__10129;
    wire N__10124;
    wire N__10121;
    wire N__10118;
    wire N__10115;
    wire N__10114;
    wire N__10111;
    wire N__10108;
    wire N__10105;
    wire N__10102;
    wire N__10097;
    wire N__10096;
    wire N__10095;
    wire N__10094;
    wire N__10091;
    wire N__10090;
    wire N__10083;
    wire N__10078;
    wire N__10077;
    wire N__10074;
    wire N__10071;
    wire N__10068;
    wire N__10065;
    wire N__10062;
    wire N__10059;
    wire N__10056;
    wire N__10051;
    wire N__10048;
    wire N__10045;
    wire N__10040;
    wire N__10037;
    wire N__10036;
    wire N__10035;
    wire N__10034;
    wire N__10027;
    wire N__10024;
    wire N__10021;
    wire N__10018;
    wire N__10015;
    wire N__10012;
    wire N__10007;
    wire N__10004;
    wire N__10001;
    wire N__10000;
    wire N__9999;
    wire N__9996;
    wire N__9993;
    wire N__9990;
    wire N__9989;
    wire N__9988;
    wire N__9987;
    wire N__9984;
    wire N__9979;
    wire N__9974;
    wire N__9971;
    wire N__9964;
    wire N__9961;
    wire N__9958;
    wire N__9955;
    wire N__9952;
    wire N__9949;
    wire N__9946;
    wire N__9943;
    wire N__9938;
    wire N__9937;
    wire N__9936;
    wire N__9933;
    wire N__9928;
    wire N__9923;
    wire N__9920;
    wire N__9917;
    wire N__9914;
    wire N__9911;
    wire N__9910;
    wire N__9907;
    wire N__9904;
    wire N__9899;
    wire N__9896;
    wire N__9893;
    wire N__9892;
    wire N__9891;
    wire N__9888;
    wire N__9885;
    wire N__9884;
    wire N__9881;
    wire N__9880;
    wire N__9877;
    wire N__9874;
    wire N__9873;
    wire N__9870;
    wire N__9867;
    wire N__9864;
    wire N__9859;
    wire N__9856;
    wire N__9855;
    wire N__9854;
    wire N__9849;
    wire N__9846;
    wire N__9843;
    wire N__9840;
    wire N__9837;
    wire N__9834;
    wire N__9821;
    wire N__9818;
    wire N__9815;
    wire N__9812;
    wire N__9809;
    wire N__9806;
    wire N__9803;
    wire N__9800;
    wire N__9797;
    wire N__9794;
    wire N__9793;
    wire N__9792;
    wire N__9789;
    wire N__9786;
    wire N__9783;
    wire N__9782;
    wire N__9775;
    wire N__9772;
    wire N__9767;
    wire N__9764;
    wire N__9761;
    wire N__9758;
    wire N__9755;
    wire N__9752;
    wire N__9749;
    wire N__9746;
    wire N__9743;
    wire N__9742;
    wire N__9741;
    wire N__9740;
    wire N__9737;
    wire N__9734;
    wire N__9729;
    wire N__9722;
    wire N__9719;
    wire N__9716;
    wire N__9713;
    wire N__9710;
    wire N__9707;
    wire N__9704;
    wire N__9701;
    wire N__9698;
    wire N__9695;
    wire N__9692;
    wire N__9689;
    wire N__9686;
    wire N__9683;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9671;
    wire N__9668;
    wire N__9667;
    wire N__9666;
    wire N__9663;
    wire N__9660;
    wire N__9657;
    wire N__9654;
    wire N__9651;
    wire N__9648;
    wire N__9647;
    wire N__9646;
    wire N__9645;
    wire N__9642;
    wire N__9637;
    wire N__9634;
    wire N__9631;
    wire N__9628;
    wire N__9617;
    wire N__9614;
    wire N__9611;
    wire N__9608;
    wire N__9605;
    wire N__9602;
    wire N__9599;
    wire N__9596;
    wire N__9593;
    wire N__9590;
    wire N__9587;
    wire N__9584;
    wire N__9581;
    wire N__9578;
    wire N__9575;
    wire N__9572;
    wire N__9569;
    wire N__9566;
    wire N__9563;
    wire N__9560;
    wire N__9557;
    wire N__9554;
    wire N__9551;
    wire N__9548;
    wire N__9547;
    wire N__9544;
    wire N__9541;
    wire N__9538;
    wire N__9535;
    wire N__9532;
    wire N__9529;
    wire N__9524;
    wire N__9521;
    wire N__9518;
    wire N__9515;
    wire N__9512;
    wire N__9509;
    wire N__9506;
    wire N__9503;
    wire N__9500;
    wire N__9497;
    wire N__9494;
    wire N__9491;
    wire N__9488;
    wire N__9485;
    wire N__9482;
    wire N__9479;
    wire N__9476;
    wire N__9473;
    wire N__9470;
    wire N__9467;
    wire N__9464;
    wire N__9461;
    wire N__9458;
    wire N__9457;
    wire N__9454;
    wire N__9453;
    wire N__9452;
    wire N__9451;
    wire N__9450;
    wire N__9447;
    wire N__9444;
    wire N__9441;
    wire N__9440;
    wire N__9439;
    wire N__9436;
    wire N__9435;
    wire N__9432;
    wire N__9431;
    wire N__9430;
    wire N__9427;
    wire N__9426;
    wire N__9425;
    wire N__9422;
    wire N__9419;
    wire N__9416;
    wire N__9415;
    wire N__9414;
    wire N__9411;
    wire N__9408;
    wire N__9405;
    wire N__9402;
    wire N__9399;
    wire N__9396;
    wire N__9389;
    wire N__9386;
    wire N__9381;
    wire N__9378;
    wire N__9373;
    wire N__9370;
    wire N__9367;
    wire N__9362;
    wire N__9341;
    wire N__9338;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9326;
    wire N__9323;
    wire N__9320;
    wire N__9317;
    wire N__9314;
    wire N__9311;
    wire N__9308;
    wire N__9305;
    wire N__9302;
    wire N__9299;
    wire N__9296;
    wire N__9293;
    wire N__9290;
    wire N__9287;
    wire N__9284;
    wire N__9281;
    wire N__9278;
    wire N__9275;
    wire N__9272;
    wire N__9269;
    wire N__9266;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9242;
    wire N__9241;
    wire N__9238;
    wire N__9235;
    wire N__9234;
    wire N__9233;
    wire N__9232;
    wire N__9229;
    wire N__9228;
    wire N__9225;
    wire N__9222;
    wire N__9221;
    wire N__9220;
    wire N__9217;
    wire N__9214;
    wire N__9211;
    wire N__9208;
    wire N__9205;
    wire N__9202;
    wire N__9199;
    wire N__9196;
    wire N__9187;
    wire N__9176;
    wire N__9173;
    wire N__9170;
    wire N__9167;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9145;
    wire N__9142;
    wire N__9139;
    wire N__9136;
    wire N__9131;
    wire N__9130;
    wire N__9127;
    wire N__9126;
    wire N__9125;
    wire N__9124;
    wire N__9123;
    wire N__9122;
    wire N__9121;
    wire N__9120;
    wire N__9119;
    wire N__9118;
    wire N__9115;
    wire N__9112;
    wire N__9107;
    wire N__9104;
    wire N__9103;
    wire N__9102;
    wire N__9099;
    wire N__9096;
    wire N__9093;
    wire N__9090;
    wire N__9089;
    wire N__9088;
    wire N__9087;
    wire N__9086;
    wire N__9081;
    wire N__9078;
    wire N__9071;
    wire N__9068;
    wire N__9065;
    wire N__9062;
    wire N__9059;
    wire N__9056;
    wire N__9049;
    wire N__9044;
    wire N__9037;
    wire N__9020;
    wire N__9017;
    wire N__9014;
    wire N__9011;
    wire N__9008;
    wire N__9005;
    wire N__9002;
    wire N__8999;
    wire N__8996;
    wire N__8993;
    wire N__8992;
    wire N__8989;
    wire N__8986;
    wire N__8981;
    wire N__8980;
    wire N__8979;
    wire N__8978;
    wire N__8977;
    wire N__8976;
    wire N__8975;
    wire N__8974;
    wire N__8967;
    wire N__8962;
    wire N__8955;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8935;
    wire N__8932;
    wire N__8929;
    wire N__8924;
    wire N__8923;
    wire N__8922;
    wire N__8921;
    wire N__8920;
    wire N__8919;
    wire N__8916;
    wire N__8915;
    wire N__8914;
    wire N__8913;
    wire N__8910;
    wire N__8907;
    wire N__8900;
    wire N__8899;
    wire N__8896;
    wire N__8889;
    wire N__8888;
    wire N__8887;
    wire N__8886;
    wire N__8885;
    wire N__8884;
    wire N__8883;
    wire N__8882;
    wire N__8875;
    wire N__8874;
    wire N__8873;
    wire N__8872;
    wire N__8871;
    wire N__8868;
    wire N__8867;
    wire N__8866;
    wire N__8861;
    wire N__8854;
    wire N__8847;
    wire N__8846;
    wire N__8845;
    wire N__8842;
    wire N__8841;
    wire N__8838;
    wire N__8833;
    wire N__8830;
    wire N__8821;
    wire N__8816;
    wire N__8813;
    wire N__8808;
    wire N__8803;
    wire N__8786;
    wire N__8785;
    wire N__8784;
    wire N__8781;
    wire N__8780;
    wire N__8779;
    wire N__8776;
    wire N__8773;
    wire N__8772;
    wire N__8771;
    wire N__8768;
    wire N__8763;
    wire N__8760;
    wire N__8757;
    wire N__8754;
    wire N__8751;
    wire N__8738;
    wire N__8735;
    wire N__8732;
    wire N__8729;
    wire N__8726;
    wire N__8723;
    wire N__8720;
    wire N__8719;
    wire N__8716;
    wire N__8713;
    wire N__8710;
    wire N__8707;
    wire N__8702;
    wire N__8699;
    wire N__8696;
    wire N__8693;
    wire N__8690;
    wire N__8687;
    wire N__8686;
    wire N__8685;
    wire N__8682;
    wire N__8681;
    wire N__8680;
    wire N__8677;
    wire N__8676;
    wire N__8673;
    wire N__8672;
    wire N__8671;
    wire N__8670;
    wire N__8669;
    wire N__8668;
    wire N__8667;
    wire N__8666;
    wire N__8665;
    wire N__8664;
    wire N__8659;
    wire N__8658;
    wire N__8655;
    wire N__8654;
    wire N__8653;
    wire N__8650;
    wire N__8647;
    wire N__8642;
    wire N__8641;
    wire N__8640;
    wire N__8639;
    wire N__8636;
    wire N__8629;
    wire N__8628;
    wire N__8627;
    wire N__8626;
    wire N__8625;
    wire N__8618;
    wire N__8615;
    wire N__8612;
    wire N__8603;
    wire N__8596;
    wire N__8595;
    wire N__8594;
    wire N__8593;
    wire N__8590;
    wire N__8589;
    wire N__8586;
    wire N__8585;
    wire N__8582;
    wire N__8577;
    wire N__8570;
    wire N__8567;
    wire N__8564;
    wire N__8555;
    wire N__8548;
    wire N__8545;
    wire N__8542;
    wire N__8539;
    wire N__8536;
    wire N__8513;
    wire N__8510;
    wire N__8507;
    wire N__8504;
    wire N__8501;
    wire N__8498;
    wire N__8497;
    wire N__8494;
    wire N__8491;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8462;
    wire N__8461;
    wire N__8458;
    wire N__8455;
    wire N__8452;
    wire N__8449;
    wire N__8446;
    wire N__8443;
    wire N__8440;
    wire N__8437;
    wire N__8432;
    wire N__8429;
    wire N__8426;
    wire N__8425;
    wire N__8422;
    wire N__8419;
    wire N__8416;
    wire N__8413;
    wire N__8410;
    wire N__8405;
    wire N__8402;
    wire N__8399;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8384;
    wire N__8381;
    wire N__8378;
    wire N__8375;
    wire N__8372;
    wire N__8371;
    wire N__8370;
    wire N__8369;
    wire N__8368;
    wire N__8365;
    wire N__8362;
    wire N__8361;
    wire N__8360;
    wire N__8357;
    wire N__8356;
    wire N__8355;
    wire N__8354;
    wire N__8351;
    wire N__8348;
    wire N__8345;
    wire N__8338;
    wire N__8335;
    wire N__8330;
    wire N__8325;
    wire N__8322;
    wire N__8317;
    wire N__8306;
    wire N__8305;
    wire N__8304;
    wire N__8303;
    wire N__8300;
    wire N__8299;
    wire N__8296;
    wire N__8295;
    wire N__8294;
    wire N__8291;
    wire N__8286;
    wire N__8283;
    wire N__8280;
    wire N__8275;
    wire N__8272;
    wire N__8269;
    wire N__8266;
    wire N__8263;
    wire N__8252;
    wire N__8249;
    wire N__8246;
    wire N__8243;
    wire N__8240;
    wire N__8237;
    wire N__8234;
    wire N__8231;
    wire N__8228;
    wire N__8225;
    wire N__8222;
    wire N__8219;
    wire N__8216;
    wire N__8213;
    wire N__8210;
    wire N__8209;
    wire N__8206;
    wire N__8203;
    wire N__8202;
    wire N__8199;
    wire N__8196;
    wire N__8193;
    wire N__8190;
    wire N__8187;
    wire N__8184;
    wire N__8177;
    wire N__8174;
    wire N__8171;
    wire N__8168;
    wire N__8167;
    wire N__8164;
    wire N__8161;
    wire N__8156;
    wire N__8155;
    wire N__8154;
    wire N__8153;
    wire N__8152;
    wire N__8149;
    wire N__8148;
    wire N__8145;
    wire N__8142;
    wire N__8135;
    wire N__8132;
    wire N__8125;
    wire N__8122;
    wire N__8119;
    wire N__8114;
    wire N__8113;
    wire N__8112;
    wire N__8111;
    wire N__8110;
    wire N__8109;
    wire N__8108;
    wire N__8101;
    wire N__8100;
    wire N__8099;
    wire N__8098;
    wire N__8097;
    wire N__8096;
    wire N__8095;
    wire N__8094;
    wire N__8087;
    wire N__8086;
    wire N__8085;
    wire N__8084;
    wire N__8081;
    wire N__8080;
    wire N__8077;
    wire N__8074;
    wire N__8065;
    wire N__8062;
    wire N__8061;
    wire N__8058;
    wire N__8057;
    wire N__8056;
    wire N__8053;
    wire N__8048;
    wire N__8047;
    wire N__8040;
    wire N__8039;
    wire N__8038;
    wire N__8037;
    wire N__8036;
    wire N__8031;
    wire N__8028;
    wire N__8025;
    wire N__8022;
    wire N__8019;
    wire N__8014;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__8000;
    wire N__7995;
    wire N__7992;
    wire N__7989;
    wire N__7984;
    wire N__7981;
    wire N__7976;
    wire N__7971;
    wire N__7964;
    wire N__7963;
    wire N__7960;
    wire N__7953;
    wire N__7946;
    wire N__7943;
    wire N__7936;
    wire N__7933;
    wire N__7930;
    wire N__7927;
    wire N__7922;
    wire N__7919;
    wire N__7916;
    wire N__7913;
    wire N__7910;
    wire N__7907;
    wire N__7904;
    wire N__7901;
    wire N__7898;
    wire N__7895;
    wire N__7892;
    wire N__7889;
    wire N__7886;
    wire N__7883;
    wire N__7880;
    wire N__7877;
    wire N__7874;
    wire N__7871;
    wire N__7868;
    wire N__7865;
    wire N__7862;
    wire N__7861;
    wire N__7858;
    wire N__7855;
    wire N__7850;
    wire N__7849;
    wire N__7844;
    wire N__7841;
    wire N__7840;
    wire N__7837;
    wire N__7834;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7816;
    wire N__7813;
    wire N__7810;
    wire N__7809;
    wire N__7806;
    wire N__7803;
    wire N__7802;
    wire N__7801;
    wire N__7800;
    wire N__7799;
    wire N__7796;
    wire N__7791;
    wire N__7786;
    wire N__7781;
    wire N__7772;
    wire N__7771;
    wire N__7770;
    wire N__7767;
    wire N__7766;
    wire N__7763;
    wire N__7760;
    wire N__7757;
    wire N__7756;
    wire N__7753;
    wire N__7752;
    wire N__7751;
    wire N__7750;
    wire N__7749;
    wire N__7748;
    wire N__7747;
    wire N__7746;
    wire N__7741;
    wire N__7738;
    wire N__7727;
    wire N__7726;
    wire N__7725;
    wire N__7724;
    wire N__7721;
    wire N__7718;
    wire N__7713;
    wire N__7710;
    wire N__7705;
    wire N__7698;
    wire N__7685;
    wire N__7682;
    wire N__7681;
    wire N__7680;
    wire N__7679;
    wire N__7676;
    wire N__7673;
    wire N__7670;
    wire N__7667;
    wire N__7666;
    wire N__7663;
    wire N__7660;
    wire N__7655;
    wire N__7652;
    wire N__7643;
    wire N__7640;
    wire N__7637;
    wire N__7634;
    wire N__7631;
    wire N__7628;
    wire N__7625;
    wire N__7622;
    wire N__7619;
    wire N__7616;
    wire N__7613;
    wire N__7610;
    wire N__7607;
    wire N__7604;
    wire N__7601;
    wire N__7598;
    wire N__7597;
    wire N__7594;
    wire N__7591;
    wire N__7586;
    wire N__7583;
    wire N__7582;
    wire N__7581;
    wire N__7580;
    wire N__7579;
    wire N__7578;
    wire N__7575;
    wire N__7568;
    wire N__7565;
    wire N__7564;
    wire N__7561;
    wire N__7558;
    wire N__7555;
    wire N__7552;
    wire N__7549;
    wire N__7546;
    wire N__7543;
    wire N__7538;
    wire N__7529;
    wire N__7528;
    wire N__7525;
    wire N__7524;
    wire N__7521;
    wire N__7518;
    wire N__7515;
    wire N__7512;
    wire N__7505;
    wire N__7504;
    wire N__7503;
    wire N__7500;
    wire N__7499;
    wire N__7494;
    wire N__7491;
    wire N__7488;
    wire N__7481;
    wire N__7478;
    wire N__7475;
    wire N__7472;
    wire N__7469;
    wire N__7466;
    wire N__7463;
    wire N__7460;
    wire N__7459;
    wire N__7456;
    wire N__7453;
    wire N__7448;
    wire N__7445;
    wire N__7442;
    wire N__7439;
    wire N__7436;
    wire N__7433;
    wire N__7430;
    wire N__7429;
    wire N__7426;
    wire N__7423;
    wire N__7420;
    wire N__7415;
    wire N__7412;
    wire N__7409;
    wire N__7406;
    wire N__7403;
    wire N__7400;
    wire N__7397;
    wire N__7394;
    wire N__7393;
    wire N__7390;
    wire N__7387;
    wire N__7384;
    wire N__7379;
    wire N__7376;
    wire N__7373;
    wire N__7370;
    wire N__7367;
    wire N__7364;
    wire N__7361;
    wire N__7360;
    wire N__7357;
    wire N__7354;
    wire N__7351;
    wire N__7346;
    wire N__7343;
    wire N__7340;
    wire N__7337;
    wire N__7336;
    wire N__7335;
    wire N__7332;
    wire N__7329;
    wire N__7326;
    wire N__7325;
    wire N__7320;
    wire N__7317;
    wire N__7314;
    wire N__7311;
    wire N__7304;
    wire N__7303;
    wire N__7300;
    wire N__7299;
    wire N__7298;
    wire N__7297;
    wire N__7294;
    wire N__7291;
    wire N__7286;
    wire N__7283;
    wire N__7282;
    wire N__7281;
    wire N__7280;
    wire N__7279;
    wire N__7276;
    wire N__7273;
    wire N__7268;
    wire N__7265;
    wire N__7262;
    wire N__7257;
    wire N__7254;
    wire N__7249;
    wire N__7238;
    wire N__7235;
    wire N__7232;
    wire N__7229;
    wire N__7226;
    wire N__7223;
    wire N__7220;
    wire N__7217;
    wire N__7216;
    wire N__7213;
    wire N__7210;
    wire N__7205;
    wire N__7202;
    wire N__7199;
    wire N__7196;
    wire N__7193;
    wire N__7192;
    wire N__7189;
    wire N__7186;
    wire N__7183;
    wire N__7180;
    wire N__7177;
    wire N__7174;
    wire N__7171;
    wire N__7168;
    wire N__7163;
    wire N__7160;
    wire N__7157;
    wire N__7154;
    wire N__7151;
    wire N__7148;
    wire N__7145;
    wire N__7142;
    wire N__7139;
    wire N__7138;
    wire N__7137;
    wire N__7136;
    wire N__7133;
    wire N__7130;
    wire N__7125;
    wire N__7118;
    wire N__7115;
    wire N__7112;
    wire N__7109;
    wire N__7106;
    wire N__7103;
    wire N__7100;
    wire N__7097;
    wire N__7096;
    wire N__7095;
    wire N__7094;
    wire N__7093;
    wire N__7090;
    wire N__7087;
    wire N__7084;
    wire N__7079;
    wire N__7070;
    wire N__7069;
    wire N__7068;
    wire N__7067;
    wire N__7064;
    wire N__7061;
    wire N__7056;
    wire N__7051;
    wire N__7046;
    wire N__7043;
    wire N__7042;
    wire N__7039;
    wire N__7036;
    wire N__7033;
    wire N__7028;
    wire N__7025;
    wire N__7024;
    wire N__7023;
    wire N__7022;
    wire N__7019;
    wire N__7018;
    wire N__7017;
    wire N__7010;
    wire N__7007;
    wire N__7002;
    wire N__6995;
    wire N__6992;
    wire N__6989;
    wire N__6986;
    wire N__6983;
    wire N__6980;
    wire N__6977;
    wire N__6976;
    wire N__6975;
    wire N__6972;
    wire N__6969;
    wire N__6966;
    wire N__6959;
    wire N__6956;
    wire N__6953;
    wire N__6950;
    wire N__6947;
    wire N__6944;
    wire N__6941;
    wire N__6938;
    wire N__6935;
    wire N__6932;
    wire N__6929;
    wire N__6926;
    wire N__6923;
    wire N__6920;
    wire N__6917;
    wire N__6914;
    wire N__6911;
    wire N__6908;
    wire N__6905;
    wire N__6902;
    wire N__6899;
    wire N__6896;
    wire N__6893;
    wire N__6890;
    wire N__6887;
    wire N__6884;
    wire N__6881;
    wire N__6878;
    wire N__6875;
    wire N__6872;
    wire N__6869;
    wire N__6868;
    wire N__6867;
    wire N__6864;
    wire N__6861;
    wire N__6858;
    wire N__6855;
    wire N__6852;
    wire N__6849;
    wire N__6842;
    wire N__6839;
    wire N__6836;
    wire N__6833;
    wire N__6832;
    wire N__6831;
    wire N__6828;
    wire N__6825;
    wire N__6822;
    wire N__6819;
    wire N__6816;
    wire N__6813;
    wire N__6810;
    wire N__6807;
    wire N__6804;
    wire N__6801;
    wire N__6798;
    wire N__6795;
    wire N__6792;
    wire N__6789;
    wire N__6786;
    wire N__6781;
    wire N__6776;
    wire N__6773;
    wire N__6770;
    wire N__6767;
    wire N__6764;
    wire N__6761;
    wire N__6758;
    wire N__6755;
    wire N__6752;
    wire N__6749;
    wire N__6746;
    wire N__6743;
    wire N__6740;
    wire N__6737;
    wire N__6734;
    wire N__6731;
    wire N__6728;
    wire N__6725;
    wire N__6722;
    wire N__6719;
    wire N__6716;
    wire N__6713;
    wire N__6710;
    wire N__6707;
    wire N__6704;
    wire N__6701;
    wire N__6698;
    wire N__6695;
    wire N__6692;
    wire N__6689;
    wire N__6686;
    wire N__6683;
    wire N__6680;
    wire N__6677;
    wire N__6674;
    wire N__6671;
    wire N__6668;
    wire N__6665;
    wire N__6662;
    wire N__6659;
    wire N__6656;
    wire N__6653;
    wire N__6650;
    wire N__6647;
    wire N__6644;
    wire N__6641;
    wire N__6638;
    wire N__6635;
    wire N__6632;
    wire N__6629;
    wire N__6626;
    wire N__6623;
    wire N__6622;
    wire N__6619;
    wire N__6616;
    wire N__6611;
    wire N__6610;
    wire N__6607;
    wire N__6604;
    wire N__6599;
    wire N__6598;
    wire N__6595;
    wire N__6592;
    wire N__6587;
    wire N__6586;
    wire N__6583;
    wire N__6580;
    wire N__6577;
    wire N__6572;
    wire N__6571;
    wire N__6568;
    wire N__6565;
    wire N__6560;
    wire N__6557;
    wire N__6556;
    wire N__6555;
    wire N__6554;
    wire N__6551;
    wire N__6546;
    wire N__6545;
    wire N__6544;
    wire N__6541;
    wire N__6538;
    wire N__6535;
    wire N__6530;
    wire N__6527;
    wire N__6518;
    wire N__6517;
    wire N__6514;
    wire N__6511;
    wire N__6508;
    wire N__6503;
    wire N__6500;
    wire N__6497;
    wire N__6494;
    wire N__6491;
    wire N__6488;
    wire N__6487;
    wire N__6486;
    wire N__6485;
    wire N__6484;
    wire N__6483;
    wire N__6482;
    wire N__6481;
    wire N__6478;
    wire N__6471;
    wire N__6464;
    wire N__6461;
    wire N__6452;
    wire N__6449;
    wire N__6446;
    wire N__6443;
    wire N__6442;
    wire N__6441;
    wire N__6440;
    wire N__6439;
    wire N__6438;
    wire N__6437;
    wire N__6434;
    wire N__6431;
    wire N__6428;
    wire N__6425;
    wire N__6418;
    wire N__6415;
    wire N__6410;
    wire N__6407;
    wire N__6406;
    wire N__6399;
    wire N__6396;
    wire N__6393;
    wire N__6386;
    wire N__6385;
    wire N__6380;
    wire N__6377;
    wire N__6374;
    wire N__6371;
    wire N__6368;
    wire N__6367;
    wire N__6364;
    wire N__6361;
    wire N__6356;
    wire N__6353;
    wire N__6350;
    wire N__6347;
    wire N__6344;
    wire N__6341;
    wire N__6338;
    wire N__6335;
    wire N__6332;
    wire N__6329;
    wire N__6326;
    wire N__6323;
    wire N__6320;
    wire N__6317;
    wire N__6314;
    wire N__6313;
    wire N__6310;
    wire N__6307;
    wire N__6304;
    wire N__6299;
    wire N__6296;
    wire N__6293;
    wire N__6290;
    wire N__6287;
    wire N__6284;
    wire N__6281;
    wire N__6278;
    wire N__6277;
    wire N__6274;
    wire N__6271;
    wire N__6268;
    wire N__6263;
    wire N__6262;
    wire N__6259;
    wire N__6256;
    wire N__6251;
    wire N__6248;
    wire N__6247;
    wire N__6244;
    wire N__6241;
    wire N__6238;
    wire N__6233;
    wire N__6232;
    wire N__6229;
    wire N__6226;
    wire N__6223;
    wire N__6218;
    wire N__6215;
    wire N__6212;
    wire N__6209;
    wire N__6206;
    wire N__6203;
    wire N__6202;
    wire N__6201;
    wire N__6198;
    wire N__6195;
    wire N__6192;
    wire N__6185;
    wire N__6182;
    wire N__6179;
    wire N__6176;
    wire N__6173;
    wire N__6170;
    wire N__6167;
    wire N__6164;
    wire N__6161;
    wire N__6158;
    wire N__6155;
    wire N__6152;
    wire N__6149;
    wire N__6146;
    wire N__6143;
    wire N__6140;
    wire N__6137;
    wire N__6134;
    wire N__6131;
    wire N__6128;
    wire N__6125;
    wire N__6122;
    wire N__6121;
    wire N__6120;
    wire N__6117;
    wire N__6112;
    wire N__6107;
    wire N__6104;
    wire N__6101;
    wire N__6098;
    wire N__6095;
    wire N__6092;
    wire N__6089;
    wire N__6086;
    wire N__6083;
    wire N__6082;
    wire N__6079;
    wire N__6076;
    wire N__6071;
    wire N__6068;
    wire N__6065;
    wire N__6064;
    wire N__6061;
    wire N__6058;
    wire N__6055;
    wire N__6052;
    wire N__6049;
    wire N__6046;
    wire N__6041;
    wire N__6038;
    wire N__6035;
    wire N__6032;
    wire N__6029;
    wire N__6026;
    wire N__6023;
    wire N__6020;
    wire N__6019;
    wire N__6016;
    wire N__6013;
    wire N__6010;
    wire N__6007;
    wire N__6004;
    wire N__6001;
    wire N__5998;
    wire N__5995;
    wire N__5992;
    wire N__5989;
    wire N__5984;
    wire N__5981;
    wire N__5978;
    wire N__5975;
    wire N__5972;
    wire N__5969;
    wire N__5966;
    wire N__5963;
    wire N__5960;
    wire N__5959;
    wire N__5956;
    wire N__5953;
    wire N__5950;
    wire N__5945;
    wire N__5942;
    wire N__5939;
    wire N__5936;
    wire N__5933;
    wire N__5930;
    wire N__5927;
    wire N__5924;
    wire N__5921;
    wire N__5918;
    wire N__5915;
    wire N__5912;
    wire N__5909;
    wire N__5906;
    wire N__5903;
    wire N__5900;
    wire N__5897;
    wire N__5894;
    wire N__5893;
    wire N__5892;
    wire N__5891;
    wire N__5890;
    wire N__5889;
    wire N__5888;
    wire N__5887;
    wire N__5884;
    wire N__5881;
    wire N__5872;
    wire N__5867;
    wire N__5858;
    wire N__5855;
    wire N__5854;
    wire N__5851;
    wire N__5850;
    wire N__5847;
    wire N__5844;
    wire N__5841;
    wire N__5838;
    wire N__5835;
    wire N__5832;
    wire N__5825;
    wire N__5822;
    wire N__5819;
    wire N__5816;
    wire N__5813;
    wire N__5810;
    wire N__5807;
    wire N__5804;
    wire N__5801;
    wire N__5798;
    wire N__5797;
    wire N__5796;
    wire N__5795;
    wire N__5792;
    wire N__5785;
    wire N__5780;
    wire N__5779;
    wire N__5776;
    wire N__5773;
    wire N__5768;
    wire N__5765;
    wire N__5762;
    wire N__5759;
    wire N__5756;
    wire N__5753;
    wire N__5750;
    wire N__5747;
    wire N__5744;
    wire N__5741;
    wire N__5738;
    wire N__5735;
    wire N__5732;
    wire N__5729;
    wire N__5726;
    wire N__5723;
    wire N__5722;
    wire N__5719;
    wire N__5716;
    wire N__5711;
    wire N__5710;
    wire N__5709;
    wire N__5706;
    wire N__5705;
    wire N__5702;
    wire N__5701;
    wire N__5700;
    wire N__5699;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5687;
    wire N__5684;
    wire N__5683;
    wire N__5682;
    wire N__5681;
    wire N__5678;
    wire N__5675;
    wire N__5668;
    wire N__5667;
    wire N__5666;
    wire N__5665;
    wire N__5662;
    wire N__5659;
    wire N__5656;
    wire N__5651;
    wire N__5646;
    wire N__5643;
    wire N__5636;
    wire N__5633;
    wire N__5618;
    wire N__5615;
    wire N__5614;
    wire N__5611;
    wire N__5608;
    wire N__5605;
    wire N__5602;
    wire N__5599;
    wire N__5596;
    wire N__5593;
    wire N__5590;
    wire N__5585;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5570;
    wire N__5567;
    wire N__5564;
    wire N__5563;
    wire N__5562;
    wire N__5559;
    wire N__5556;
    wire N__5553;
    wire N__5550;
    wire N__5547;
    wire N__5544;
    wire N__5541;
    wire N__5538;
    wire N__5535;
    wire N__5532;
    wire N__5529;
    wire N__5526;
    wire N__5523;
    wire N__5520;
    wire N__5517;
    wire N__5516;
    wire N__5513;
    wire N__5510;
    wire N__5507;
    wire N__5504;
    wire N__5495;
    wire N__5494;
    wire N__5493;
    wire N__5490;
    wire N__5485;
    wire N__5480;
    wire N__5479;
    wire N__5476;
    wire N__5473;
    wire N__5470;
    wire N__5465;
    wire N__5464;
    wire N__5463;
    wire N__5462;
    wire N__5461;
    wire N__5458;
    wire N__5449;
    wire N__5444;
    wire N__5441;
    wire N__5440;
    wire N__5439;
    wire N__5436;
    wire N__5431;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5416;
    wire N__5415;
    wire N__5412;
    wire N__5411;
    wire N__5410;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5396;
    wire N__5387;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5375;
    wire N__5374;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5362;
    wire N__5357;
    wire N__5354;
    wire N__5351;
    wire N__5348;
    wire N__5345;
    wire N__5342;
    wire N__5339;
    wire N__5336;
    wire N__5333;
    wire N__5332;
    wire N__5327;
    wire N__5324;
    wire N__5321;
    wire N__5320;
    wire N__5315;
    wire N__5312;
    wire N__5309;
    wire N__5306;
    wire N__5303;
    wire N__5302;
    wire N__5297;
    wire N__5294;
    wire N__5293;
    wire N__5290;
    wire N__5287;
    wire N__5284;
    wire N__5281;
    wire N__5278;
    wire N__5275;
    wire N__5272;
    wire N__5269;
    wire N__5266;
    wire N__5263;
    wire N__5258;
    wire N__5255;
    wire N__5252;
    wire N__5249;
    wire N__5246;
    wire N__5243;
    wire N__5240;
    wire N__5239;
    wire N__5238;
    wire N__5235;
    wire N__5232;
    wire N__5229;
    wire N__5224;
    wire N__5219;
    wire N__5216;
    wire N__5215;
    wire N__5212;
    wire N__5209;
    wire N__5208;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5196;
    wire N__5189;
    wire N__5188;
    wire N__5183;
    wire N__5180;
    wire N__5177;
    wire N__5174;
    wire N__5171;
    wire N__5168;
    wire N__5165;
    wire N__5162;
    wire N__5161;
    wire N__5158;
    wire N__5155;
    wire N__5152;
    wire N__5149;
    wire N__5146;
    wire N__5143;
    wire N__5138;
    wire N__5137;
    wire N__5134;
    wire N__5129;
    wire N__5126;
    wire N__5123;
    wire N__5120;
    wire N__5117;
    wire N__5114;
    wire N__5111;
    wire N__5108;
    wire N__5105;
    wire N__5102;
    wire N__5101;
    wire N__5098;
    wire N__5095;
    wire N__5090;
    wire N__5087;
    wire N__5084;
    wire N__5081;
    wire N__5080;
    wire N__5077;
    wire N__5074;
    wire N__5069;
    wire N__5066;
    wire N__5065;
    wire N__5062;
    wire N__5059;
    wire N__5054;
    wire N__5051;
    wire N__5050;
    wire N__5047;
    wire N__5044;
    wire N__5039;
    wire N__5036;
    wire N__5035;
    wire N__5032;
    wire N__5029;
    wire N__5026;
    wire N__5021;
    wire N__5018;
    wire N__5015;
    wire N__5012;
    wire N__5009;
    wire N__5008;
    wire N__5007;
    wire N__5006;
    wire N__5005;
    wire N__5004;
    wire N__5003;
    wire N__5002;
    wire N__5001;
    wire N__4982;
    wire N__4979;
    wire N__4976;
    wire N__4973;
    wire N__4970;
    wire N__4967;
    wire N__4964;
    wire N__4961;
    wire N__4958;
    wire N__4955;
    wire N__4954;
    wire N__4953;
    wire N__4950;
    wire N__4949;
    wire N__4944;
    wire N__4941;
    wire N__4938;
    wire N__4931;
    wire N__4928;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4916;
    wire N__4915;
    wire N__4912;
    wire N__4909;
    wire N__4904;
    wire N__4901;
    wire N__4898;
    wire N__4895;
    wire N__4892;
    wire N__4889;
    wire N__4886;
    wire N__4883;
    wire N__4882;
    wire N__4879;
    wire N__4878;
    wire N__4875;
    wire N__4872;
    wire N__4869;
    wire N__4866;
    wire N__4863;
    wire N__4860;
    wire N__4857;
    wire N__4854;
    wire N__4851;
    wire N__4848;
    wire N__4845;
    wire N__4842;
    wire N__4841;
    wire N__4840;
    wire N__4837;
    wire N__4834;
    wire N__4831;
    wire N__4828;
    wire N__4825;
    wire N__4816;
    wire N__4811;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4799;
    wire N__4798;
    wire N__4797;
    wire N__4796;
    wire N__4791;
    wire N__4786;
    wire N__4781;
    wire N__4778;
    wire N__4775;
    wire N__4774;
    wire N__4771;
    wire N__4768;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4750;
    wire N__4749;
    wire N__4748;
    wire N__4747;
    wire N__4746;
    wire N__4741;
    wire N__4736;
    wire N__4731;
    wire N__4724;
    wire N__4721;
    wire N__4718;
    wire N__4715;
    wire N__4712;
    wire N__4709;
    wire N__4706;
    wire N__4705;
    wire N__4702;
    wire N__4699;
    wire N__4696;
    wire N__4693;
    wire N__4690;
    wire N__4687;
    wire N__4682;
    wire N__4679;
    wire N__4676;
    wire N__4673;
    wire N__4670;
    wire N__4667;
    wire N__4666;
    wire N__4663;
    wire N__4660;
    wire N__4655;
    wire N__4652;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4640;
    wire N__4637;
    wire N__4634;
    wire N__4631;
    wire N__4628;
    wire N__4625;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4615;
    wire N__4614;
    wire N__4613;
    wire N__4608;
    wire N__4603;
    wire N__4598;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4586;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4573;
    wire N__4570;
    wire N__4567;
    wire N__4564;
    wire N__4561;
    wire N__4558;
    wire N__4555;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4541;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4523;
    wire N__4520;
    wire N__4517;
    wire N__4514;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire DBRn_c_i_0;
    wire CLK80_PLL_i_i;
    wire N_112_0;
    wire U712_REG_SM_REG_TACK_7_0;
    wire N_19_0_cascade_;
    wire U712_REG_SM_STATE_COUNT_3;
    wire N_19_0;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire C3_c;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire DBRn_c;
    wire DBR_SYNCZ0Z_0;
    wire VBENn_c;
    wire REG_TACK;
    wire U712_CHIP_RAM_m113_0;
    wire \U712_CHIP_RAM.N_87_0 ;
    wire \U712_CHIP_RAM.N_87_0_cascade_ ;
    wire \U712_CHIP_RAM.N_97_0_cascade_ ;
    wire U712_REG_SM_STATE_COUNT_7;
    wire U712_REG_SM_STATE_COUNT_0;
    wire \U712_CHIP_RAM.N_79_0 ;
    wire U712_REG_SM_STATE_COUNT_5;
    wire \U712_REG_SM.STATE_COUNTZ0Z_6 ;
    wire \U712_CHIP_RAM.N_103_0 ;
    wire U712_REG_SM_STATE_COUNT_8;
    wire \U712_CHIP_RAM.N_103_0_cascade_ ;
    wire \U712_CHIP_RAM.m106_nsZ0Z_1 ;
    wire i62_mux;
    wire U712_REG_SM_WRITE_CYCLE;
    wire PRnW_c;
    wire \U712_CHIP_RAM.N_332 ;
    wire \INVU712_CYCLE_TERM.TACK_ENC_net ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_2 ;
    wire TACK_EN;
    wire \U712_CYCLE_TERM.TACK_RST_0_i ;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire bfn_9_11_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire C1_c_g;
    wire REGSPACEn_c;
    wire U712_REG_SM_REG_CYCLE_START;
    wire U712_REG_SM_START_RST;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_3 ;
    wire RAMENn_c;
    wire TSn_c;
    wire \U712_CHIP_RAM.m223_ns_1_cascade_ ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_5 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_4 ;
    wire C1_c;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.m231_0 ;
    wire \U712_CHIP_RAM.N_236 ;
    wire U712_REG_SM_STATE_COUNT_0_sqmuxa_1;
    wire \U712_CHIP_RAM.N_83_0_cascade_ ;
    wire \U712_CHIP_RAM.N_83_0 ;
    wire \U712_CHIP_RAM.N_94_0_cascade_ ;
    wire U712_REG_SM_STATE_COUNT_1;
    wire U712_REG_SM_STATE_COUNT_2;
    wire DBR_SYNC_i_1;
    wire bfn_9_16_0_;
    wire \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1 ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2 ;
    wire \U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ;
    wire \U712_CHIP_RAM.CAS_COUNTERZ1Z_1 ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3 ;
    wire \U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.N_7_0 ;
    wire N_86_0;
    wire U712_REG_SM_C3_SYNC_1;
    wire BLSn_c;
    wire \U712_REG_SM.N_86_0_0 ;
    wire \U712_CYCLE_TERM.N_36_0_cascade_ ;
    wire TACK_OUT;
    wire \U712_CYCLE_TERM.TACK_STARTZ0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \INVU712_CYCLE_TERM.TACK_OUTC_net ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0 ;
    wire \U712_CHIP_RAM.N_146_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_3_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_3 ;
    wire \U712_CHIP_RAM.N_154_0_cascade_ ;
    wire \U712_CHIP_RAM.m38_1 ;
    wire \U712_CHIP_RAM.N_34_0_cascade_ ;
    wire \U712_CHIP_RAM.N_359 ;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_28_0_cascade_ ;
    wire \U712_CHIP_RAM.N_47_0_cascade_ ;
    wire \U712_CHIP_RAM.N_215 ;
    wire bfn_10_14_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.N_56_0_i ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire \U712_CHIP_RAM.N_330 ;
    wire \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ;
    wire U712_REG_SM_UDSn_6_0;
    wire UDSn_c;
    wire DBRn_c_i;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ;
    wire CMA_c_8;
    wire A_c_9;
    wire \U712_CHIP_RAM.m186_0_cascade_ ;
    wire A_c_17;
    wire \U712_CHIP_RAM.m192_0_cascade_ ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.m192_1 ;
    wire \U712_CHIP_RAM.d_N_6_5 ;
    wire \U712_CHIP_RAM.d_N_6_1 ;
    wire \U712_CHIP_RAM.N_353_mux ;
    wire \U712_CHIP_RAM.N_168_0_cascade_ ;
    wire \U712_CHIP_RAM.m64_ns_1 ;
    wire \U712_CHIP_RAM.i67_mux_cascade_ ;
    wire \U712_CHIP_RAM.m66_ns_1 ;
    wire \U712_CHIP_RAM.N_146_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_2_cascade_ ;
    wire \U712_CHIP_RAM.N_151_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_2 ;
    wire A_c_2;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ;
    wire A_c_20;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH5lt7 ;
    wire \U712_CHIP_RAM.N_28_0 ;
    wire \U712_CHIP_RAM.N_219 ;
    wire \U712_CHIP_RAM.m41_1 ;
    wire \U712_CHIP_RAM.N_31_0_cascade_ ;
    wire \U712_CHIP_RAM.m217_ns_1_cascade_ ;
    wire \U712_CHIP_RAM.N_218 ;
    wire \U712_CHIP_RAM.m212_ns_1_cascade_ ;
    wire \U712_CHIP_RAM.N_30_0_cascade_ ;
    wire \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0 ;
    wire \U712_CHIP_RAM.N_213 ;
    wire CPU_TACKm;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.N_333_mux_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.N_51_0 ;
    wire \U712_CHIP_RAM.N_51_0_cascade_ ;
    wire \U712_CHIP_RAM.N_54_0 ;
    wire \U712_CHIP_RAM.m53_ns_1 ;
    wire \U712_CHIP_RAM.N_333_mux ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0 ;
    wire DBR_SYNCZ0Z_1;
    wire \U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ;
    wire CMA_c_4;
    wire CMA_c_3;
    wire CMA_c_10;
    wire \U712_CHIP_RAM.m189_1 ;
    wire \U712_CHIP_RAM.m188_1 ;
    wire \U712_CHIP_RAM.d_N_6_2 ;
    wire A_c_12;
    wire \U712_CHIP_RAM.m188_0 ;
    wire \U712_CHIP_RAM.d_N_6 ;
    wire A_c_13;
    wire \U712_CHIP_RAM.m189_0 ;
    wire A_c_14;
    wire CMA_c_2;
    wire \U712_CHIP_RAM.m186_1 ;
    wire CMA_c_0;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.N_198_cascade_ ;
    wire CLK40_PLL;
    wire CLK40_PLL_iso_i;
    wire \U712_CHIP_RAM.m187_1 ;
    wire A_c_11;
    wire \U712_CHIP_RAM.N_3_0_cascade_ ;
    wire \U712_CHIP_RAM.m187_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_1 ;
    wire \U712_CHIP_RAM.N_163_0_cascade_ ;
    wire \U712_CHIP_RAM.N_67_0 ;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.N_48_0 ;
    wire \U712_CHIP_RAM.N_363 ;
    wire \U712_CHIP_RAM.N_158_0_cascade_ ;
    wire \U712_CHIP_RAM.N_58_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_1 ;
    wire \U712_CHIP_RAM.d_N_6_0 ;
    wire \U712_CHIP_RAM.N_43_0 ;
    wire A_c_4;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ;
    wire A_c_5;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ;
    wire A_c_6;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ;
    wire A_c_7;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_START_RNIJD6OZ0Z3_cascade_ ;
    wire \U712_CHIP_RAM.N_204_cascade_ ;
    wire \U712_CHIP_RAM.N_364 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_ ;
    wire DBDIR_c;
    wire \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ;
    wire AWEn_c;
    wire \U712_CHIP_RAM.N_26_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.N_30_0 ;
    wire \U712_CHIP_RAM.N_62_0_cascade_ ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_RNI9THUZ0Z5 ;
    wire \U712_CHIP_RAM.CLK_EN_RNOZ0Z_2_cascade_ ;
    wire \U712_CHIP_RAM.CLK_EN_RNOZ0Z_3 ;
    wire \U712_CHIP_RAM.N_174_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER43 ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.WRITE_CYCLEZ0 ;
    wire \U712_CHIP_RAM.N_62_0 ;
    wire \U712_CHIP_RAM.N_52_0 ;
    wire \U712_CHIP_RAM.N_208_cascade_ ;
    wire N_99_0;
    wire LDSn_c;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire RESETn_c;
    wire RESETn_c_i;
    wire RASn_c;
    wire \U712_CHIP_RAM.d_N_7 ;
    wire \U712_CHIP_RAM.m185_0 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ;
    wire A_c_16;
    wire \U712_CHIP_RAM.m191_0_cascade_ ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.d_N_6_4 ;
    wire A_c_10;
    wire \U712_CHIP_RAM.m184_m2_0_a2_0 ;
    wire \U712_CHIP_RAM.m184_0_cascade_ ;
    wire \U712_CHIP_RAM.m184_1 ;
    wire A_c_15;
    wire \U712_CHIP_RAM.N_3_0 ;
    wire \U712_CHIP_RAM.m186_m2_0_a2_0 ;
    wire \U712_CHIP_RAM.m190_0_cascade_ ;
    wire \U712_CHIP_RAM.m190_1 ;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.d_N_6_3 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire \U712_CHIP_RAM.d_N_7_0 ;
    wire A_c_18;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.N_204 ;
    wire A_c_3;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ;
    wire A_c_8;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.N_31_0 ;
    wire \U712_CHIP_RAM.DBENn_8_0 ;
    wire CONSTANT_ONE_NET;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0 ;
    wire LATCH_CLK_c;
    wire ASn_c;
    wire \U712_REG_SM.N_99_0_0 ;
    wire U712_REG_SM_C1_SYNC_1;
    wire U712_REG_SM_LDSn_6_0;
    wire \U712_CHIP_RAM.m185_1 ;
    wire CMA_c_5;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire A_c_19;
    wire \U712_CHIP_RAM.m194_0 ;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.m191_1 ;
    wire CMA_c_7;
    wire \U712_CHIP_RAM.N_198_0 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire CUMBEn_c;
    wire LMBEn_c;
    wire CLMBEn_c;
    wire CUUBEn_c;
    wire \U712_CHIP_RAM.N_346 ;
    wire DBENn_c;
    wire \U712_CHIP_RAM.N_346_cascade_ ;
    wire CLLBEn_c;
    wire LLBEn_c;
    wire A_c_0;
    wire UUBEn_c;
    wire SIZ_c_0;
    wire A_c_1;
    wire SIZ_c_1;
    wire \U712_CHIP_RAM.N_325_mux ;
    wire UMBEn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire WEn_c;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ;
    wire DRA_c_6;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire DRA_c_0;
    wire DRA_c_1;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \INVU712_CHIP_RAM.DMA_A1_nesrC_net ;
    wire \U712_CHIP_RAM.DMA_CYCLEm ;
    wire \U712_CHIP_RAM.N_345 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire DMA_LATCH_EN_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire CASn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CRCSn_c;
    wire DRA_c_8;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire DRA_c_9;
    wire AGNUS_REV_c;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire C3_c_g;
    wire DBRn_c_i_0_g;
    wire RAS0n_c;
    wire RAS1n_c;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_0 ;
    wire CLK80_PLL;
    wire RESETn_c_i_g;
    wire REG_CYCLEm;
    wire \U712_CHIP_RAM.CPU_CYCLEm ;
    wire N_338_mux;
    wire CASLn_c;
    wire RnW_c;
    wire \U712_CHIP_RAM.DMA_WRITE_CYCLEZ0 ;
    wire CASUn_c;
    wire N_328_mux;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL),
            .REFERENCECLK(N__4511),
            .RESETB(N__8729),
            .BYPASS(GNDG0),
            .PLLOUTCOREA(),
            .SDI(GNDG0),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(GNDG0),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK(GNDG0));
    IO_PAD DBENn_obuf_iopad (
            .OE(N__13161),
            .DIN(N__13160),
            .DOUT(N__13159),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__13161),
            .PADOUT(N__13160),
            .PADIN(N__13159),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10274),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__13152),
            .DIN(N__13151),
            .DOUT(N__13150),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__13152),
            .PADOUT(N__13151),
            .PADIN(N__13150),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__13143),
            .DIN(N__13142),
            .DOUT(N__13141),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__13143),
            .PADOUT(N__13142),
            .PADIN(N__13141),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12026),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__13134),
            .DIN(N__13133),
            .DOUT(N__13132),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__13134),
            .PADOUT(N__13133),
            .PADIN(N__13132),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10661),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__13125),
            .DIN(N__13124),
            .DOUT(N__13123),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__13125),
            .PADOUT(N__13124),
            .PADIN(N__13123),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__13116),
            .DIN(N__13115),
            .DOUT(N__13114),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__13116),
            .PADOUT(N__13115),
            .PADIN(N__13114),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__13107),
            .DIN(N__13106),
            .DOUT(N__13105),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__13107),
            .PADOUT(N__13106),
            .PADIN(N__13105),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__13098),
            .DIN(N__13097),
            .DOUT(N__13096),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__13098),
            .PADOUT(N__13097),
            .PADIN(N__13096),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__13089),
            .DIN(N__13088),
            .DOUT(N__13087),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__13089),
            .PADOUT(N__13088),
            .PADIN(N__13087),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS1n_ibuf_iopad (
            .OE(N__13080),
            .DIN(N__13079),
            .DOUT(N__13078),
            .PACKAGEPIN(RAS1n));
    defparam RAS1n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS1n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS1n_ibuf_preio (
            .PADOEN(N__13080),
            .PADOUT(N__13079),
            .PADIN(N__13078),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS1n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__13071),
            .DIN(N__13070),
            .DOUT(N__13069),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__13071),
            .PADOUT(N__13070),
            .PADIN(N__13069),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__13062),
            .DIN(N__13061),
            .DOUT(N__13060),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__13062),
            .PADOUT(N__13061),
            .PADIN(N__13060),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9692),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__13053),
            .DIN(N__13052),
            .DOUT(N__13051),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__13053),
            .PADOUT(N__13052),
            .PADIN(N__13051),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10121),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__13044),
            .DIN(N__13043),
            .DOUT(N__13042),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__13044),
            .PADOUT(N__13043),
            .PADIN(N__13042),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMENn_obuf_iopad (
            .OE(N__13035),
            .DIN(N__13034),
            .DOUT(N__13033),
            .PACKAGEPIN(RAMENn));
    defparam RAMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMENn_obuf_preio (
            .PADOEN(N__13035),
            .PADOUT(N__13034),
            .PADIN(N__13033),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5161),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__13026),
            .DIN(N__13025),
            .DOUT(N__13024),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__13026),
            .PADOUT(N__13025),
            .PADIN(N__13024),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__13017),
            .DIN(N__13016),
            .DOUT(N__13015),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__13017),
            .PADOUT(N__13016),
            .PADIN(N__13015),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__13008),
            .DIN(N__13007),
            .DOUT(N__13006),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__13008),
            .PADOUT(N__13007),
            .PADIN(N__13006),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4676),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__12999),
            .DIN(N__12998),
            .DOUT(N__12997),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__12999),
            .PADOUT(N__12998),
            .PADIN(N__12997),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__12990),
            .DIN(N__12989),
            .DOUT(N__12988),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__12990),
            .PADOUT(N__12989),
            .PADIN(N__12988),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__12981),
            .DIN(N__12980),
            .DOUT(N__12979),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__12981),
            .PADOUT(N__12980),
            .PADIN(N__12979),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6905),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__12972),
            .DIN(N__12971),
            .DOUT(N__12970),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__12972),
            .PADOUT(N__12971),
            .PADIN(N__12970),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__12963),
            .DIN(N__12962),
            .DOUT(N__12961),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__12963),
            .PADOUT(N__12962),
            .PADIN(N__12961),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11960),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__12954),
            .DIN(N__12953),
            .DOUT(N__12952),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__12954),
            .PADOUT(N__12953),
            .PADIN(N__12952),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__12945),
            .DIN(N__12944),
            .DOUT(N__12943),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__12945),
            .PADOUT(N__12944),
            .PADIN(N__12943),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10193),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_obuft_iopad (
            .OE(N__12936),
            .DIN(N__12935),
            .DOUT(N__12934),
            .PACKAGEPIN(TBIn));
    defparam TBIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TBIn_obuft_preio (
            .PADOEN(N__12936),
            .PADOUT(N__12935),
            .PADIN(N__12934),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4878),
            .DIN0(),
            .DOUT0(N__5562),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__12927),
            .DIN(N__12926),
            .DOUT(N__12925),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__12927),
            .PADOUT(N__12926),
            .PADIN(N__12925),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__12918),
            .DIN(N__12917),
            .DOUT(N__12916),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__12918),
            .PADOUT(N__12917),
            .PADIN(N__12916),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__12909),
            .DIN(N__12908),
            .DOUT(N__12907),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__12909),
            .PADOUT(N__12908),
            .PADIN(N__12907),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__12900),
            .DIN(N__12899),
            .DOUT(N__12898),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__12900),
            .PADOUT(N__12899),
            .PADIN(N__12898),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__12891),
            .DIN(N__12890),
            .DOUT(N__12889),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__12891),
            .PADOUT(N__12890),
            .PADIN(N__12889),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_EN_obuf_iopad (
            .OE(N__12882),
            .DIN(N__12881),
            .DOUT(N__12880),
            .PACKAGEPIN(DMA_LATCH_EN));
    defparam DMA_LATCH_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_EN_obuf_preio (
            .PADOEN(N__12882),
            .PADOUT(N__12881),
            .PADIN(N__12880),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12269),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__12873),
            .DIN(N__12872),
            .DOUT(N__12871),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__12873),
            .PADOUT(N__12872),
            .PADIN(N__12871),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__12864),
            .DIN(N__12863),
            .DOUT(N__12862),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__12864),
            .PADOUT(N__12863),
            .PADIN(N__12862),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__12855),
            .DIN(N__12854),
            .DOUT(N__12853),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__12855),
            .PADOUT(N__12854),
            .PADIN(N__12853),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__12846),
            .DIN(N__12845),
            .DOUT(N__12844),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__12846),
            .PADOUT(N__12845),
            .PADIN(N__12844),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__12837),
            .DIN(N__12836),
            .DOUT(N__12835),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__12837),
            .PADOUT(N__12836),
            .PADIN(N__12835),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__12828),
            .DIN(N__12827),
            .DOUT(N__12826),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__12828),
            .PADOUT(N__12827),
            .PADIN(N__12826),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7910),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__12819),
            .DIN(N__12818),
            .DOUT(N__12817),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__12819),
            .PADOUT(N__12818),
            .PADIN(N__12817),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__12810),
            .DIN(N__12809),
            .DOUT(N__12808),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__12810),
            .PADOUT(N__12809),
            .PADIN(N__12808),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__12801),
            .DIN(N__12800),
            .DOUT(N__12799),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__12801),
            .PADOUT(N__12800),
            .PADIN(N__12799),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9485),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_0_iopad (
            .OE(N__12792),
            .DIN(N__12791),
            .DOUT(N__12790),
            .PACKAGEPIN(DA[0]));
    defparam DA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_0_preio (
            .PADOEN(N__12792),
            .PADOUT(N__12791),
            .PADIN(N__12790),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6020),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__12783),
            .DIN(N__12782),
            .DOUT(N__12781),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__12783),
            .PADOUT(N__12782),
            .PADIN(N__12781),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__12774),
            .DIN(N__12773),
            .DOUT(N__12772),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__12774),
            .PADOUT(N__12773),
            .PADIN(N__12772),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6722),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__12765),
            .DIN(N__12764),
            .DOUT(N__12763),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__12765),
            .PADOUT(N__12764),
            .PADIN(N__12763),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6770),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__12756),
            .DIN(N__12755),
            .DOUT(N__12754),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__12756),
            .PADOUT(N__12755),
            .PADIN(N__12754),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5614),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__12747),
            .DIN(N__12746),
            .DOUT(N__12745),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__12747),
            .PADOUT(N__12746),
            .PADIN(N__12745),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__12738),
            .DIN(N__12737),
            .DOUT(N__12736),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__12738),
            .PADOUT(N__12737),
            .PADIN(N__12736),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9524),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_obuft_iopad (
            .OE(N__12729),
            .DIN(N__12728),
            .DOUT(N__12727),
            .PACKAGEPIN(TCIn));
    defparam TCIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TCIn_obuft_preio (
            .PADOEN(N__12729),
            .PADOUT(N__12728),
            .PADIN(N__12727),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4883),
            .DIN0(),
            .DOUT0(N__5563),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__12720),
            .DIN(N__12719),
            .DOUT(N__12718),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__12720),
            .PADOUT(N__12719),
            .PADIN(N__12718),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9821),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__12711),
            .DIN(N__12710),
            .DOUT(N__12709),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__12711),
            .PADOUT(N__12710),
            .PADIN(N__12709),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7235),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__12702),
            .DIN(N__12701),
            .DOUT(N__12700),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__12702),
            .PADOUT(N__12701),
            .PADIN(N__12700),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9578),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__12693),
            .DIN(N__12692),
            .DOUT(N__12691),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__12693),
            .PADOUT(N__12692),
            .PADIN(N__12691),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__12684),
            .DIN(N__12683),
            .DOUT(N__12682),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__12684),
            .PADOUT(N__12683),
            .PADIN(N__12682),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_2_iopad (
            .OE(N__12675),
            .DIN(N__12674),
            .DOUT(N__12673),
            .PACKAGEPIN(DA[2]));
    defparam DA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_2_preio (
            .PADOEN(N__12675),
            .PADOUT(N__12674),
            .PADIN(N__12673),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7205),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__12666),
            .DIN(N__12665),
            .DOUT(N__12664),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__12666),
            .PADOUT(N__12665),
            .PADIN(N__12664),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__12657),
            .DIN(N__12656),
            .DOUT(N__12655),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__12657),
            .PADOUT(N__12656),
            .PADIN(N__12655),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__12648),
            .DIN(N__12647),
            .DOUT(N__12646),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__12648),
            .PADOUT(N__12647),
            .PADIN(N__12646),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6884),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__12639),
            .DIN(N__12638),
            .DOUT(N__12637),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__12639),
            .PADOUT(N__12638),
            .PADIN(N__12637),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9554),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__12630),
            .DIN(N__12629),
            .DOUT(N__12628),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__12630),
            .PADOUT(N__12629),
            .PADIN(N__12628),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__12621),
            .DIN(N__12620),
            .DOUT(N__12619),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__12621),
            .PADOUT(N__12620),
            .PADIN(N__12619),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9503),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__12612),
            .DIN(N__12611),
            .DOUT(N__12610),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__12612),
            .PADOUT(N__12611),
            .PADIN(N__12610),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4882),
            .DIN0(),
            .DOUT0(N__5564),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__12603),
            .DIN(N__12602),
            .DOUT(N__12601),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__12603),
            .PADOUT(N__12602),
            .PADIN(N__12601),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6929),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__12594),
            .DIN(N__12593),
            .DOUT(N__12592),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__12594),
            .PADOUT(N__12593),
            .PADIN(N__12592),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__12585),
            .DIN(N__12584),
            .DOUT(N__12583),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__12585),
            .PADOUT(N__12584),
            .PADIN(N__12583),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__12576),
            .DIN(N__12575),
            .DOUT(N__12574),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__12576),
            .PADOUT(N__12575),
            .PADIN(N__12574),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6041),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__12567),
            .DIN(N__12566),
            .DOUT(N__12565),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__12567),
            .PADOUT(N__12566),
            .PADIN(N__12565),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__12558),
            .DIN(N__12557),
            .DOUT(N__12556),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__12558),
            .PADOUT(N__12557),
            .PADIN(N__12556),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_1_iopad (
            .OE(N__12549),
            .DIN(N__12548),
            .DOUT(N__12547),
            .PACKAGEPIN(DA[1]));
    defparam DA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_1_preio (
            .PADOEN(N__12549),
            .PADOUT(N__12548),
            .PADIN(N__12547),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8471),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__12540),
            .DIN(N__12539),
            .DOUT(N__12538),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__12540),
            .PADOUT(N__12539),
            .PADIN(N__12538),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__12531),
            .DIN(N__12530),
            .DOUT(N__12529),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__12531),
            .PADOUT(N__12530),
            .PADIN(N__12529),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__12522),
            .DIN(N__12521),
            .DOUT(N__12520),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__12522),
            .PADOUT(N__12521),
            .PADIN(N__12520),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9329),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__12513),
            .DIN(N__12512),
            .DOUT(N__12511),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__12513),
            .PADOUT(N__12512),
            .PADIN(N__12511),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6098),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__12504),
            .DIN(N__12503),
            .DOUT(N__12502),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__12504),
            .PADOUT(N__12503),
            .PADIN(N__12502),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9923),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__12495),
            .DIN(N__12494),
            .DOUT(N__12493),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__12495),
            .PADOUT(N__12494),
            .PADIN(N__12493),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7613),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__12486),
            .DIN(N__12485),
            .DOUT(N__12484),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__12486),
            .PADOUT(N__12485),
            .PADIN(N__12484),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__12477),
            .DIN(N__12476),
            .DOUT(N__12475),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__12477),
            .PADOUT(N__12476),
            .PADIN(N__12475),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__12468),
            .DIN(N__12467),
            .DOUT(N__12466),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__12468),
            .PADOUT(N__12467),
            .PADIN(N__12466),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8243),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__12459),
            .DIN(N__12458),
            .DOUT(N__12457),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__12459),
            .PADOUT(N__12458),
            .PADIN(N__12457),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__12450),
            .DIN(N__12449),
            .DOUT(N__12448),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__12450),
            .PADOUT(N__12449),
            .PADIN(N__12448),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__12441),
            .DIN(N__12440),
            .DOUT(N__12439),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__12441),
            .PADOUT(N__12440),
            .PADIN(N__12439),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8507),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__12432),
            .DIN(N__12431),
            .DOUT(N__12430),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__12432),
            .PADOUT(N__12431),
            .PADIN(N__12430),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8177),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__12423),
            .DIN(N__12422),
            .DOUT(N__12421),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__12423),
            .PADOUT(N__12422),
            .PADIN(N__12421),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6831),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PRnW_obuf_iopad (
            .OE(N__12414),
            .DIN(N__12413),
            .DOUT(N__12412),
            .PACKAGEPIN(PRnW));
    defparam PRnW_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PRnW_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PRnW_obuf_preio (
            .PADOEN(N__12414),
            .PADOUT(N__12413),
            .PADIN(N__12412),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4931),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__12405),
            .DIN(N__12404),
            .DOUT(N__12403),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__12405),
            .PADOUT(N__12404),
            .PADIN(N__12403),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__12396),
            .DIN(N__12395),
            .DOUT(N__12394),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__12396),
            .PADOUT(N__12395),
            .PADIN(N__12394),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6833),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__12387),
            .DIN(N__12386),
            .DOUT(N__12385),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__12387),
            .PADOUT(N__12386),
            .PADIN(N__12385),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4526),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__12378),
            .DIN(N__12377),
            .DOUT(N__12376),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__12378),
            .PADOUT(N__12377),
            .PADIN(N__12376),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6746),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__12369),
            .DIN(N__12368),
            .DOUT(N__12367),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__12369),
            .PADOUT(N__12368),
            .PADIN(N__12367),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__12360),
            .DIN(N__12359),
            .DOUT(N__12358),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__12360),
            .PADOUT(N__12359),
            .PADIN(N__12358),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__12351),
            .DIN(N__12350),
            .DOUT(N__12349),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__12351),
            .PADOUT(N__12350),
            .PADIN(N__12349),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BLSn_obuf_iopad (
            .OE(N__12342),
            .DIN(N__12341),
            .DOUT(N__12340),
            .PACKAGEPIN(BLSn));
    defparam BLSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BLSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BLSn_obuf_preio (
            .PADOEN(N__12342),
            .PADOUT(N__12341),
            .PADIN(N__12340),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5618),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__12333),
            .DIN(N__12332),
            .DOUT(N__12331),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__12333),
            .PADOUT(N__12332),
            .PADIN(N__12331),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__12324),
            .DIN(N__12323),
            .DOUT(N__12322),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__12324),
            .PADOUT(N__12323),
            .PADIN(N__12322),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6832),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__12315),
            .DIN(N__12314),
            .DOUT(N__12313),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__12315),
            .PADOUT(N__12314),
            .PADIN(N__12313),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10871),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__12306),
            .DIN(N__12305),
            .DOUT(N__12304),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__12306),
            .PADOUT(N__12305),
            .PADIN(N__12304),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10214),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__12297),
            .DIN(N__12296),
            .DOUT(N__12295),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__12297),
            .PADOUT(N__12296),
            .PADIN(N__12295),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9263),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__12288),
            .DIN(N__12287),
            .DOUT(N__12286),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__12288),
            .PADOUT(N__12287),
            .PADIN(N__12286),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IoInMux I__2982 (
            .O(N__12269),
            .I(N__12266));
    LocalMux I__2981 (
            .O(N__12266),
            .I(N__12263));
    Span4Mux_s3_v I__2980 (
            .O(N__12263),
            .I(N__12260));
    Span4Mux_v I__2979 (
            .O(N__12260),
            .I(N__12257));
    Sp12to4 I__2978 (
            .O(N__12257),
            .I(N__12254));
    Span12Mux_h I__2977 (
            .O(N__12254),
            .I(N__12251));
    Odrv12 I__2976 (
            .O(N__12251),
            .I(DMA_LATCH_EN_c));
    CascadeMux I__2975 (
            .O(N__12248),
            .I(N__12244));
    InMux I__2974 (
            .O(N__12247),
            .I(N__12237));
    InMux I__2973 (
            .O(N__12244),
            .I(N__12234));
    CascadeMux I__2972 (
            .O(N__12243),
            .I(N__12231));
    CascadeMux I__2971 (
            .O(N__12242),
            .I(N__12221));
    CascadeMux I__2970 (
            .O(N__12241),
            .I(N__12218));
    CascadeMux I__2969 (
            .O(N__12240),
            .I(N__12215));
    LocalMux I__2968 (
            .O(N__12237),
            .I(N__12209));
    LocalMux I__2967 (
            .O(N__12234),
            .I(N__12209));
    InMux I__2966 (
            .O(N__12231),
            .I(N__12206));
    InMux I__2965 (
            .O(N__12230),
            .I(N__12203));
    CascadeMux I__2964 (
            .O(N__12229),
            .I(N__12200));
    CascadeMux I__2963 (
            .O(N__12228),
            .I(N__12196));
    CascadeMux I__2962 (
            .O(N__12227),
            .I(N__12193));
    CascadeMux I__2961 (
            .O(N__12226),
            .I(N__12190));
    CascadeMux I__2960 (
            .O(N__12225),
            .I(N__12187));
    CascadeMux I__2959 (
            .O(N__12224),
            .I(N__12178));
    InMux I__2958 (
            .O(N__12221),
            .I(N__12171));
    InMux I__2957 (
            .O(N__12218),
            .I(N__12171));
    InMux I__2956 (
            .O(N__12215),
            .I(N__12171));
    InMux I__2955 (
            .O(N__12214),
            .I(N__12168));
    Span4Mux_h I__2954 (
            .O(N__12209),
            .I(N__12165));
    LocalMux I__2953 (
            .O(N__12206),
            .I(N__12160));
    LocalMux I__2952 (
            .O(N__12203),
            .I(N__12157));
    InMux I__2951 (
            .O(N__12200),
            .I(N__12154));
    InMux I__2950 (
            .O(N__12199),
            .I(N__12141));
    InMux I__2949 (
            .O(N__12196),
            .I(N__12141));
    InMux I__2948 (
            .O(N__12193),
            .I(N__12141));
    InMux I__2947 (
            .O(N__12190),
            .I(N__12134));
    InMux I__2946 (
            .O(N__12187),
            .I(N__12134));
    InMux I__2945 (
            .O(N__12186),
            .I(N__12134));
    InMux I__2944 (
            .O(N__12185),
            .I(N__12127));
    InMux I__2943 (
            .O(N__12184),
            .I(N__12127));
    InMux I__2942 (
            .O(N__12183),
            .I(N__12127));
    CascadeMux I__2941 (
            .O(N__12182),
            .I(N__12124));
    CascadeMux I__2940 (
            .O(N__12181),
            .I(N__12115));
    InMux I__2939 (
            .O(N__12178),
            .I(N__12112));
    LocalMux I__2938 (
            .O(N__12171),
            .I(N__12107));
    LocalMux I__2937 (
            .O(N__12168),
            .I(N__12107));
    Span4Mux_v I__2936 (
            .O(N__12165),
            .I(N__12104));
    InMux I__2935 (
            .O(N__12164),
            .I(N__12099));
    InMux I__2934 (
            .O(N__12163),
            .I(N__12099));
    Span4Mux_h I__2933 (
            .O(N__12160),
            .I(N__12092));
    Span4Mux_v I__2932 (
            .O(N__12157),
            .I(N__12092));
    LocalMux I__2931 (
            .O(N__12154),
            .I(N__12092));
    InMux I__2930 (
            .O(N__12153),
            .I(N__12085));
    InMux I__2929 (
            .O(N__12152),
            .I(N__12085));
    InMux I__2928 (
            .O(N__12151),
            .I(N__12085));
    InMux I__2927 (
            .O(N__12150),
            .I(N__12080));
    InMux I__2926 (
            .O(N__12149),
            .I(N__12080));
    InMux I__2925 (
            .O(N__12148),
            .I(N__12077));
    LocalMux I__2924 (
            .O(N__12141),
            .I(N__12070));
    LocalMux I__2923 (
            .O(N__12134),
            .I(N__12070));
    LocalMux I__2922 (
            .O(N__12127),
            .I(N__12070));
    InMux I__2921 (
            .O(N__12124),
            .I(N__12063));
    InMux I__2920 (
            .O(N__12123),
            .I(N__12063));
    InMux I__2919 (
            .O(N__12122),
            .I(N__12063));
    InMux I__2918 (
            .O(N__12121),
            .I(N__12056));
    InMux I__2917 (
            .O(N__12120),
            .I(N__12056));
    InMux I__2916 (
            .O(N__12119),
            .I(N__12056));
    InMux I__2915 (
            .O(N__12118),
            .I(N__12051));
    InMux I__2914 (
            .O(N__12115),
            .I(N__12051));
    LocalMux I__2913 (
            .O(N__12112),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2912 (
            .O(N__12107),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2911 (
            .O(N__12104),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2910 (
            .O(N__12099),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2909 (
            .O(N__12092),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2908 (
            .O(N__12085),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2907 (
            .O(N__12080),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2906 (
            .O(N__12077),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv12 I__2905 (
            .O(N__12070),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2904 (
            .O(N__12063),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2903 (
            .O(N__12056),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2902 (
            .O(N__12051),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    IoInMux I__2901 (
            .O(N__12026),
            .I(N__12023));
    LocalMux I__2900 (
            .O(N__12023),
            .I(N__12020));
    Span12Mux_s9_v I__2899 (
            .O(N__12020),
            .I(N__12017));
    Odrv12 I__2898 (
            .O(N__12017),
            .I(CASn_c));
    InMux I__2897 (
            .O(N__12014),
            .I(N__12010));
    InMux I__2896 (
            .O(N__12013),
            .I(N__12007));
    LocalMux I__2895 (
            .O(N__12010),
            .I(N__12003));
    LocalMux I__2894 (
            .O(N__12007),
            .I(N__12000));
    CascadeMux I__2893 (
            .O(N__12006),
            .I(N__11997));
    Span4Mux_h I__2892 (
            .O(N__12003),
            .I(N__11991));
    Span4Mux_h I__2891 (
            .O(N__12000),
            .I(N__11991));
    InMux I__2890 (
            .O(N__11997),
            .I(N__11988));
    InMux I__2889 (
            .O(N__11996),
            .I(N__11985));
    Span4Mux_v I__2888 (
            .O(N__11991),
            .I(N__11979));
    LocalMux I__2887 (
            .O(N__11988),
            .I(N__11979));
    LocalMux I__2886 (
            .O(N__11985),
            .I(N__11976));
    InMux I__2885 (
            .O(N__11984),
            .I(N__11973));
    Span4Mux_h I__2884 (
            .O(N__11979),
            .I(N__11970));
    Span4Mux_h I__2883 (
            .O(N__11976),
            .I(N__11967));
    LocalMux I__2882 (
            .O(N__11973),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__2881 (
            .O(N__11970),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__2880 (
            .O(N__11967),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__2879 (
            .O(N__11960),
            .I(N__11957));
    LocalMux I__2878 (
            .O(N__11957),
            .I(N__11954));
    Span4Mux_s1_v I__2877 (
            .O(N__11954),
            .I(N__11951));
    Span4Mux_v I__2876 (
            .O(N__11951),
            .I(N__11948));
    Span4Mux_v I__2875 (
            .O(N__11948),
            .I(N__11945));
    Odrv4 I__2874 (
            .O(N__11945),
            .I(CRCSn_c));
    InMux I__2873 (
            .O(N__11942),
            .I(N__11939));
    LocalMux I__2872 (
            .O(N__11939),
            .I(N__11933));
    InMux I__2871 (
            .O(N__11938),
            .I(N__11930));
    InMux I__2870 (
            .O(N__11937),
            .I(N__11927));
    InMux I__2869 (
            .O(N__11936),
            .I(N__11924));
    Span4Mux_v I__2868 (
            .O(N__11933),
            .I(N__11921));
    LocalMux I__2867 (
            .O(N__11930),
            .I(N__11918));
    LocalMux I__2866 (
            .O(N__11927),
            .I(N__11913));
    LocalMux I__2865 (
            .O(N__11924),
            .I(N__11913));
    Span4Mux_h I__2864 (
            .O(N__11921),
            .I(N__11908));
    Span4Mux_v I__2863 (
            .O(N__11918),
            .I(N__11908));
    Span12Mux_v I__2862 (
            .O(N__11913),
            .I(N__11905));
    Sp12to4 I__2861 (
            .O(N__11908),
            .I(N__11902));
    Span12Mux_h I__2860 (
            .O(N__11905),
            .I(N__11899));
    Odrv12 I__2859 (
            .O(N__11902),
            .I(DRA_c_8));
    Odrv12 I__2858 (
            .O(N__11899),
            .I(DRA_c_8));
    InMux I__2857 (
            .O(N__11894),
            .I(N__11890));
    InMux I__2856 (
            .O(N__11893),
            .I(N__11887));
    LocalMux I__2855 (
            .O(N__11890),
            .I(N__11880));
    LocalMux I__2854 (
            .O(N__11887),
            .I(N__11880));
    InMux I__2853 (
            .O(N__11886),
            .I(N__11877));
    InMux I__2852 (
            .O(N__11885),
            .I(N__11874));
    Span4Mux_h I__2851 (
            .O(N__11880),
            .I(N__11867));
    LocalMux I__2850 (
            .O(N__11877),
            .I(N__11867));
    LocalMux I__2849 (
            .O(N__11874),
            .I(N__11867));
    Span4Mux_v I__2848 (
            .O(N__11867),
            .I(N__11864));
    Sp12to4 I__2847 (
            .O(N__11864),
            .I(N__11861));
    Span12Mux_h I__2846 (
            .O(N__11861),
            .I(N__11858));
    Odrv12 I__2845 (
            .O(N__11858),
            .I(DRA_c_7));
    InMux I__2844 (
            .O(N__11855),
            .I(N__11852));
    LocalMux I__2843 (
            .O(N__11852),
            .I(N__11849));
    Odrv4 I__2842 (
            .O(N__11849),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__2841 (
            .O(N__11846),
            .I(N__11842));
    InMux I__2840 (
            .O(N__11845),
            .I(N__11838));
    LocalMux I__2839 (
            .O(N__11842),
            .I(N__11835));
    InMux I__2838 (
            .O(N__11841),
            .I(N__11832));
    LocalMux I__2837 (
            .O(N__11838),
            .I(N__11829));
    Span4Mux_v I__2836 (
            .O(N__11835),
            .I(N__11825));
    LocalMux I__2835 (
            .O(N__11832),
            .I(N__11822));
    Span4Mux_h I__2834 (
            .O(N__11829),
            .I(N__11819));
    InMux I__2833 (
            .O(N__11828),
            .I(N__11816));
    Span4Mux_h I__2832 (
            .O(N__11825),
            .I(N__11811));
    Span4Mux_v I__2831 (
            .O(N__11822),
            .I(N__11811));
    Sp12to4 I__2830 (
            .O(N__11819),
            .I(N__11806));
    LocalMux I__2829 (
            .O(N__11816),
            .I(N__11806));
    Span4Mux_v I__2828 (
            .O(N__11811),
            .I(N__11803));
    Span12Mux_v I__2827 (
            .O(N__11806),
            .I(N__11798));
    Sp12to4 I__2826 (
            .O(N__11803),
            .I(N__11798));
    Span12Mux_h I__2825 (
            .O(N__11798),
            .I(N__11795));
    Span12Mux_v I__2824 (
            .O(N__11795),
            .I(N__11792));
    Odrv12 I__2823 (
            .O(N__11792),
            .I(DRA_c_9));
    CascadeMux I__2822 (
            .O(N__11789),
            .I(N__11786));
    InMux I__2821 (
            .O(N__11786),
            .I(N__11783));
    LocalMux I__2820 (
            .O(N__11783),
            .I(N__11772));
    CascadeMux I__2819 (
            .O(N__11782),
            .I(N__11769));
    InMux I__2818 (
            .O(N__11781),
            .I(N__11766));
    InMux I__2817 (
            .O(N__11780),
            .I(N__11761));
    InMux I__2816 (
            .O(N__11779),
            .I(N__11761));
    InMux I__2815 (
            .O(N__11778),
            .I(N__11756));
    InMux I__2814 (
            .O(N__11777),
            .I(N__11756));
    InMux I__2813 (
            .O(N__11776),
            .I(N__11753));
    InMux I__2812 (
            .O(N__11775),
            .I(N__11743));
    Span4Mux_v I__2811 (
            .O(N__11772),
            .I(N__11740));
    InMux I__2810 (
            .O(N__11769),
            .I(N__11737));
    LocalMux I__2809 (
            .O(N__11766),
            .I(N__11728));
    LocalMux I__2808 (
            .O(N__11761),
            .I(N__11728));
    LocalMux I__2807 (
            .O(N__11756),
            .I(N__11728));
    LocalMux I__2806 (
            .O(N__11753),
            .I(N__11728));
    InMux I__2805 (
            .O(N__11752),
            .I(N__11723));
    InMux I__2804 (
            .O(N__11751),
            .I(N__11723));
    InMux I__2803 (
            .O(N__11750),
            .I(N__11720));
    InMux I__2802 (
            .O(N__11749),
            .I(N__11717));
    InMux I__2801 (
            .O(N__11748),
            .I(N__11714));
    InMux I__2800 (
            .O(N__11747),
            .I(N__11711));
    InMux I__2799 (
            .O(N__11746),
            .I(N__11707));
    LocalMux I__2798 (
            .O(N__11743),
            .I(N__11702));
    Span4Mux_v I__2797 (
            .O(N__11740),
            .I(N__11695));
    LocalMux I__2796 (
            .O(N__11737),
            .I(N__11695));
    Span4Mux_v I__2795 (
            .O(N__11728),
            .I(N__11682));
    LocalMux I__2794 (
            .O(N__11723),
            .I(N__11682));
    LocalMux I__2793 (
            .O(N__11720),
            .I(N__11682));
    LocalMux I__2792 (
            .O(N__11717),
            .I(N__11682));
    LocalMux I__2791 (
            .O(N__11714),
            .I(N__11682));
    LocalMux I__2790 (
            .O(N__11711),
            .I(N__11682));
    CascadeMux I__2789 (
            .O(N__11710),
            .I(N__11679));
    LocalMux I__2788 (
            .O(N__11707),
            .I(N__11676));
    InMux I__2787 (
            .O(N__11706),
            .I(N__11671));
    InMux I__2786 (
            .O(N__11705),
            .I(N__11671));
    Span4Mux_v I__2785 (
            .O(N__11702),
            .I(N__11668));
    InMux I__2784 (
            .O(N__11701),
            .I(N__11665));
    InMux I__2783 (
            .O(N__11700),
            .I(N__11662));
    Span4Mux_h I__2782 (
            .O(N__11695),
            .I(N__11657));
    Span4Mux_v I__2781 (
            .O(N__11682),
            .I(N__11657));
    InMux I__2780 (
            .O(N__11679),
            .I(N__11654));
    Sp12to4 I__2779 (
            .O(N__11676),
            .I(N__11651));
    LocalMux I__2778 (
            .O(N__11671),
            .I(N__11642));
    Sp12to4 I__2777 (
            .O(N__11668),
            .I(N__11642));
    LocalMux I__2776 (
            .O(N__11665),
            .I(N__11642));
    LocalMux I__2775 (
            .O(N__11662),
            .I(N__11642));
    Sp12to4 I__2774 (
            .O(N__11657),
            .I(N__11637));
    LocalMux I__2773 (
            .O(N__11654),
            .I(N__11637));
    Span12Mux_v I__2772 (
            .O(N__11651),
            .I(N__11634));
    Span12Mux_h I__2771 (
            .O(N__11642),
            .I(N__11631));
    Span12Mux_h I__2770 (
            .O(N__11637),
            .I(N__11628));
    Span12Mux_h I__2769 (
            .O(N__11634),
            .I(N__11623));
    Span12Mux_v I__2768 (
            .O(N__11631),
            .I(N__11623));
    Span12Mux_v I__2767 (
            .O(N__11628),
            .I(N__11620));
    Odrv12 I__2766 (
            .O(N__11623),
            .I(AGNUS_REV_c));
    Odrv12 I__2765 (
            .O(N__11620),
            .I(AGNUS_REV_c));
    InMux I__2764 (
            .O(N__11615),
            .I(N__11612));
    LocalMux I__2763 (
            .O(N__11612),
            .I(N__11609));
    Span4Mux_v I__2762 (
            .O(N__11609),
            .I(N__11606));
    Odrv4 I__2761 (
            .O(N__11606),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    ClkMux I__2760 (
            .O(N__11603),
            .I(N__11579));
    ClkMux I__2759 (
            .O(N__11602),
            .I(N__11579));
    ClkMux I__2758 (
            .O(N__11601),
            .I(N__11579));
    ClkMux I__2757 (
            .O(N__11600),
            .I(N__11579));
    ClkMux I__2756 (
            .O(N__11599),
            .I(N__11579));
    ClkMux I__2755 (
            .O(N__11598),
            .I(N__11579));
    ClkMux I__2754 (
            .O(N__11597),
            .I(N__11579));
    ClkMux I__2753 (
            .O(N__11596),
            .I(N__11579));
    GlobalMux I__2752 (
            .O(N__11579),
            .I(N__11576));
    gio2CtrlBuf I__2751 (
            .O(N__11576),
            .I(C3_c_g));
    CEMux I__2750 (
            .O(N__11573),
            .I(N__11528));
    CEMux I__2749 (
            .O(N__11572),
            .I(N__11528));
    CEMux I__2748 (
            .O(N__11571),
            .I(N__11528));
    CEMux I__2747 (
            .O(N__11570),
            .I(N__11528));
    CEMux I__2746 (
            .O(N__11569),
            .I(N__11528));
    CEMux I__2745 (
            .O(N__11568),
            .I(N__11528));
    CEMux I__2744 (
            .O(N__11567),
            .I(N__11528));
    CEMux I__2743 (
            .O(N__11566),
            .I(N__11528));
    CEMux I__2742 (
            .O(N__11565),
            .I(N__11528));
    CEMux I__2741 (
            .O(N__11564),
            .I(N__11528));
    CEMux I__2740 (
            .O(N__11563),
            .I(N__11528));
    CEMux I__2739 (
            .O(N__11562),
            .I(N__11528));
    CEMux I__2738 (
            .O(N__11561),
            .I(N__11528));
    CEMux I__2737 (
            .O(N__11560),
            .I(N__11528));
    CEMux I__2736 (
            .O(N__11559),
            .I(N__11528));
    GlobalMux I__2735 (
            .O(N__11528),
            .I(N__11525));
    gio2CtrlBuf I__2734 (
            .O(N__11525),
            .I(DBRn_c_i_0_g));
    InMux I__2733 (
            .O(N__11522),
            .I(N__11518));
    InMux I__2732 (
            .O(N__11521),
            .I(N__11515));
    LocalMux I__2731 (
            .O(N__11518),
            .I(N__11512));
    LocalMux I__2730 (
            .O(N__11515),
            .I(N__11509));
    Span4Mux_v I__2729 (
            .O(N__11512),
            .I(N__11504));
    Span4Mux_v I__2728 (
            .O(N__11509),
            .I(N__11504));
    Sp12to4 I__2727 (
            .O(N__11504),
            .I(N__11501));
    Odrv12 I__2726 (
            .O(N__11501),
            .I(RAS0n_c));
    InMux I__2725 (
            .O(N__11498),
            .I(N__11495));
    LocalMux I__2724 (
            .O(N__11495),
            .I(N__11492));
    Span12Mux_h I__2723 (
            .O(N__11492),
            .I(N__11489));
    Odrv12 I__2722 (
            .O(N__11489),
            .I(RAS1n_c));
    InMux I__2721 (
            .O(N__11486),
            .I(N__11483));
    LocalMux I__2720 (
            .O(N__11483),
            .I(N__11480));
    Span12Mux_h I__2719 (
            .O(N__11480),
            .I(N__11477));
    Odrv12 I__2718 (
            .O(N__11477),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ));
    InMux I__2717 (
            .O(N__11474),
            .I(N__11471));
    LocalMux I__2716 (
            .O(N__11471),
            .I(N__11432));
    ClkMux I__2715 (
            .O(N__11470),
            .I(N__11330));
    ClkMux I__2714 (
            .O(N__11469),
            .I(N__11330));
    ClkMux I__2713 (
            .O(N__11468),
            .I(N__11330));
    ClkMux I__2712 (
            .O(N__11467),
            .I(N__11330));
    ClkMux I__2711 (
            .O(N__11466),
            .I(N__11330));
    ClkMux I__2710 (
            .O(N__11465),
            .I(N__11330));
    ClkMux I__2709 (
            .O(N__11464),
            .I(N__11330));
    ClkMux I__2708 (
            .O(N__11463),
            .I(N__11330));
    ClkMux I__2707 (
            .O(N__11462),
            .I(N__11330));
    ClkMux I__2706 (
            .O(N__11461),
            .I(N__11330));
    ClkMux I__2705 (
            .O(N__11460),
            .I(N__11330));
    ClkMux I__2704 (
            .O(N__11459),
            .I(N__11330));
    ClkMux I__2703 (
            .O(N__11458),
            .I(N__11330));
    ClkMux I__2702 (
            .O(N__11457),
            .I(N__11330));
    ClkMux I__2701 (
            .O(N__11456),
            .I(N__11330));
    ClkMux I__2700 (
            .O(N__11455),
            .I(N__11330));
    ClkMux I__2699 (
            .O(N__11454),
            .I(N__11330));
    ClkMux I__2698 (
            .O(N__11453),
            .I(N__11330));
    ClkMux I__2697 (
            .O(N__11452),
            .I(N__11330));
    ClkMux I__2696 (
            .O(N__11451),
            .I(N__11330));
    ClkMux I__2695 (
            .O(N__11450),
            .I(N__11330));
    ClkMux I__2694 (
            .O(N__11449),
            .I(N__11330));
    ClkMux I__2693 (
            .O(N__11448),
            .I(N__11330));
    ClkMux I__2692 (
            .O(N__11447),
            .I(N__11330));
    ClkMux I__2691 (
            .O(N__11446),
            .I(N__11330));
    ClkMux I__2690 (
            .O(N__11445),
            .I(N__11330));
    ClkMux I__2689 (
            .O(N__11444),
            .I(N__11330));
    ClkMux I__2688 (
            .O(N__11443),
            .I(N__11330));
    ClkMux I__2687 (
            .O(N__11442),
            .I(N__11330));
    ClkMux I__2686 (
            .O(N__11441),
            .I(N__11330));
    ClkMux I__2685 (
            .O(N__11440),
            .I(N__11330));
    ClkMux I__2684 (
            .O(N__11439),
            .I(N__11330));
    ClkMux I__2683 (
            .O(N__11438),
            .I(N__11330));
    ClkMux I__2682 (
            .O(N__11437),
            .I(N__11330));
    ClkMux I__2681 (
            .O(N__11436),
            .I(N__11330));
    ClkMux I__2680 (
            .O(N__11435),
            .I(N__11330));
    Glb2LocalMux I__2679 (
            .O(N__11432),
            .I(N__11330));
    ClkMux I__2678 (
            .O(N__11431),
            .I(N__11330));
    ClkMux I__2677 (
            .O(N__11430),
            .I(N__11330));
    ClkMux I__2676 (
            .O(N__11429),
            .I(N__11330));
    ClkMux I__2675 (
            .O(N__11428),
            .I(N__11330));
    ClkMux I__2674 (
            .O(N__11427),
            .I(N__11330));
    ClkMux I__2673 (
            .O(N__11426),
            .I(N__11330));
    ClkMux I__2672 (
            .O(N__11425),
            .I(N__11330));
    ClkMux I__2671 (
            .O(N__11424),
            .I(N__11330));
    ClkMux I__2670 (
            .O(N__11423),
            .I(N__11330));
    GlobalMux I__2669 (
            .O(N__11330),
            .I(CLK80_PLL));
    InMux I__2668 (
            .O(N__11327),
            .I(N__11320));
    InMux I__2667 (
            .O(N__11326),
            .I(N__11317));
    InMux I__2666 (
            .O(N__11325),
            .I(N__11314));
    InMux I__2665 (
            .O(N__11324),
            .I(N__11311));
    InMux I__2664 (
            .O(N__11323),
            .I(N__11308));
    LocalMux I__2663 (
            .O(N__11320),
            .I(N__11303));
    LocalMux I__2662 (
            .O(N__11317),
            .I(N__11272));
    LocalMux I__2661 (
            .O(N__11314),
            .I(N__11269));
    LocalMux I__2660 (
            .O(N__11311),
            .I(N__11251));
    LocalMux I__2659 (
            .O(N__11308),
            .I(N__11247));
    SRMux I__2658 (
            .O(N__11307),
            .I(N__11135));
    SRMux I__2657 (
            .O(N__11306),
            .I(N__11135));
    Glb2LocalMux I__2656 (
            .O(N__11303),
            .I(N__11135));
    SRMux I__2655 (
            .O(N__11302),
            .I(N__11135));
    SRMux I__2654 (
            .O(N__11301),
            .I(N__11135));
    SRMux I__2653 (
            .O(N__11300),
            .I(N__11135));
    SRMux I__2652 (
            .O(N__11299),
            .I(N__11135));
    SRMux I__2651 (
            .O(N__11298),
            .I(N__11135));
    SRMux I__2650 (
            .O(N__11297),
            .I(N__11135));
    SRMux I__2649 (
            .O(N__11296),
            .I(N__11135));
    SRMux I__2648 (
            .O(N__11295),
            .I(N__11135));
    SRMux I__2647 (
            .O(N__11294),
            .I(N__11135));
    SRMux I__2646 (
            .O(N__11293),
            .I(N__11135));
    SRMux I__2645 (
            .O(N__11292),
            .I(N__11135));
    SRMux I__2644 (
            .O(N__11291),
            .I(N__11135));
    SRMux I__2643 (
            .O(N__11290),
            .I(N__11135));
    SRMux I__2642 (
            .O(N__11289),
            .I(N__11135));
    SRMux I__2641 (
            .O(N__11288),
            .I(N__11135));
    SRMux I__2640 (
            .O(N__11287),
            .I(N__11135));
    SRMux I__2639 (
            .O(N__11286),
            .I(N__11135));
    SRMux I__2638 (
            .O(N__11285),
            .I(N__11135));
    SRMux I__2637 (
            .O(N__11284),
            .I(N__11135));
    SRMux I__2636 (
            .O(N__11283),
            .I(N__11135));
    SRMux I__2635 (
            .O(N__11282),
            .I(N__11135));
    SRMux I__2634 (
            .O(N__11281),
            .I(N__11135));
    SRMux I__2633 (
            .O(N__11280),
            .I(N__11135));
    SRMux I__2632 (
            .O(N__11279),
            .I(N__11135));
    SRMux I__2631 (
            .O(N__11278),
            .I(N__11135));
    SRMux I__2630 (
            .O(N__11277),
            .I(N__11135));
    SRMux I__2629 (
            .O(N__11276),
            .I(N__11135));
    SRMux I__2628 (
            .O(N__11275),
            .I(N__11135));
    Glb2LocalMux I__2627 (
            .O(N__11272),
            .I(N__11135));
    Glb2LocalMux I__2626 (
            .O(N__11269),
            .I(N__11135));
    SRMux I__2625 (
            .O(N__11268),
            .I(N__11135));
    SRMux I__2624 (
            .O(N__11267),
            .I(N__11135));
    SRMux I__2623 (
            .O(N__11266),
            .I(N__11135));
    SRMux I__2622 (
            .O(N__11265),
            .I(N__11135));
    SRMux I__2621 (
            .O(N__11264),
            .I(N__11135));
    SRMux I__2620 (
            .O(N__11263),
            .I(N__11135));
    SRMux I__2619 (
            .O(N__11262),
            .I(N__11135));
    SRMux I__2618 (
            .O(N__11261),
            .I(N__11135));
    SRMux I__2617 (
            .O(N__11260),
            .I(N__11135));
    SRMux I__2616 (
            .O(N__11259),
            .I(N__11135));
    SRMux I__2615 (
            .O(N__11258),
            .I(N__11135));
    SRMux I__2614 (
            .O(N__11257),
            .I(N__11135));
    SRMux I__2613 (
            .O(N__11256),
            .I(N__11135));
    SRMux I__2612 (
            .O(N__11255),
            .I(N__11135));
    SRMux I__2611 (
            .O(N__11254),
            .I(N__11135));
    Glb2LocalMux I__2610 (
            .O(N__11251),
            .I(N__11135));
    SRMux I__2609 (
            .O(N__11250),
            .I(N__11135));
    Glb2LocalMux I__2608 (
            .O(N__11247),
            .I(N__11135));
    SRMux I__2607 (
            .O(N__11246),
            .I(N__11135));
    SRMux I__2606 (
            .O(N__11245),
            .I(N__11135));
    SRMux I__2605 (
            .O(N__11244),
            .I(N__11135));
    GlobalMux I__2604 (
            .O(N__11135),
            .I(N__11132));
    gio2CtrlBuf I__2603 (
            .O(N__11132),
            .I(RESETn_c_i_g));
    InMux I__2602 (
            .O(N__11129),
            .I(N__11126));
    LocalMux I__2601 (
            .O(N__11126),
            .I(N__11123));
    Sp12to4 I__2600 (
            .O(N__11123),
            .I(N__11119));
    InMux I__2599 (
            .O(N__11122),
            .I(N__11116));
    Span12Mux_v I__2598 (
            .O(N__11119),
            .I(N__11113));
    LocalMux I__2597 (
            .O(N__11116),
            .I(N__11110));
    Span12Mux_h I__2596 (
            .O(N__11113),
            .I(N__11105));
    Span12Mux_v I__2595 (
            .O(N__11110),
            .I(N__11102));
    InMux I__2594 (
            .O(N__11109),
            .I(N__11099));
    InMux I__2593 (
            .O(N__11108),
            .I(N__11096));
    Odrv12 I__2592 (
            .O(N__11105),
            .I(REG_CYCLEm));
    Odrv12 I__2591 (
            .O(N__11102),
            .I(REG_CYCLEm));
    LocalMux I__2590 (
            .O(N__11099),
            .I(REG_CYCLEm));
    LocalMux I__2589 (
            .O(N__11096),
            .I(REG_CYCLEm));
    InMux I__2588 (
            .O(N__11087),
            .I(N__11084));
    LocalMux I__2587 (
            .O(N__11084),
            .I(N__11081));
    Span4Mux_v I__2586 (
            .O(N__11081),
            .I(N__11077));
    CascadeMux I__2585 (
            .O(N__11080),
            .I(N__11073));
    Span4Mux_h I__2584 (
            .O(N__11077),
            .I(N__11067));
    InMux I__2583 (
            .O(N__11076),
            .I(N__11057));
    InMux I__2582 (
            .O(N__11073),
            .I(N__11052));
    InMux I__2581 (
            .O(N__11072),
            .I(N__11052));
    InMux I__2580 (
            .O(N__11071),
            .I(N__11047));
    InMux I__2579 (
            .O(N__11070),
            .I(N__11047));
    Span4Mux_h I__2578 (
            .O(N__11067),
            .I(N__11040));
    InMux I__2577 (
            .O(N__11066),
            .I(N__11031));
    InMux I__2576 (
            .O(N__11065),
            .I(N__11031));
    InMux I__2575 (
            .O(N__11064),
            .I(N__11031));
    InMux I__2574 (
            .O(N__11063),
            .I(N__11031));
    CascadeMux I__2573 (
            .O(N__11062),
            .I(N__11026));
    CascadeMux I__2572 (
            .O(N__11061),
            .I(N__11023));
    InMux I__2571 (
            .O(N__11060),
            .I(N__11019));
    LocalMux I__2570 (
            .O(N__11057),
            .I(N__11016));
    LocalMux I__2569 (
            .O(N__11052),
            .I(N__11013));
    LocalMux I__2568 (
            .O(N__11047),
            .I(N__11010));
    InMux I__2567 (
            .O(N__11046),
            .I(N__11005));
    InMux I__2566 (
            .O(N__11045),
            .I(N__11005));
    CascadeMux I__2565 (
            .O(N__11044),
            .I(N__11001));
    InMux I__2564 (
            .O(N__11043),
            .I(N__10995));
    Span4Mux_v I__2563 (
            .O(N__11040),
            .I(N__10987));
    LocalMux I__2562 (
            .O(N__11031),
            .I(N__10987));
    InMux I__2561 (
            .O(N__11030),
            .I(N__10984));
    InMux I__2560 (
            .O(N__11029),
            .I(N__10981));
    InMux I__2559 (
            .O(N__11026),
            .I(N__10976));
    InMux I__2558 (
            .O(N__11023),
            .I(N__10976));
    InMux I__2557 (
            .O(N__11022),
            .I(N__10973));
    LocalMux I__2556 (
            .O(N__11019),
            .I(N__10970));
    Span4Mux_v I__2555 (
            .O(N__11016),
            .I(N__10961));
    Span4Mux_h I__2554 (
            .O(N__11013),
            .I(N__10961));
    Span4Mux_v I__2553 (
            .O(N__11010),
            .I(N__10961));
    LocalMux I__2552 (
            .O(N__11005),
            .I(N__10961));
    InMux I__2551 (
            .O(N__11004),
            .I(N__10958));
    InMux I__2550 (
            .O(N__11001),
            .I(N__10955));
    InMux I__2549 (
            .O(N__11000),
            .I(N__10948));
    InMux I__2548 (
            .O(N__10999),
            .I(N__10948));
    InMux I__2547 (
            .O(N__10998),
            .I(N__10948));
    LocalMux I__2546 (
            .O(N__10995),
            .I(N__10945));
    InMux I__2545 (
            .O(N__10994),
            .I(N__10940));
    InMux I__2544 (
            .O(N__10993),
            .I(N__10940));
    InMux I__2543 (
            .O(N__10992),
            .I(N__10934));
    Span4Mux_h I__2542 (
            .O(N__10987),
            .I(N__10929));
    LocalMux I__2541 (
            .O(N__10984),
            .I(N__10929));
    LocalMux I__2540 (
            .O(N__10981),
            .I(N__10916));
    LocalMux I__2539 (
            .O(N__10976),
            .I(N__10916));
    LocalMux I__2538 (
            .O(N__10973),
            .I(N__10916));
    Span4Mux_h I__2537 (
            .O(N__10970),
            .I(N__10916));
    Span4Mux_h I__2536 (
            .O(N__10961),
            .I(N__10916));
    LocalMux I__2535 (
            .O(N__10958),
            .I(N__10916));
    LocalMux I__2534 (
            .O(N__10955),
            .I(N__10908));
    LocalMux I__2533 (
            .O(N__10948),
            .I(N__10908));
    Span4Mux_v I__2532 (
            .O(N__10945),
            .I(N__10908));
    LocalMux I__2531 (
            .O(N__10940),
            .I(N__10905));
    InMux I__2530 (
            .O(N__10939),
            .I(N__10898));
    InMux I__2529 (
            .O(N__10938),
            .I(N__10898));
    InMux I__2528 (
            .O(N__10937),
            .I(N__10898));
    LocalMux I__2527 (
            .O(N__10934),
            .I(N__10895));
    Span4Mux_v I__2526 (
            .O(N__10929),
            .I(N__10890));
    Span4Mux_v I__2525 (
            .O(N__10916),
            .I(N__10890));
    InMux I__2524 (
            .O(N__10915),
            .I(N__10887));
    Span4Mux_h I__2523 (
            .O(N__10908),
            .I(N__10880));
    Span4Mux_v I__2522 (
            .O(N__10905),
            .I(N__10880));
    LocalMux I__2521 (
            .O(N__10898),
            .I(N__10880));
    Odrv4 I__2520 (
            .O(N__10895),
            .I(\U712_CHIP_RAM.CPU_CYCLEm ));
    Odrv4 I__2519 (
            .O(N__10890),
            .I(\U712_CHIP_RAM.CPU_CYCLEm ));
    LocalMux I__2518 (
            .O(N__10887),
            .I(\U712_CHIP_RAM.CPU_CYCLEm ));
    Odrv4 I__2517 (
            .O(N__10880),
            .I(\U712_CHIP_RAM.CPU_CYCLEm ));
    IoInMux I__2516 (
            .O(N__10871),
            .I(N__10868));
    LocalMux I__2515 (
            .O(N__10868),
            .I(N__10865));
    Span4Mux_s3_v I__2514 (
            .O(N__10865),
            .I(N__10862));
    Span4Mux_v I__2513 (
            .O(N__10862),
            .I(N__10859));
    Odrv4 I__2512 (
            .O(N__10859),
            .I(N_338_mux));
    InMux I__2511 (
            .O(N__10856),
            .I(N__10853));
    LocalMux I__2510 (
            .O(N__10853),
            .I(N__10849));
    InMux I__2509 (
            .O(N__10852),
            .I(N__10846));
    Span4Mux_h I__2508 (
            .O(N__10849),
            .I(N__10840));
    LocalMux I__2507 (
            .O(N__10846),
            .I(N__10840));
    InMux I__2506 (
            .O(N__10845),
            .I(N__10837));
    Span4Mux_v I__2505 (
            .O(N__10840),
            .I(N__10831));
    LocalMux I__2504 (
            .O(N__10837),
            .I(N__10831));
    CascadeMux I__2503 (
            .O(N__10836),
            .I(N__10827));
    Sp12to4 I__2502 (
            .O(N__10831),
            .I(N__10824));
    InMux I__2501 (
            .O(N__10830),
            .I(N__10819));
    InMux I__2500 (
            .O(N__10827),
            .I(N__10819));
    Span12Mux_v I__2499 (
            .O(N__10824),
            .I(N__10816));
    LocalMux I__2498 (
            .O(N__10819),
            .I(N__10813));
    Span12Mux_h I__2497 (
            .O(N__10816),
            .I(N__10810));
    Span12Mux_v I__2496 (
            .O(N__10813),
            .I(N__10807));
    Odrv12 I__2495 (
            .O(N__10810),
            .I(CASLn_c));
    Odrv12 I__2494 (
            .O(N__10807),
            .I(CASLn_c));
    InMux I__2493 (
            .O(N__10802),
            .I(N__10798));
    InMux I__2492 (
            .O(N__10801),
            .I(N__10795));
    LocalMux I__2491 (
            .O(N__10798),
            .I(N__10789));
    LocalMux I__2490 (
            .O(N__10795),
            .I(N__10786));
    InMux I__2489 (
            .O(N__10794),
            .I(N__10781));
    InMux I__2488 (
            .O(N__10793),
            .I(N__10781));
    InMux I__2487 (
            .O(N__10792),
            .I(N__10778));
    Span4Mux_v I__2486 (
            .O(N__10789),
            .I(N__10775));
    Span4Mux_v I__2485 (
            .O(N__10786),
            .I(N__10772));
    LocalMux I__2484 (
            .O(N__10781),
            .I(N__10769));
    LocalMux I__2483 (
            .O(N__10778),
            .I(N__10766));
    Sp12to4 I__2482 (
            .O(N__10775),
            .I(N__10763));
    Span4Mux_h I__2481 (
            .O(N__10772),
            .I(N__10758));
    Span4Mux_v I__2480 (
            .O(N__10769),
            .I(N__10758));
    Span4Mux_v I__2479 (
            .O(N__10766),
            .I(N__10755));
    Span12Mux_h I__2478 (
            .O(N__10763),
            .I(N__10748));
    Sp12to4 I__2477 (
            .O(N__10758),
            .I(N__10748));
    Sp12to4 I__2476 (
            .O(N__10755),
            .I(N__10748));
    Span12Mux_h I__2475 (
            .O(N__10748),
            .I(N__10745));
    Odrv12 I__2474 (
            .O(N__10745),
            .I(RnW_c));
    CascadeMux I__2473 (
            .O(N__10742),
            .I(N__10739));
    InMux I__2472 (
            .O(N__10739),
            .I(N__10736));
    LocalMux I__2471 (
            .O(N__10736),
            .I(N__10732));
    InMux I__2470 (
            .O(N__10735),
            .I(N__10729));
    Sp12to4 I__2469 (
            .O(N__10732),
            .I(N__10724));
    LocalMux I__2468 (
            .O(N__10729),
            .I(N__10724));
    Span12Mux_h I__2467 (
            .O(N__10724),
            .I(N__10720));
    InMux I__2466 (
            .O(N__10723),
            .I(N__10717));
    Odrv12 I__2465 (
            .O(N__10720),
            .I(\U712_CHIP_RAM.DMA_WRITE_CYCLEZ0 ));
    LocalMux I__2464 (
            .O(N__10717),
            .I(\U712_CHIP_RAM.DMA_WRITE_CYCLEZ0 ));
    InMux I__2463 (
            .O(N__10712),
            .I(N__10709));
    LocalMux I__2462 (
            .O(N__10709),
            .I(N__10704));
    InMux I__2461 (
            .O(N__10708),
            .I(N__10701));
    InMux I__2460 (
            .O(N__10707),
            .I(N__10698));
    Span4Mux_v I__2459 (
            .O(N__10704),
            .I(N__10693));
    LocalMux I__2458 (
            .O(N__10701),
            .I(N__10693));
    LocalMux I__2457 (
            .O(N__10698),
            .I(N__10690));
    Span4Mux_v I__2456 (
            .O(N__10693),
            .I(N__10685));
    Span4Mux_h I__2455 (
            .O(N__10690),
            .I(N__10685));
    Span4Mux_h I__2454 (
            .O(N__10685),
            .I(N__10680));
    InMux I__2453 (
            .O(N__10684),
            .I(N__10675));
    InMux I__2452 (
            .O(N__10683),
            .I(N__10675));
    Span4Mux_h I__2451 (
            .O(N__10680),
            .I(N__10670));
    LocalMux I__2450 (
            .O(N__10675),
            .I(N__10670));
    Span4Mux_h I__2449 (
            .O(N__10670),
            .I(N__10667));
    Span4Mux_v I__2448 (
            .O(N__10667),
            .I(N__10664));
    Odrv4 I__2447 (
            .O(N__10664),
            .I(CASUn_c));
    IoInMux I__2446 (
            .O(N__10661),
            .I(N__10658));
    LocalMux I__2445 (
            .O(N__10658),
            .I(N__10655));
    IoSpan4Mux I__2444 (
            .O(N__10655),
            .I(N__10652));
    Span4Mux_s3_h I__2443 (
            .O(N__10652),
            .I(N__10649));
    Odrv4 I__2442 (
            .O(N__10649),
            .I(N_328_mux));
    InMux I__2441 (
            .O(N__10646),
            .I(N__10643));
    LocalMux I__2440 (
            .O(N__10643),
            .I(N__10639));
    InMux I__2439 (
            .O(N__10642),
            .I(N__10636));
    Span4Mux_h I__2438 (
            .O(N__10639),
            .I(N__10631));
    LocalMux I__2437 (
            .O(N__10636),
            .I(N__10631));
    Span4Mux_v I__2436 (
            .O(N__10631),
            .I(N__10626));
    InMux I__2435 (
            .O(N__10630),
            .I(N__10623));
    InMux I__2434 (
            .O(N__10629),
            .I(N__10620));
    Span4Mux_v I__2433 (
            .O(N__10626),
            .I(N__10617));
    LocalMux I__2432 (
            .O(N__10623),
            .I(N__10612));
    LocalMux I__2431 (
            .O(N__10620),
            .I(N__10612));
    Sp12to4 I__2430 (
            .O(N__10617),
            .I(N__10607));
    Span12Mux_v I__2429 (
            .O(N__10612),
            .I(N__10607));
    Span12Mux_h I__2428 (
            .O(N__10607),
            .I(N__10604));
    Odrv12 I__2427 (
            .O(N__10604),
            .I(DRA_c_6));
    InMux I__2426 (
            .O(N__10601),
            .I(N__10598));
    LocalMux I__2425 (
            .O(N__10598),
            .I(N__10595));
    Span4Mux_h I__2424 (
            .O(N__10595),
            .I(N__10592));
    Odrv4 I__2423 (
            .O(N__10592),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__2422 (
            .O(N__10589),
            .I(N__10586));
    LocalMux I__2421 (
            .O(N__10586),
            .I(N__10583));
    Odrv4 I__2420 (
            .O(N__10583),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__2419 (
            .O(N__10580),
            .I(N__10576));
    InMux I__2418 (
            .O(N__10579),
            .I(N__10573));
    LocalMux I__2417 (
            .O(N__10576),
            .I(N__10566));
    LocalMux I__2416 (
            .O(N__10573),
            .I(N__10566));
    InMux I__2415 (
            .O(N__10572),
            .I(N__10563));
    InMux I__2414 (
            .O(N__10571),
            .I(N__10560));
    Span4Mux_v I__2413 (
            .O(N__10566),
            .I(N__10557));
    LocalMux I__2412 (
            .O(N__10563),
            .I(N__10552));
    LocalMux I__2411 (
            .O(N__10560),
            .I(N__10552));
    Span4Mux_v I__2410 (
            .O(N__10557),
            .I(N__10549));
    Span12Mux_v I__2409 (
            .O(N__10552),
            .I(N__10544));
    Sp12to4 I__2408 (
            .O(N__10549),
            .I(N__10544));
    Span12Mux_h I__2407 (
            .O(N__10544),
            .I(N__10541));
    Odrv12 I__2406 (
            .O(N__10541),
            .I(DRA_c_3));
    InMux I__2405 (
            .O(N__10538),
            .I(N__10535));
    LocalMux I__2404 (
            .O(N__10535),
            .I(N__10532));
    Odrv4 I__2403 (
            .O(N__10532),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__2402 (
            .O(N__10529),
            .I(N__10524));
    InMux I__2401 (
            .O(N__10528),
            .I(N__10521));
    InMux I__2400 (
            .O(N__10527),
            .I(N__10518));
    LocalMux I__2399 (
            .O(N__10524),
            .I(N__10510));
    LocalMux I__2398 (
            .O(N__10521),
            .I(N__10510));
    LocalMux I__2397 (
            .O(N__10518),
            .I(N__10510));
    InMux I__2396 (
            .O(N__10517),
            .I(N__10507));
    Span4Mux_v I__2395 (
            .O(N__10510),
            .I(N__10504));
    LocalMux I__2394 (
            .O(N__10507),
            .I(N__10501));
    Sp12to4 I__2393 (
            .O(N__10504),
            .I(N__10498));
    Span4Mux_h I__2392 (
            .O(N__10501),
            .I(N__10495));
    Span12Mux_h I__2391 (
            .O(N__10498),
            .I(N__10492));
    Sp12to4 I__2390 (
            .O(N__10495),
            .I(N__10489));
    Span12Mux_v I__2389 (
            .O(N__10492),
            .I(N__10486));
    Span12Mux_v I__2388 (
            .O(N__10489),
            .I(N__10483));
    Odrv12 I__2387 (
            .O(N__10486),
            .I(DRA_c_2));
    Odrv12 I__2386 (
            .O(N__10483),
            .I(DRA_c_2));
    InMux I__2385 (
            .O(N__10478),
            .I(N__10475));
    LocalMux I__2384 (
            .O(N__10475),
            .I(N__10472));
    Span4Mux_h I__2383 (
            .O(N__10472),
            .I(N__10469));
    Span4Mux_h I__2382 (
            .O(N__10469),
            .I(N__10466));
    Odrv4 I__2381 (
            .O(N__10466),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__2380 (
            .O(N__10463),
            .I(N__10460));
    LocalMux I__2379 (
            .O(N__10460),
            .I(N__10457));
    Span4Mux_h I__2378 (
            .O(N__10457),
            .I(N__10454));
    Odrv4 I__2377 (
            .O(N__10454),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__2376 (
            .O(N__10451),
            .I(N__10447));
    InMux I__2375 (
            .O(N__10450),
            .I(N__10444));
    LocalMux I__2374 (
            .O(N__10447),
            .I(N__10441));
    LocalMux I__2373 (
            .O(N__10444),
            .I(N__10438));
    Sp12to4 I__2372 (
            .O(N__10441),
            .I(N__10435));
    Span12Mux_h I__2371 (
            .O(N__10438),
            .I(N__10432));
    Span12Mux_v I__2370 (
            .O(N__10435),
            .I(N__10429));
    Span12Mux_v I__2369 (
            .O(N__10432),
            .I(N__10426));
    Span12Mux_h I__2368 (
            .O(N__10429),
            .I(N__10423));
    Odrv12 I__2367 (
            .O(N__10426),
            .I(DRA_c_0));
    Odrv12 I__2366 (
            .O(N__10423),
            .I(DRA_c_0));
    InMux I__2365 (
            .O(N__10418),
            .I(N__10414));
    InMux I__2364 (
            .O(N__10417),
            .I(N__10410));
    LocalMux I__2363 (
            .O(N__10414),
            .I(N__10406));
    InMux I__2362 (
            .O(N__10413),
            .I(N__10403));
    LocalMux I__2361 (
            .O(N__10410),
            .I(N__10400));
    InMux I__2360 (
            .O(N__10409),
            .I(N__10397));
    Span4Mux_v I__2359 (
            .O(N__10406),
            .I(N__10390));
    LocalMux I__2358 (
            .O(N__10403),
            .I(N__10390));
    Span4Mux_v I__2357 (
            .O(N__10400),
            .I(N__10390));
    LocalMux I__2356 (
            .O(N__10397),
            .I(N__10387));
    Sp12to4 I__2355 (
            .O(N__10390),
            .I(N__10384));
    Span4Mux_h I__2354 (
            .O(N__10387),
            .I(N__10381));
    Span12Mux_h I__2353 (
            .O(N__10384),
            .I(N__10378));
    Sp12to4 I__2352 (
            .O(N__10381),
            .I(N__10375));
    Span12Mux_v I__2351 (
            .O(N__10378),
            .I(N__10372));
    Span12Mux_v I__2350 (
            .O(N__10375),
            .I(N__10369));
    Odrv12 I__2349 (
            .O(N__10372),
            .I(DRA_c_1));
    Odrv12 I__2348 (
            .O(N__10369),
            .I(DRA_c_1));
    InMux I__2347 (
            .O(N__10364),
            .I(N__10361));
    LocalMux I__2346 (
            .O(N__10361),
            .I(N__10358));
    Span4Mux_h I__2345 (
            .O(N__10358),
            .I(N__10355));
    Odrv4 I__2344 (
            .O(N__10355),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    CascadeMux I__2343 (
            .O(N__10352),
            .I(N__10347));
    InMux I__2342 (
            .O(N__10351),
            .I(N__10344));
    InMux I__2341 (
            .O(N__10350),
            .I(N__10341));
    InMux I__2340 (
            .O(N__10347),
            .I(N__10338));
    LocalMux I__2339 (
            .O(N__10344),
            .I(N__10332));
    LocalMux I__2338 (
            .O(N__10341),
            .I(N__10332));
    LocalMux I__2337 (
            .O(N__10338),
            .I(N__10327));
    InMux I__2336 (
            .O(N__10337),
            .I(N__10324));
    Span4Mux_v I__2335 (
            .O(N__10332),
            .I(N__10321));
    InMux I__2334 (
            .O(N__10331),
            .I(N__10318));
    InMux I__2333 (
            .O(N__10330),
            .I(N__10315));
    Span4Mux_v I__2332 (
            .O(N__10327),
            .I(N__10312));
    LocalMux I__2331 (
            .O(N__10324),
            .I(N__10309));
    Odrv4 I__2330 (
            .O(N__10321),
            .I(\U712_CHIP_RAM.DMA_CYCLEm ));
    LocalMux I__2329 (
            .O(N__10318),
            .I(\U712_CHIP_RAM.DMA_CYCLEm ));
    LocalMux I__2328 (
            .O(N__10315),
            .I(\U712_CHIP_RAM.DMA_CYCLEm ));
    Odrv4 I__2327 (
            .O(N__10312),
            .I(\U712_CHIP_RAM.DMA_CYCLEm ));
    Odrv4 I__2326 (
            .O(N__10309),
            .I(\U712_CHIP_RAM.DMA_CYCLEm ));
    InMux I__2325 (
            .O(N__10298),
            .I(N__10292));
    InMux I__2324 (
            .O(N__10297),
            .I(N__10292));
    LocalMux I__2323 (
            .O(N__10292),
            .I(\U712_CHIP_RAM.N_345 ));
    InMux I__2322 (
            .O(N__10289),
            .I(N__10286));
    LocalMux I__2321 (
            .O(N__10286),
            .I(N__10283));
    Odrv4 I__2320 (
            .O(N__10283),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    InMux I__2319 (
            .O(N__10280),
            .I(N__10277));
    LocalMux I__2318 (
            .O(N__10277),
            .I(\U712_CHIP_RAM.N_346 ));
    IoInMux I__2317 (
            .O(N__10274),
            .I(N__10271));
    LocalMux I__2316 (
            .O(N__10271),
            .I(N__10268));
    IoSpan4Mux I__2315 (
            .O(N__10268),
            .I(N__10265));
    Sp12to4 I__2314 (
            .O(N__10265),
            .I(N__10259));
    CascadeMux I__2313 (
            .O(N__10264),
            .I(N__10256));
    CascadeMux I__2312 (
            .O(N__10263),
            .I(N__10253));
    CascadeMux I__2311 (
            .O(N__10262),
            .I(N__10249));
    Span12Mux_s7_v I__2310 (
            .O(N__10259),
            .I(N__10246));
    InMux I__2309 (
            .O(N__10256),
            .I(N__10243));
    InMux I__2308 (
            .O(N__10253),
            .I(N__10236));
    InMux I__2307 (
            .O(N__10252),
            .I(N__10236));
    InMux I__2306 (
            .O(N__10249),
            .I(N__10236));
    Span12Mux_h I__2305 (
            .O(N__10246),
            .I(N__10232));
    LocalMux I__2304 (
            .O(N__10243),
            .I(N__10227));
    LocalMux I__2303 (
            .O(N__10236),
            .I(N__10227));
    InMux I__2302 (
            .O(N__10235),
            .I(N__10224));
    Odrv12 I__2301 (
            .O(N__10232),
            .I(DBENn_c));
    Odrv4 I__2300 (
            .O(N__10227),
            .I(DBENn_c));
    LocalMux I__2299 (
            .O(N__10224),
            .I(DBENn_c));
    CascadeMux I__2298 (
            .O(N__10217),
            .I(\U712_CHIP_RAM.N_346_cascade_ ));
    IoInMux I__2297 (
            .O(N__10214),
            .I(N__10211));
    LocalMux I__2296 (
            .O(N__10211),
            .I(N__10208));
    IoSpan4Mux I__2295 (
            .O(N__10208),
            .I(N__10205));
    Sp12to4 I__2294 (
            .O(N__10205),
            .I(N__10202));
    Span12Mux_s7_v I__2293 (
            .O(N__10202),
            .I(N__10199));
    Span12Mux_v I__2292 (
            .O(N__10199),
            .I(N__10196));
    Odrv12 I__2291 (
            .O(N__10196),
            .I(CLLBEn_c));
    IoInMux I__2290 (
            .O(N__10193),
            .I(N__10190));
    LocalMux I__2289 (
            .O(N__10190),
            .I(N__10187));
    IoSpan4Mux I__2288 (
            .O(N__10187),
            .I(N__10183));
    InMux I__2287 (
            .O(N__10186),
            .I(N__10180));
    Sp12to4 I__2286 (
            .O(N__10183),
            .I(N__10177));
    LocalMux I__2285 (
            .O(N__10180),
            .I(N__10174));
    Odrv12 I__2284 (
            .O(N__10177),
            .I(LLBEn_c));
    Odrv4 I__2283 (
            .O(N__10174),
            .I(LLBEn_c));
    CascadeMux I__2282 (
            .O(N__10169),
            .I(N__10164));
    InMux I__2281 (
            .O(N__10168),
            .I(N__10161));
    InMux I__2280 (
            .O(N__10167),
            .I(N__10156));
    InMux I__2279 (
            .O(N__10164),
            .I(N__10156));
    LocalMux I__2278 (
            .O(N__10161),
            .I(N__10152));
    LocalMux I__2277 (
            .O(N__10156),
            .I(N__10149));
    InMux I__2276 (
            .O(N__10155),
            .I(N__10146));
    Span4Mux_v I__2275 (
            .O(N__10152),
            .I(N__10143));
    Span4Mux_v I__2274 (
            .O(N__10149),
            .I(N__10140));
    LocalMux I__2273 (
            .O(N__10146),
            .I(N__10137));
    Sp12to4 I__2272 (
            .O(N__10143),
            .I(N__10134));
    Span4Mux_h I__2271 (
            .O(N__10140),
            .I(N__10129));
    Span4Mux_v I__2270 (
            .O(N__10137),
            .I(N__10129));
    Span12Mux_h I__2269 (
            .O(N__10134),
            .I(N__10124));
    Sp12to4 I__2268 (
            .O(N__10129),
            .I(N__10124));
    Odrv12 I__2267 (
            .O(N__10124),
            .I(A_c_0));
    IoInMux I__2266 (
            .O(N__10121),
            .I(N__10118));
    LocalMux I__2265 (
            .O(N__10118),
            .I(N__10115));
    Span4Mux_s2_v I__2264 (
            .O(N__10115),
            .I(N__10111));
    InMux I__2263 (
            .O(N__10114),
            .I(N__10108));
    Span4Mux_v I__2262 (
            .O(N__10111),
            .I(N__10105));
    LocalMux I__2261 (
            .O(N__10108),
            .I(N__10102));
    Odrv4 I__2260 (
            .O(N__10105),
            .I(UUBEn_c));
    Odrv12 I__2259 (
            .O(N__10102),
            .I(UUBEn_c));
    CascadeMux I__2258 (
            .O(N__10097),
            .I(N__10091));
    InMux I__2257 (
            .O(N__10096),
            .I(N__10083));
    InMux I__2256 (
            .O(N__10095),
            .I(N__10083));
    InMux I__2255 (
            .O(N__10094),
            .I(N__10083));
    InMux I__2254 (
            .O(N__10091),
            .I(N__10078));
    InMux I__2253 (
            .O(N__10090),
            .I(N__10078));
    LocalMux I__2252 (
            .O(N__10083),
            .I(N__10074));
    LocalMux I__2251 (
            .O(N__10078),
            .I(N__10071));
    InMux I__2250 (
            .O(N__10077),
            .I(N__10068));
    Span4Mux_v I__2249 (
            .O(N__10074),
            .I(N__10065));
    Span4Mux_v I__2248 (
            .O(N__10071),
            .I(N__10062));
    LocalMux I__2247 (
            .O(N__10068),
            .I(N__10059));
    Span4Mux_v I__2246 (
            .O(N__10065),
            .I(N__10056));
    Span4Mux_h I__2245 (
            .O(N__10062),
            .I(N__10051));
    Span4Mux_v I__2244 (
            .O(N__10059),
            .I(N__10051));
    Sp12to4 I__2243 (
            .O(N__10056),
            .I(N__10048));
    Span4Mux_v I__2242 (
            .O(N__10051),
            .I(N__10045));
    Span12Mux_h I__2241 (
            .O(N__10048),
            .I(N__10040));
    Sp12to4 I__2240 (
            .O(N__10045),
            .I(N__10040));
    Odrv12 I__2239 (
            .O(N__10040),
            .I(SIZ_c_0));
    InMux I__2238 (
            .O(N__10037),
            .I(N__10027));
    InMux I__2237 (
            .O(N__10036),
            .I(N__10027));
    InMux I__2236 (
            .O(N__10035),
            .I(N__10027));
    InMux I__2235 (
            .O(N__10034),
            .I(N__10024));
    LocalMux I__2234 (
            .O(N__10027),
            .I(N__10021));
    LocalMux I__2233 (
            .O(N__10024),
            .I(N__10018));
    Span4Mux_v I__2232 (
            .O(N__10021),
            .I(N__10015));
    Span4Mux_v I__2231 (
            .O(N__10018),
            .I(N__10012));
    Sp12to4 I__2230 (
            .O(N__10015),
            .I(N__10007));
    Sp12to4 I__2229 (
            .O(N__10012),
            .I(N__10007));
    Span12Mux_h I__2228 (
            .O(N__10007),
            .I(N__10004));
    Odrv12 I__2227 (
            .O(N__10004),
            .I(A_c_1));
    CascadeMux I__2226 (
            .O(N__10001),
            .I(N__9996));
    CascadeMux I__2225 (
            .O(N__10000),
            .I(N__9993));
    CascadeMux I__2224 (
            .O(N__9999),
            .I(N__9990));
    InMux I__2223 (
            .O(N__9996),
            .I(N__9984));
    InMux I__2222 (
            .O(N__9993),
            .I(N__9979));
    InMux I__2221 (
            .O(N__9990),
            .I(N__9979));
    InMux I__2220 (
            .O(N__9989),
            .I(N__9974));
    InMux I__2219 (
            .O(N__9988),
            .I(N__9974));
    InMux I__2218 (
            .O(N__9987),
            .I(N__9971));
    LocalMux I__2217 (
            .O(N__9984),
            .I(N__9964));
    LocalMux I__2216 (
            .O(N__9979),
            .I(N__9964));
    LocalMux I__2215 (
            .O(N__9974),
            .I(N__9964));
    LocalMux I__2214 (
            .O(N__9971),
            .I(N__9961));
    Sp12to4 I__2213 (
            .O(N__9964),
            .I(N__9958));
    Sp12to4 I__2212 (
            .O(N__9961),
            .I(N__9955));
    Span12Mux_v I__2211 (
            .O(N__9958),
            .I(N__9952));
    Span12Mux_v I__2210 (
            .O(N__9955),
            .I(N__9949));
    Span12Mux_h I__2209 (
            .O(N__9952),
            .I(N__9946));
    Span12Mux_h I__2208 (
            .O(N__9949),
            .I(N__9943));
    Odrv12 I__2207 (
            .O(N__9946),
            .I(SIZ_c_1));
    Odrv12 I__2206 (
            .O(N__9943),
            .I(SIZ_c_1));
    InMux I__2205 (
            .O(N__9938),
            .I(N__9933));
    InMux I__2204 (
            .O(N__9937),
            .I(N__9928));
    InMux I__2203 (
            .O(N__9936),
            .I(N__9928));
    LocalMux I__2202 (
            .O(N__9933),
            .I(\U712_CHIP_RAM.N_325_mux ));
    LocalMux I__2201 (
            .O(N__9928),
            .I(\U712_CHIP_RAM.N_325_mux ));
    IoInMux I__2200 (
            .O(N__9923),
            .I(N__9920));
    LocalMux I__2199 (
            .O(N__9920),
            .I(N__9917));
    IoSpan4Mux I__2198 (
            .O(N__9917),
            .I(N__9914));
    Span4Mux_s1_v I__2197 (
            .O(N__9914),
            .I(N__9911));
    Span4Mux_h I__2196 (
            .O(N__9911),
            .I(N__9907));
    InMux I__2195 (
            .O(N__9910),
            .I(N__9904));
    Sp12to4 I__2194 (
            .O(N__9907),
            .I(N__9899));
    LocalMux I__2193 (
            .O(N__9904),
            .I(N__9899));
    Odrv12 I__2192 (
            .O(N__9899),
            .I(UMBEn_c));
    InMux I__2191 (
            .O(N__9896),
            .I(N__9893));
    LocalMux I__2190 (
            .O(N__9893),
            .I(N__9888));
    CascadeMux I__2189 (
            .O(N__9892),
            .I(N__9885));
    CascadeMux I__2188 (
            .O(N__9891),
            .I(N__9881));
    Span4Mux_h I__2187 (
            .O(N__9888),
            .I(N__9877));
    InMux I__2186 (
            .O(N__9885),
            .I(N__9874));
    InMux I__2185 (
            .O(N__9884),
            .I(N__9870));
    InMux I__2184 (
            .O(N__9881),
            .I(N__9867));
    InMux I__2183 (
            .O(N__9880),
            .I(N__9864));
    Span4Mux_v I__2182 (
            .O(N__9877),
            .I(N__9859));
    LocalMux I__2181 (
            .O(N__9874),
            .I(N__9859));
    CascadeMux I__2180 (
            .O(N__9873),
            .I(N__9856));
    LocalMux I__2179 (
            .O(N__9870),
            .I(N__9849));
    LocalMux I__2178 (
            .O(N__9867),
            .I(N__9849));
    LocalMux I__2177 (
            .O(N__9864),
            .I(N__9846));
    Span4Mux_h I__2176 (
            .O(N__9859),
            .I(N__9843));
    InMux I__2175 (
            .O(N__9856),
            .I(N__9840));
    InMux I__2174 (
            .O(N__9855),
            .I(N__9837));
    InMux I__2173 (
            .O(N__9854),
            .I(N__9834));
    Odrv4 I__2172 (
            .O(N__9849),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__2171 (
            .O(N__9846),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__2170 (
            .O(N__9843),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__2169 (
            .O(N__9840),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__2168 (
            .O(N__9837),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__2167 (
            .O(N__9834),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    IoInMux I__2166 (
            .O(N__9821),
            .I(N__9818));
    LocalMux I__2165 (
            .O(N__9818),
            .I(N__9815));
    IoSpan4Mux I__2164 (
            .O(N__9815),
            .I(N__9812));
    Sp12to4 I__2163 (
            .O(N__9812),
            .I(N__9809));
    Span12Mux_s7_v I__2162 (
            .O(N__9809),
            .I(N__9806));
    Odrv12 I__2161 (
            .O(N__9806),
            .I(WEn_c));
    InMux I__2160 (
            .O(N__9803),
            .I(N__9800));
    LocalMux I__2159 (
            .O(N__9800),
            .I(N__9797));
    Odrv4 I__2158 (
            .O(N__9797),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__2157 (
            .O(N__9794),
            .I(N__9789));
    InMux I__2156 (
            .O(N__9793),
            .I(N__9786));
    InMux I__2155 (
            .O(N__9792),
            .I(N__9783));
    LocalMux I__2154 (
            .O(N__9789),
            .I(N__9775));
    LocalMux I__2153 (
            .O(N__9786),
            .I(N__9775));
    LocalMux I__2152 (
            .O(N__9783),
            .I(N__9775));
    InMux I__2151 (
            .O(N__9782),
            .I(N__9772));
    Span4Mux_v I__2150 (
            .O(N__9775),
            .I(N__9767));
    LocalMux I__2149 (
            .O(N__9772),
            .I(N__9767));
    Span4Mux_v I__2148 (
            .O(N__9767),
            .I(N__9764));
    Span4Mux_v I__2147 (
            .O(N__9764),
            .I(N__9761));
    Sp12to4 I__2146 (
            .O(N__9761),
            .I(N__9758));
    Span12Mux_h I__2145 (
            .O(N__9758),
            .I(N__9755));
    Odrv12 I__2144 (
            .O(N__9755),
            .I(DRA_c_4));
    InMux I__2143 (
            .O(N__9752),
            .I(N__9749));
    LocalMux I__2142 (
            .O(N__9749),
            .I(N__9746));
    Odrv12 I__2141 (
            .O(N__9746),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__2140 (
            .O(N__9743),
            .I(N__9737));
    InMux I__2139 (
            .O(N__9742),
            .I(N__9734));
    InMux I__2138 (
            .O(N__9741),
            .I(N__9729));
    InMux I__2137 (
            .O(N__9740),
            .I(N__9729));
    LocalMux I__2136 (
            .O(N__9737),
            .I(N__9722));
    LocalMux I__2135 (
            .O(N__9734),
            .I(N__9722));
    LocalMux I__2134 (
            .O(N__9729),
            .I(N__9722));
    Span4Mux_v I__2133 (
            .O(N__9722),
            .I(N__9719));
    Sp12to4 I__2132 (
            .O(N__9719),
            .I(N__9716));
    Span12Mux_h I__2131 (
            .O(N__9716),
            .I(N__9713));
    Span12Mux_v I__2130 (
            .O(N__9713),
            .I(N__9710));
    Odrv12 I__2129 (
            .O(N__9710),
            .I(DRA_c_5));
    InMux I__2128 (
            .O(N__9707),
            .I(N__9704));
    LocalMux I__2127 (
            .O(N__9704),
            .I(N__9701));
    Odrv4 I__2126 (
            .O(N__9701),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__2125 (
            .O(N__9698),
            .I(N__9695));
    LocalMux I__2124 (
            .O(N__9695),
            .I(\U712_CHIP_RAM.m191_1 ));
    IoInMux I__2123 (
            .O(N__9692),
            .I(N__9689));
    LocalMux I__2122 (
            .O(N__9689),
            .I(N__9686));
    IoSpan4Mux I__2121 (
            .O(N__9686),
            .I(N__9683));
    IoSpan4Mux I__2120 (
            .O(N__9683),
            .I(N__9680));
    Span4Mux_s3_h I__2119 (
            .O(N__9680),
            .I(N__9677));
    Sp12to4 I__2118 (
            .O(N__9677),
            .I(N__9674));
    Odrv12 I__2117 (
            .O(N__9674),
            .I(CMA_c_7));
    CEMux I__2116 (
            .O(N__9671),
            .I(N__9668));
    LocalMux I__2115 (
            .O(N__9668),
            .I(N__9663));
    CEMux I__2114 (
            .O(N__9667),
            .I(N__9660));
    CEMux I__2113 (
            .O(N__9666),
            .I(N__9657));
    Span4Mux_v I__2112 (
            .O(N__9663),
            .I(N__9654));
    LocalMux I__2111 (
            .O(N__9660),
            .I(N__9651));
    LocalMux I__2110 (
            .O(N__9657),
            .I(N__9648));
    Span4Mux_h I__2109 (
            .O(N__9654),
            .I(N__9642));
    Span4Mux_h I__2108 (
            .O(N__9651),
            .I(N__9637));
    Span4Mux_h I__2107 (
            .O(N__9648),
            .I(N__9637));
    CEMux I__2106 (
            .O(N__9647),
            .I(N__9634));
    CEMux I__2105 (
            .O(N__9646),
            .I(N__9631));
    CEMux I__2104 (
            .O(N__9645),
            .I(N__9628));
    Odrv4 I__2103 (
            .O(N__9642),
            .I(\U712_CHIP_RAM.N_198_0 ));
    Odrv4 I__2102 (
            .O(N__9637),
            .I(\U712_CHIP_RAM.N_198_0 ));
    LocalMux I__2101 (
            .O(N__9634),
            .I(\U712_CHIP_RAM.N_198_0 ));
    LocalMux I__2100 (
            .O(N__9631),
            .I(\U712_CHIP_RAM.N_198_0 ));
    LocalMux I__2099 (
            .O(N__9628),
            .I(\U712_CHIP_RAM.N_198_0 ));
    InMux I__2098 (
            .O(N__9617),
            .I(N__9614));
    LocalMux I__2097 (
            .O(N__9614),
            .I(N__9611));
    Odrv12 I__2096 (
            .O(N__9611),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__2095 (
            .O(N__9608),
            .I(N__9605));
    LocalMux I__2094 (
            .O(N__9605),
            .I(N__9602));
    Odrv4 I__2093 (
            .O(N__9602),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__2092 (
            .O(N__9599),
            .I(N__9596));
    LocalMux I__2091 (
            .O(N__9596),
            .I(N__9593));
    Odrv4 I__2090 (
            .O(N__9593),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__2089 (
            .O(N__9590),
            .I(N__9587));
    LocalMux I__2088 (
            .O(N__9587),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__2087 (
            .O(N__9584),
            .I(N__9581));
    LocalMux I__2086 (
            .O(N__9581),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    IoInMux I__2085 (
            .O(N__9578),
            .I(N__9575));
    LocalMux I__2084 (
            .O(N__9575),
            .I(N__9572));
    Span4Mux_s2_h I__2083 (
            .O(N__9572),
            .I(N__9569));
    Span4Mux_v I__2082 (
            .O(N__9569),
            .I(N__9566));
    Sp12to4 I__2081 (
            .O(N__9566),
            .I(N__9563));
    Span12Mux_h I__2080 (
            .O(N__9563),
            .I(N__9560));
    Span12Mux_v I__2079 (
            .O(N__9560),
            .I(N__9557));
    Odrv12 I__2078 (
            .O(N__9557),
            .I(CUMBEn_c));
    IoInMux I__2077 (
            .O(N__9554),
            .I(N__9551));
    LocalMux I__2076 (
            .O(N__9551),
            .I(N__9548));
    Span4Mux_s1_v I__2075 (
            .O(N__9548),
            .I(N__9544));
    InMux I__2074 (
            .O(N__9547),
            .I(N__9541));
    Span4Mux_v I__2073 (
            .O(N__9544),
            .I(N__9538));
    LocalMux I__2072 (
            .O(N__9541),
            .I(N__9535));
    Span4Mux_v I__2071 (
            .O(N__9538),
            .I(N__9532));
    Span4Mux_v I__2070 (
            .O(N__9535),
            .I(N__9529));
    Odrv4 I__2069 (
            .O(N__9532),
            .I(LMBEn_c));
    Odrv4 I__2068 (
            .O(N__9529),
            .I(LMBEn_c));
    IoInMux I__2067 (
            .O(N__9524),
            .I(N__9521));
    LocalMux I__2066 (
            .O(N__9521),
            .I(N__9518));
    Span4Mux_s2_h I__2065 (
            .O(N__9518),
            .I(N__9515));
    Sp12to4 I__2064 (
            .O(N__9515),
            .I(N__9512));
    Span12Mux_s10_v I__2063 (
            .O(N__9512),
            .I(N__9509));
    Span12Mux_h I__2062 (
            .O(N__9509),
            .I(N__9506));
    Odrv12 I__2061 (
            .O(N__9506),
            .I(CLMBEn_c));
    IoInMux I__2060 (
            .O(N__9503),
            .I(N__9500));
    LocalMux I__2059 (
            .O(N__9500),
            .I(N__9497));
    Span4Mux_s2_h I__2058 (
            .O(N__9497),
            .I(N__9494));
    Sp12to4 I__2057 (
            .O(N__9494),
            .I(N__9491));
    Span12Mux_v I__2056 (
            .O(N__9491),
            .I(N__9488));
    Odrv12 I__2055 (
            .O(N__9488),
            .I(CUUBEn_c));
    IoInMux I__2054 (
            .O(N__9485),
            .I(N__9482));
    LocalMux I__2053 (
            .O(N__9482),
            .I(N__9479));
    Span12Mux_s7_v I__2052 (
            .O(N__9479),
            .I(N__9476));
    Span12Mux_h I__2051 (
            .O(N__9476),
            .I(N__9473));
    Odrv12 I__2050 (
            .O(N__9473),
            .I(ASn_c));
    CEMux I__2049 (
            .O(N__9470),
            .I(N__9467));
    LocalMux I__2048 (
            .O(N__9467),
            .I(N__9464));
    Span4Mux_v I__2047 (
            .O(N__9464),
            .I(N__9461));
    Odrv4 I__2046 (
            .O(N__9461),
            .I(\U712_REG_SM.N_99_0_0 ));
    CascadeMux I__2045 (
            .O(N__9458),
            .I(N__9454));
    InMux I__2044 (
            .O(N__9457),
            .I(N__9447));
    InMux I__2043 (
            .O(N__9454),
            .I(N__9444));
    InMux I__2042 (
            .O(N__9453),
            .I(N__9441));
    InMux I__2041 (
            .O(N__9452),
            .I(N__9436));
    InMux I__2040 (
            .O(N__9451),
            .I(N__9432));
    CascadeMux I__2039 (
            .O(N__9450),
            .I(N__9427));
    LocalMux I__2038 (
            .O(N__9447),
            .I(N__9422));
    LocalMux I__2037 (
            .O(N__9444),
            .I(N__9419));
    LocalMux I__2036 (
            .O(N__9441),
            .I(N__9416));
    InMux I__2035 (
            .O(N__9440),
            .I(N__9411));
    CascadeMux I__2034 (
            .O(N__9439),
            .I(N__9408));
    LocalMux I__2033 (
            .O(N__9436),
            .I(N__9405));
    InMux I__2032 (
            .O(N__9435),
            .I(N__9402));
    LocalMux I__2031 (
            .O(N__9432),
            .I(N__9399));
    InMux I__2030 (
            .O(N__9431),
            .I(N__9396));
    InMux I__2029 (
            .O(N__9430),
            .I(N__9389));
    InMux I__2028 (
            .O(N__9427),
            .I(N__9389));
    InMux I__2027 (
            .O(N__9426),
            .I(N__9389));
    InMux I__2026 (
            .O(N__9425),
            .I(N__9386));
    Span4Mux_h I__2025 (
            .O(N__9422),
            .I(N__9381));
    Span4Mux_v I__2024 (
            .O(N__9419),
            .I(N__9381));
    Span4Mux_v I__2023 (
            .O(N__9416),
            .I(N__9378));
    InMux I__2022 (
            .O(N__9415),
            .I(N__9373));
    InMux I__2021 (
            .O(N__9414),
            .I(N__9373));
    LocalMux I__2020 (
            .O(N__9411),
            .I(N__9370));
    InMux I__2019 (
            .O(N__9408),
            .I(N__9367));
    Span4Mux_h I__2018 (
            .O(N__9405),
            .I(N__9362));
    LocalMux I__2017 (
            .O(N__9402),
            .I(N__9362));
    Odrv12 I__2016 (
            .O(N__9399),
            .I(U712_REG_SM_C1_SYNC_1));
    LocalMux I__2015 (
            .O(N__9396),
            .I(U712_REG_SM_C1_SYNC_1));
    LocalMux I__2014 (
            .O(N__9389),
            .I(U712_REG_SM_C1_SYNC_1));
    LocalMux I__2013 (
            .O(N__9386),
            .I(U712_REG_SM_C1_SYNC_1));
    Odrv4 I__2012 (
            .O(N__9381),
            .I(U712_REG_SM_C1_SYNC_1));
    Odrv4 I__2011 (
            .O(N__9378),
            .I(U712_REG_SM_C1_SYNC_1));
    LocalMux I__2010 (
            .O(N__9373),
            .I(U712_REG_SM_C1_SYNC_1));
    Odrv4 I__2009 (
            .O(N__9370),
            .I(U712_REG_SM_C1_SYNC_1));
    LocalMux I__2008 (
            .O(N__9367),
            .I(U712_REG_SM_C1_SYNC_1));
    Odrv4 I__2007 (
            .O(N__9362),
            .I(U712_REG_SM_C1_SYNC_1));
    InMux I__2006 (
            .O(N__9341),
            .I(N__9338));
    LocalMux I__2005 (
            .O(N__9338),
            .I(U712_REG_SM_LDSn_6_0));
    InMux I__2004 (
            .O(N__9335),
            .I(N__9332));
    LocalMux I__2003 (
            .O(N__9332),
            .I(\U712_CHIP_RAM.m185_1 ));
    IoInMux I__2002 (
            .O(N__9329),
            .I(N__9326));
    LocalMux I__2001 (
            .O(N__9326),
            .I(N__9323));
    Span4Mux_s3_h I__2000 (
            .O(N__9323),
            .I(N__9320));
    Span4Mux_v I__1999 (
            .O(N__9320),
            .I(N__9317));
    Sp12to4 I__1998 (
            .O(N__9317),
            .I(N__9314));
    Span12Mux_h I__1997 (
            .O(N__9314),
            .I(N__9311));
    Odrv12 I__1996 (
            .O(N__9311),
            .I(CMA_c_5));
    InMux I__1995 (
            .O(N__9308),
            .I(N__9305));
    LocalMux I__1994 (
            .O(N__9305),
            .I(N__9302));
    Span4Mux_h I__1993 (
            .O(N__9302),
            .I(N__9299));
    Odrv4 I__1992 (
            .O(N__9299),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__1991 (
            .O(N__9296),
            .I(N__9293));
    LocalMux I__1990 (
            .O(N__9293),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__1989 (
            .O(N__9290),
            .I(N__9287));
    LocalMux I__1988 (
            .O(N__9287),
            .I(N__9284));
    Span4Mux_v I__1987 (
            .O(N__9284),
            .I(N__9281));
    Span4Mux_v I__1986 (
            .O(N__9281),
            .I(N__9278));
    Sp12to4 I__1985 (
            .O(N__9278),
            .I(N__9275));
    Span12Mux_h I__1984 (
            .O(N__9275),
            .I(N__9272));
    Odrv12 I__1983 (
            .O(N__9272),
            .I(A_c_19));
    InMux I__1982 (
            .O(N__9269),
            .I(N__9266));
    LocalMux I__1981 (
            .O(N__9266),
            .I(\U712_CHIP_RAM.m194_0 ));
    IoInMux I__1980 (
            .O(N__9263),
            .I(N__9260));
    LocalMux I__1979 (
            .O(N__9260),
            .I(N__9257));
    Span4Mux_s3_h I__1978 (
            .O(N__9257),
            .I(N__9254));
    Span4Mux_v I__1977 (
            .O(N__9254),
            .I(N__9251));
    Sp12to4 I__1976 (
            .O(N__9251),
            .I(N__9248));
    Span12Mux_h I__1975 (
            .O(N__9248),
            .I(N__9245));
    Odrv12 I__1974 (
            .O(N__9245),
            .I(CMA_c_9));
    InMux I__1973 (
            .O(N__9242),
            .I(N__9238));
    InMux I__1972 (
            .O(N__9241),
            .I(N__9235));
    LocalMux I__1971 (
            .O(N__9238),
            .I(N__9229));
    LocalMux I__1970 (
            .O(N__9235),
            .I(N__9225));
    InMux I__1969 (
            .O(N__9234),
            .I(N__9222));
    InMux I__1968 (
            .O(N__9233),
            .I(N__9217));
    InMux I__1967 (
            .O(N__9232),
            .I(N__9214));
    Span4Mux_h I__1966 (
            .O(N__9229),
            .I(N__9211));
    InMux I__1965 (
            .O(N__9228),
            .I(N__9208));
    Span12Mux_v I__1964 (
            .O(N__9225),
            .I(N__9205));
    LocalMux I__1963 (
            .O(N__9222),
            .I(N__9202));
    InMux I__1962 (
            .O(N__9221),
            .I(N__9199));
    InMux I__1961 (
            .O(N__9220),
            .I(N__9196));
    LocalMux I__1960 (
            .O(N__9217),
            .I(N__9187));
    LocalMux I__1959 (
            .O(N__9214),
            .I(N__9187));
    Span4Mux_v I__1958 (
            .O(N__9211),
            .I(N__9187));
    LocalMux I__1957 (
            .O(N__9208),
            .I(N__9187));
    Odrv12 I__1956 (
            .O(N__9205),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1955 (
            .O(N__9202),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1954 (
            .O(N__9199),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1953 (
            .O(N__9196),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1952 (
            .O(N__9187),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    InMux I__1951 (
            .O(N__9176),
            .I(N__9173));
    LocalMux I__1950 (
            .O(N__9173),
            .I(N__9170));
    Odrv4 I__1949 (
            .O(N__9170),
            .I(\U712_CHIP_RAM.d_N_7_0 ));
    InMux I__1948 (
            .O(N__9167),
            .I(N__9164));
    LocalMux I__1947 (
            .O(N__9164),
            .I(N__9161));
    Span4Mux_v I__1946 (
            .O(N__9161),
            .I(N__9158));
    Sp12to4 I__1945 (
            .O(N__9158),
            .I(N__9155));
    Span12Mux_v I__1944 (
            .O(N__9155),
            .I(N__9152));
    Span12Mux_h I__1943 (
            .O(N__9152),
            .I(N__9149));
    Odrv12 I__1942 (
            .O(N__9149),
            .I(A_c_18));
    InMux I__1941 (
            .O(N__9146),
            .I(N__9142));
    InMux I__1940 (
            .O(N__9145),
            .I(N__9139));
    LocalMux I__1939 (
            .O(N__9142),
            .I(N__9136));
    LocalMux I__1938 (
            .O(N__9139),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ));
    Odrv4 I__1937 (
            .O(N__9136),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ));
    CascadeMux I__1936 (
            .O(N__9131),
            .I(N__9127));
    InMux I__1935 (
            .O(N__9130),
            .I(N__9115));
    InMux I__1934 (
            .O(N__9127),
            .I(N__9112));
    InMux I__1933 (
            .O(N__9126),
            .I(N__9107));
    InMux I__1932 (
            .O(N__9125),
            .I(N__9107));
    InMux I__1931 (
            .O(N__9124),
            .I(N__9104));
    InMux I__1930 (
            .O(N__9123),
            .I(N__9099));
    InMux I__1929 (
            .O(N__9122),
            .I(N__9096));
    CascadeMux I__1928 (
            .O(N__9121),
            .I(N__9093));
    CascadeMux I__1927 (
            .O(N__9120),
            .I(N__9090));
    InMux I__1926 (
            .O(N__9119),
            .I(N__9081));
    InMux I__1925 (
            .O(N__9118),
            .I(N__9081));
    LocalMux I__1924 (
            .O(N__9115),
            .I(N__9078));
    LocalMux I__1923 (
            .O(N__9112),
            .I(N__9071));
    LocalMux I__1922 (
            .O(N__9107),
            .I(N__9071));
    LocalMux I__1921 (
            .O(N__9104),
            .I(N__9071));
    InMux I__1920 (
            .O(N__9103),
            .I(N__9068));
    InMux I__1919 (
            .O(N__9102),
            .I(N__9065));
    LocalMux I__1918 (
            .O(N__9099),
            .I(N__9062));
    LocalMux I__1917 (
            .O(N__9096),
            .I(N__9059));
    InMux I__1916 (
            .O(N__9093),
            .I(N__9056));
    InMux I__1915 (
            .O(N__9090),
            .I(N__9049));
    InMux I__1914 (
            .O(N__9089),
            .I(N__9049));
    InMux I__1913 (
            .O(N__9088),
            .I(N__9049));
    InMux I__1912 (
            .O(N__9087),
            .I(N__9044));
    InMux I__1911 (
            .O(N__9086),
            .I(N__9044));
    LocalMux I__1910 (
            .O(N__9081),
            .I(N__9037));
    Span4Mux_h I__1909 (
            .O(N__9078),
            .I(N__9037));
    Span4Mux_h I__1908 (
            .O(N__9071),
            .I(N__9037));
    LocalMux I__1907 (
            .O(N__9068),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1906 (
            .O(N__9065),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1905 (
            .O(N__9062),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1904 (
            .O(N__9059),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1903 (
            .O(N__9056),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1902 (
            .O(N__9049),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1901 (
            .O(N__9044),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1900 (
            .O(N__9037),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    InMux I__1899 (
            .O(N__9020),
            .I(N__9017));
    LocalMux I__1898 (
            .O(N__9017),
            .I(\U712_CHIP_RAM.N_204 ));
    InMux I__1897 (
            .O(N__9014),
            .I(N__9011));
    LocalMux I__1896 (
            .O(N__9011),
            .I(N__9008));
    Span4Mux_h I__1895 (
            .O(N__9008),
            .I(N__9005));
    Sp12to4 I__1894 (
            .O(N__9005),
            .I(N__9002));
    Span12Mux_v I__1893 (
            .O(N__9002),
            .I(N__8999));
    Span12Mux_h I__1892 (
            .O(N__8999),
            .I(N__8996));
    Odrv12 I__1891 (
            .O(N__8996),
            .I(A_c_3));
    InMux I__1890 (
            .O(N__8993),
            .I(N__8989));
    InMux I__1889 (
            .O(N__8992),
            .I(N__8986));
    LocalMux I__1888 (
            .O(N__8989),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ));
    LocalMux I__1887 (
            .O(N__8986),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ));
    InMux I__1886 (
            .O(N__8981),
            .I(N__8967));
    InMux I__1885 (
            .O(N__8980),
            .I(N__8967));
    InMux I__1884 (
            .O(N__8979),
            .I(N__8967));
    InMux I__1883 (
            .O(N__8978),
            .I(N__8962));
    InMux I__1882 (
            .O(N__8977),
            .I(N__8962));
    InMux I__1881 (
            .O(N__8976),
            .I(N__8955));
    InMux I__1880 (
            .O(N__8975),
            .I(N__8955));
    InMux I__1879 (
            .O(N__8974),
            .I(N__8955));
    LocalMux I__1878 (
            .O(N__8967),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ));
    LocalMux I__1877 (
            .O(N__8962),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ));
    LocalMux I__1876 (
            .O(N__8955),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ));
    InMux I__1875 (
            .O(N__8948),
            .I(N__8945));
    LocalMux I__1874 (
            .O(N__8945),
            .I(N__8942));
    Span12Mux_h I__1873 (
            .O(N__8942),
            .I(N__8939));
    Odrv12 I__1872 (
            .O(N__8939),
            .I(A_c_8));
    InMux I__1871 (
            .O(N__8936),
            .I(N__8932));
    InMux I__1870 (
            .O(N__8935),
            .I(N__8929));
    LocalMux I__1869 (
            .O(N__8932),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ));
    LocalMux I__1868 (
            .O(N__8929),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ));
    InMux I__1867 (
            .O(N__8924),
            .I(N__8916));
    InMux I__1866 (
            .O(N__8923),
            .I(N__8910));
    InMux I__1865 (
            .O(N__8922),
            .I(N__8907));
    InMux I__1864 (
            .O(N__8921),
            .I(N__8900));
    InMux I__1863 (
            .O(N__8920),
            .I(N__8900));
    InMux I__1862 (
            .O(N__8919),
            .I(N__8900));
    LocalMux I__1861 (
            .O(N__8916),
            .I(N__8896));
    InMux I__1860 (
            .O(N__8915),
            .I(N__8889));
    InMux I__1859 (
            .O(N__8914),
            .I(N__8889));
    InMux I__1858 (
            .O(N__8913),
            .I(N__8889));
    LocalMux I__1857 (
            .O(N__8910),
            .I(N__8875));
    LocalMux I__1856 (
            .O(N__8907),
            .I(N__8875));
    LocalMux I__1855 (
            .O(N__8900),
            .I(N__8875));
    CascadeMux I__1854 (
            .O(N__8899),
            .I(N__8868));
    Span4Mux_v I__1853 (
            .O(N__8896),
            .I(N__8861));
    LocalMux I__1852 (
            .O(N__8889),
            .I(N__8861));
    InMux I__1851 (
            .O(N__8888),
            .I(N__8854));
    InMux I__1850 (
            .O(N__8887),
            .I(N__8854));
    InMux I__1849 (
            .O(N__8886),
            .I(N__8854));
    InMux I__1848 (
            .O(N__8885),
            .I(N__8847));
    InMux I__1847 (
            .O(N__8884),
            .I(N__8847));
    InMux I__1846 (
            .O(N__8883),
            .I(N__8847));
    CascadeMux I__1845 (
            .O(N__8882),
            .I(N__8842));
    Span4Mux_v I__1844 (
            .O(N__8875),
            .I(N__8838));
    InMux I__1843 (
            .O(N__8874),
            .I(N__8833));
    InMux I__1842 (
            .O(N__8873),
            .I(N__8833));
    InMux I__1841 (
            .O(N__8872),
            .I(N__8830));
    InMux I__1840 (
            .O(N__8871),
            .I(N__8821));
    InMux I__1839 (
            .O(N__8868),
            .I(N__8821));
    InMux I__1838 (
            .O(N__8867),
            .I(N__8821));
    InMux I__1837 (
            .O(N__8866),
            .I(N__8821));
    Span4Mux_h I__1836 (
            .O(N__8861),
            .I(N__8816));
    LocalMux I__1835 (
            .O(N__8854),
            .I(N__8816));
    LocalMux I__1834 (
            .O(N__8847),
            .I(N__8813));
    InMux I__1833 (
            .O(N__8846),
            .I(N__8808));
    InMux I__1832 (
            .O(N__8845),
            .I(N__8808));
    InMux I__1831 (
            .O(N__8842),
            .I(N__8803));
    InMux I__1830 (
            .O(N__8841),
            .I(N__8803));
    Odrv4 I__1829 (
            .O(N__8838),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1828 (
            .O(N__8833),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1827 (
            .O(N__8830),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1826 (
            .O(N__8821),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1825 (
            .O(N__8816),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1824 (
            .O(N__8813),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1823 (
            .O(N__8808),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1822 (
            .O(N__8803),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__1821 (
            .O(N__8786),
            .I(N__8781));
    InMux I__1820 (
            .O(N__8785),
            .I(N__8776));
    CascadeMux I__1819 (
            .O(N__8784),
            .I(N__8773));
    LocalMux I__1818 (
            .O(N__8781),
            .I(N__8768));
    InMux I__1817 (
            .O(N__8780),
            .I(N__8763));
    InMux I__1816 (
            .O(N__8779),
            .I(N__8763));
    LocalMux I__1815 (
            .O(N__8776),
            .I(N__8760));
    InMux I__1814 (
            .O(N__8773),
            .I(N__8757));
    InMux I__1813 (
            .O(N__8772),
            .I(N__8754));
    InMux I__1812 (
            .O(N__8771),
            .I(N__8751));
    Odrv4 I__1811 (
            .O(N__8768),
            .I(\U712_CHIP_RAM.N_31_0 ));
    LocalMux I__1810 (
            .O(N__8763),
            .I(\U712_CHIP_RAM.N_31_0 ));
    Odrv4 I__1809 (
            .O(N__8760),
            .I(\U712_CHIP_RAM.N_31_0 ));
    LocalMux I__1808 (
            .O(N__8757),
            .I(\U712_CHIP_RAM.N_31_0 ));
    LocalMux I__1807 (
            .O(N__8754),
            .I(\U712_CHIP_RAM.N_31_0 ));
    LocalMux I__1806 (
            .O(N__8751),
            .I(\U712_CHIP_RAM.N_31_0 ));
    CascadeMux I__1805 (
            .O(N__8738),
            .I(N__8735));
    InMux I__1804 (
            .O(N__8735),
            .I(N__8732));
    LocalMux I__1803 (
            .O(N__8732),
            .I(\U712_CHIP_RAM.DBENn_8_0 ));
    IoInMux I__1802 (
            .O(N__8729),
            .I(N__8726));
    LocalMux I__1801 (
            .O(N__8726),
            .I(N__8723));
    IoSpan4Mux I__1800 (
            .O(N__8723),
            .I(N__8720));
    Sp12to4 I__1799 (
            .O(N__8720),
            .I(N__8716));
    InMux I__1798 (
            .O(N__8719),
            .I(N__8713));
    Span12Mux_s7_v I__1797 (
            .O(N__8716),
            .I(N__8710));
    LocalMux I__1796 (
            .O(N__8713),
            .I(N__8707));
    Odrv12 I__1795 (
            .O(N__8710),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1794 (
            .O(N__8707),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__1793 (
            .O(N__8702),
            .I(N__8699));
    InMux I__1792 (
            .O(N__8699),
            .I(N__8696));
    LocalMux I__1791 (
            .O(N__8696),
            .I(N__8693));
    Span4Mux_h I__1790 (
            .O(N__8693),
            .I(N__8690));
    Odrv4 I__1789 (
            .O(N__8690),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ));
    CascadeMux I__1788 (
            .O(N__8687),
            .I(N__8682));
    CascadeMux I__1787 (
            .O(N__8686),
            .I(N__8677));
    CascadeMux I__1786 (
            .O(N__8685),
            .I(N__8673));
    InMux I__1785 (
            .O(N__8682),
            .I(N__8659));
    InMux I__1784 (
            .O(N__8681),
            .I(N__8659));
    CascadeMux I__1783 (
            .O(N__8680),
            .I(N__8655));
    InMux I__1782 (
            .O(N__8677),
            .I(N__8650));
    InMux I__1781 (
            .O(N__8676),
            .I(N__8647));
    InMux I__1780 (
            .O(N__8673),
            .I(N__8642));
    InMux I__1779 (
            .O(N__8672),
            .I(N__8642));
    InMux I__1778 (
            .O(N__8671),
            .I(N__8636));
    InMux I__1777 (
            .O(N__8670),
            .I(N__8629));
    InMux I__1776 (
            .O(N__8669),
            .I(N__8629));
    InMux I__1775 (
            .O(N__8668),
            .I(N__8629));
    InMux I__1774 (
            .O(N__8667),
            .I(N__8618));
    InMux I__1773 (
            .O(N__8666),
            .I(N__8618));
    InMux I__1772 (
            .O(N__8665),
            .I(N__8618));
    InMux I__1771 (
            .O(N__8664),
            .I(N__8615));
    LocalMux I__1770 (
            .O(N__8659),
            .I(N__8612));
    InMux I__1769 (
            .O(N__8658),
            .I(N__8603));
    InMux I__1768 (
            .O(N__8655),
            .I(N__8603));
    InMux I__1767 (
            .O(N__8654),
            .I(N__8603));
    InMux I__1766 (
            .O(N__8653),
            .I(N__8603));
    LocalMux I__1765 (
            .O(N__8650),
            .I(N__8596));
    LocalMux I__1764 (
            .O(N__8647),
            .I(N__8596));
    LocalMux I__1763 (
            .O(N__8642),
            .I(N__8596));
    CascadeMux I__1762 (
            .O(N__8641),
            .I(N__8590));
    InMux I__1761 (
            .O(N__8640),
            .I(N__8586));
    InMux I__1760 (
            .O(N__8639),
            .I(N__8582));
    LocalMux I__1759 (
            .O(N__8636),
            .I(N__8577));
    LocalMux I__1758 (
            .O(N__8629),
            .I(N__8577));
    InMux I__1757 (
            .O(N__8628),
            .I(N__8570));
    InMux I__1756 (
            .O(N__8627),
            .I(N__8570));
    InMux I__1755 (
            .O(N__8626),
            .I(N__8570));
    InMux I__1754 (
            .O(N__8625),
            .I(N__8567));
    LocalMux I__1753 (
            .O(N__8618),
            .I(N__8564));
    LocalMux I__1752 (
            .O(N__8615),
            .I(N__8555));
    Span4Mux_v I__1751 (
            .O(N__8612),
            .I(N__8555));
    LocalMux I__1750 (
            .O(N__8603),
            .I(N__8555));
    Span4Mux_v I__1749 (
            .O(N__8596),
            .I(N__8555));
    InMux I__1748 (
            .O(N__8595),
            .I(N__8548));
    InMux I__1747 (
            .O(N__8594),
            .I(N__8548));
    InMux I__1746 (
            .O(N__8593),
            .I(N__8548));
    InMux I__1745 (
            .O(N__8590),
            .I(N__8545));
    InMux I__1744 (
            .O(N__8589),
            .I(N__8542));
    LocalMux I__1743 (
            .O(N__8586),
            .I(N__8539));
    InMux I__1742 (
            .O(N__8585),
            .I(N__8536));
    LocalMux I__1741 (
            .O(N__8582),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1740 (
            .O(N__8577),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1739 (
            .O(N__8570),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1738 (
            .O(N__8567),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1737 (
            .O(N__8564),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1736 (
            .O(N__8555),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1735 (
            .O(N__8548),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1734 (
            .O(N__8545),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1733 (
            .O(N__8542),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv12 I__1732 (
            .O(N__8539),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1731 (
            .O(N__8536),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    InMux I__1730 (
            .O(N__8513),
            .I(N__8510));
    LocalMux I__1729 (
            .O(N__8510),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0 ));
    IoInMux I__1728 (
            .O(N__8507),
            .I(N__8504));
    LocalMux I__1727 (
            .O(N__8504),
            .I(N__8501));
    Span12Mux_s1_v I__1726 (
            .O(N__8501),
            .I(N__8498));
    Span12Mux_v I__1725 (
            .O(N__8498),
            .I(N__8494));
    InMux I__1724 (
            .O(N__8497),
            .I(N__8491));
    Odrv12 I__1723 (
            .O(N__8494),
            .I(LATCH_CLK_c));
    LocalMux I__1722 (
            .O(N__8491),
            .I(LATCH_CLK_c));
    CascadeMux I__1721 (
            .O(N__8486),
            .I(\U712_CHIP_RAM.m191_0_cascade_ ));
    InMux I__1720 (
            .O(N__8483),
            .I(N__8480));
    LocalMux I__1719 (
            .O(N__8480),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__1718 (
            .O(N__8477),
            .I(N__8474));
    LocalMux I__1717 (
            .O(N__8474),
            .I(\U712_CHIP_RAM.d_N_6_4 ));
    IoInMux I__1716 (
            .O(N__8471),
            .I(N__8468));
    LocalMux I__1715 (
            .O(N__8468),
            .I(N__8465));
    Span4Mux_s0_v I__1714 (
            .O(N__8465),
            .I(N__8462));
    Span4Mux_v I__1713 (
            .O(N__8462),
            .I(N__8458));
    InMux I__1712 (
            .O(N__8461),
            .I(N__8455));
    Span4Mux_v I__1711 (
            .O(N__8458),
            .I(N__8452));
    LocalMux I__1710 (
            .O(N__8455),
            .I(N__8449));
    Sp12to4 I__1709 (
            .O(N__8452),
            .I(N__8446));
    Span4Mux_v I__1708 (
            .O(N__8449),
            .I(N__8443));
    Span12Mux_h I__1707 (
            .O(N__8446),
            .I(N__8440));
    Sp12to4 I__1706 (
            .O(N__8443),
            .I(N__8437));
    Span12Mux_v I__1705 (
            .O(N__8440),
            .I(N__8432));
    Span12Mux_h I__1704 (
            .O(N__8437),
            .I(N__8432));
    Odrv12 I__1703 (
            .O(N__8432),
            .I(A_c_10));
    CascadeMux I__1702 (
            .O(N__8429),
            .I(N__8426));
    InMux I__1701 (
            .O(N__8426),
            .I(N__8422));
    InMux I__1700 (
            .O(N__8425),
            .I(N__8419));
    LocalMux I__1699 (
            .O(N__8422),
            .I(N__8416));
    LocalMux I__1698 (
            .O(N__8419),
            .I(N__8413));
    Span4Mux_h I__1697 (
            .O(N__8416),
            .I(N__8410));
    Span4Mux_v I__1696 (
            .O(N__8413),
            .I(N__8405));
    Span4Mux_v I__1695 (
            .O(N__8410),
            .I(N__8405));
    Odrv4 I__1694 (
            .O(N__8405),
            .I(\U712_CHIP_RAM.m184_m2_0_a2_0 ));
    CascadeMux I__1693 (
            .O(N__8402),
            .I(\U712_CHIP_RAM.m184_0_cascade_ ));
    InMux I__1692 (
            .O(N__8399),
            .I(N__8396));
    LocalMux I__1691 (
            .O(N__8396),
            .I(\U712_CHIP_RAM.m184_1 ));
    InMux I__1690 (
            .O(N__8393),
            .I(N__8390));
    LocalMux I__1689 (
            .O(N__8390),
            .I(N__8387));
    Span4Mux_v I__1688 (
            .O(N__8387),
            .I(N__8384));
    Span4Mux_v I__1687 (
            .O(N__8384),
            .I(N__8381));
    Sp12to4 I__1686 (
            .O(N__8381),
            .I(N__8378));
    Span12Mux_h I__1685 (
            .O(N__8378),
            .I(N__8375));
    Odrv12 I__1684 (
            .O(N__8375),
            .I(A_c_15));
    InMux I__1683 (
            .O(N__8372),
            .I(N__8365));
    CascadeMux I__1682 (
            .O(N__8371),
            .I(N__8362));
    InMux I__1681 (
            .O(N__8370),
            .I(N__8357));
    CascadeMux I__1680 (
            .O(N__8369),
            .I(N__8351));
    InMux I__1679 (
            .O(N__8368),
            .I(N__8348));
    LocalMux I__1678 (
            .O(N__8365),
            .I(N__8345));
    InMux I__1677 (
            .O(N__8362),
            .I(N__8338));
    InMux I__1676 (
            .O(N__8361),
            .I(N__8338));
    InMux I__1675 (
            .O(N__8360),
            .I(N__8338));
    LocalMux I__1674 (
            .O(N__8357),
            .I(N__8335));
    InMux I__1673 (
            .O(N__8356),
            .I(N__8330));
    InMux I__1672 (
            .O(N__8355),
            .I(N__8330));
    InMux I__1671 (
            .O(N__8354),
            .I(N__8325));
    InMux I__1670 (
            .O(N__8351),
            .I(N__8325));
    LocalMux I__1669 (
            .O(N__8348),
            .I(N__8322));
    Span4Mux_h I__1668 (
            .O(N__8345),
            .I(N__8317));
    LocalMux I__1667 (
            .O(N__8338),
            .I(N__8317));
    Odrv12 I__1666 (
            .O(N__8335),
            .I(\U712_CHIP_RAM.N_3_0 ));
    LocalMux I__1665 (
            .O(N__8330),
            .I(\U712_CHIP_RAM.N_3_0 ));
    LocalMux I__1664 (
            .O(N__8325),
            .I(\U712_CHIP_RAM.N_3_0 ));
    Odrv4 I__1663 (
            .O(N__8322),
            .I(\U712_CHIP_RAM.N_3_0 ));
    Odrv4 I__1662 (
            .O(N__8317),
            .I(\U712_CHIP_RAM.N_3_0 ));
    CascadeMux I__1661 (
            .O(N__8306),
            .I(N__8300));
    InMux I__1660 (
            .O(N__8305),
            .I(N__8296));
    CascadeMux I__1659 (
            .O(N__8304),
            .I(N__8291));
    InMux I__1658 (
            .O(N__8303),
            .I(N__8286));
    InMux I__1657 (
            .O(N__8300),
            .I(N__8286));
    InMux I__1656 (
            .O(N__8299),
            .I(N__8283));
    LocalMux I__1655 (
            .O(N__8296),
            .I(N__8280));
    InMux I__1654 (
            .O(N__8295),
            .I(N__8275));
    InMux I__1653 (
            .O(N__8294),
            .I(N__8275));
    InMux I__1652 (
            .O(N__8291),
            .I(N__8272));
    LocalMux I__1651 (
            .O(N__8286),
            .I(N__8269));
    LocalMux I__1650 (
            .O(N__8283),
            .I(N__8266));
    Span4Mux_h I__1649 (
            .O(N__8280),
            .I(N__8263));
    LocalMux I__1648 (
            .O(N__8275),
            .I(\U712_CHIP_RAM.m186_m2_0_a2_0 ));
    LocalMux I__1647 (
            .O(N__8272),
            .I(\U712_CHIP_RAM.m186_m2_0_a2_0 ));
    Odrv4 I__1646 (
            .O(N__8269),
            .I(\U712_CHIP_RAM.m186_m2_0_a2_0 ));
    Odrv4 I__1645 (
            .O(N__8266),
            .I(\U712_CHIP_RAM.m186_m2_0_a2_0 ));
    Odrv4 I__1644 (
            .O(N__8263),
            .I(\U712_CHIP_RAM.m186_m2_0_a2_0 ));
    CascadeMux I__1643 (
            .O(N__8252),
            .I(\U712_CHIP_RAM.m190_0_cascade_ ));
    InMux I__1642 (
            .O(N__8249),
            .I(N__8246));
    LocalMux I__1641 (
            .O(N__8246),
            .I(\U712_CHIP_RAM.m190_1 ));
    IoInMux I__1640 (
            .O(N__8243),
            .I(N__8240));
    LocalMux I__1639 (
            .O(N__8240),
            .I(N__8237));
    Span4Mux_s0_h I__1638 (
            .O(N__8237),
            .I(N__8234));
    Sp12to4 I__1637 (
            .O(N__8234),
            .I(N__8231));
    Span12Mux_v I__1636 (
            .O(N__8231),
            .I(N__8228));
    Span12Mux_h I__1635 (
            .O(N__8228),
            .I(N__8225));
    Odrv12 I__1634 (
            .O(N__8225),
            .I(CMA_c_6));
    InMux I__1633 (
            .O(N__8222),
            .I(N__8219));
    LocalMux I__1632 (
            .O(N__8219),
            .I(N__8216));
    Odrv4 I__1631 (
            .O(N__8216),
            .I(\U712_CHIP_RAM.d_N_6_3 ));
    CascadeMux I__1630 (
            .O(N__8213),
            .I(\U712_CHIP_RAM.N_208_cascade_ ));
    InMux I__1629 (
            .O(N__8210),
            .I(N__8206));
    InMux I__1628 (
            .O(N__8209),
            .I(N__8203));
    LocalMux I__1627 (
            .O(N__8206),
            .I(N__8199));
    LocalMux I__1626 (
            .O(N__8203),
            .I(N__8196));
    InMux I__1625 (
            .O(N__8202),
            .I(N__8193));
    Span4Mux_h I__1624 (
            .O(N__8199),
            .I(N__8190));
    Span4Mux_v I__1623 (
            .O(N__8196),
            .I(N__8187));
    LocalMux I__1622 (
            .O(N__8193),
            .I(N__8184));
    Odrv4 I__1621 (
            .O(N__8190),
            .I(N_99_0));
    Odrv4 I__1620 (
            .O(N__8187),
            .I(N_99_0));
    Odrv12 I__1619 (
            .O(N__8184),
            .I(N_99_0));
    IoInMux I__1618 (
            .O(N__8177),
            .I(N__8174));
    LocalMux I__1617 (
            .O(N__8174),
            .I(N__8171));
    Span12Mux_s5_v I__1616 (
            .O(N__8171),
            .I(N__8168));
    Span12Mux_h I__1615 (
            .O(N__8168),
            .I(N__8164));
    InMux I__1614 (
            .O(N__8167),
            .I(N__8161));
    Odrv12 I__1613 (
            .O(N__8164),
            .I(LDSn_c));
    LocalMux I__1612 (
            .O(N__8161),
            .I(LDSn_c));
    CascadeMux I__1611 (
            .O(N__8156),
            .I(N__8149));
    InMux I__1610 (
            .O(N__8155),
            .I(N__8145));
    InMux I__1609 (
            .O(N__8154),
            .I(N__8142));
    InMux I__1608 (
            .O(N__8153),
            .I(N__8135));
    InMux I__1607 (
            .O(N__8152),
            .I(N__8135));
    InMux I__1606 (
            .O(N__8149),
            .I(N__8135));
    CascadeMux I__1605 (
            .O(N__8148),
            .I(N__8132));
    LocalMux I__1604 (
            .O(N__8145),
            .I(N__8125));
    LocalMux I__1603 (
            .O(N__8142),
            .I(N__8125));
    LocalMux I__1602 (
            .O(N__8135),
            .I(N__8125));
    InMux I__1601 (
            .O(N__8132),
            .I(N__8122));
    Span4Mux_v I__1600 (
            .O(N__8125),
            .I(N__8119));
    LocalMux I__1599 (
            .O(N__8122),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    Odrv4 I__1598 (
            .O(N__8119),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    InMux I__1597 (
            .O(N__8114),
            .I(N__8101));
    InMux I__1596 (
            .O(N__8113),
            .I(N__8101));
    InMux I__1595 (
            .O(N__8112),
            .I(N__8101));
    InMux I__1594 (
            .O(N__8111),
            .I(N__8087));
    InMux I__1593 (
            .O(N__8110),
            .I(N__8087));
    InMux I__1592 (
            .O(N__8109),
            .I(N__8087));
    CascadeMux I__1591 (
            .O(N__8108),
            .I(N__8081));
    LocalMux I__1590 (
            .O(N__8101),
            .I(N__8077));
    InMux I__1589 (
            .O(N__8100),
            .I(N__8074));
    InMux I__1588 (
            .O(N__8099),
            .I(N__8065));
    InMux I__1587 (
            .O(N__8098),
            .I(N__8065));
    InMux I__1586 (
            .O(N__8097),
            .I(N__8065));
    InMux I__1585 (
            .O(N__8096),
            .I(N__8065));
    InMux I__1584 (
            .O(N__8095),
            .I(N__8062));
    InMux I__1583 (
            .O(N__8094),
            .I(N__8058));
    LocalMux I__1582 (
            .O(N__8087),
            .I(N__8053));
    InMux I__1581 (
            .O(N__8086),
            .I(N__8048));
    InMux I__1580 (
            .O(N__8085),
            .I(N__8048));
    InMux I__1579 (
            .O(N__8084),
            .I(N__8040));
    InMux I__1578 (
            .O(N__8081),
            .I(N__8040));
    InMux I__1577 (
            .O(N__8080),
            .I(N__8040));
    Span4Mux_v I__1576 (
            .O(N__8077),
            .I(N__8031));
    LocalMux I__1575 (
            .O(N__8074),
            .I(N__8031));
    LocalMux I__1574 (
            .O(N__8065),
            .I(N__8028));
    LocalMux I__1573 (
            .O(N__8062),
            .I(N__8025));
    InMux I__1572 (
            .O(N__8061),
            .I(N__8022));
    LocalMux I__1571 (
            .O(N__8058),
            .I(N__8019));
    InMux I__1570 (
            .O(N__8057),
            .I(N__8014));
    InMux I__1569 (
            .O(N__8056),
            .I(N__8014));
    Span4Mux_v I__1568 (
            .O(N__8053),
            .I(N__8009));
    LocalMux I__1567 (
            .O(N__8048),
            .I(N__8009));
    InMux I__1566 (
            .O(N__8047),
            .I(N__8006));
    LocalMux I__1565 (
            .O(N__8040),
            .I(N__8003));
    InMux I__1564 (
            .O(N__8039),
            .I(N__8000));
    InMux I__1563 (
            .O(N__8038),
            .I(N__7995));
    InMux I__1562 (
            .O(N__8037),
            .I(N__7995));
    InMux I__1561 (
            .O(N__8036),
            .I(N__7992));
    Span4Mux_v I__1560 (
            .O(N__8031),
            .I(N__7989));
    Span4Mux_v I__1559 (
            .O(N__8028),
            .I(N__7984));
    Span4Mux_v I__1558 (
            .O(N__8025),
            .I(N__7984));
    LocalMux I__1557 (
            .O(N__8022),
            .I(N__7981));
    Span4Mux_v I__1556 (
            .O(N__8019),
            .I(N__7976));
    LocalMux I__1555 (
            .O(N__8014),
            .I(N__7976));
    Span4Mux_h I__1554 (
            .O(N__8009),
            .I(N__7971));
    LocalMux I__1553 (
            .O(N__8006),
            .I(N__7971));
    Span4Mux_v I__1552 (
            .O(N__8003),
            .I(N__7964));
    LocalMux I__1551 (
            .O(N__8000),
            .I(N__7964));
    LocalMux I__1550 (
            .O(N__7995),
            .I(N__7964));
    LocalMux I__1549 (
            .O(N__7992),
            .I(N__7960));
    Span4Mux_h I__1548 (
            .O(N__7989),
            .I(N__7953));
    Span4Mux_h I__1547 (
            .O(N__7984),
            .I(N__7953));
    Span4Mux_v I__1546 (
            .O(N__7981),
            .I(N__7953));
    Span4Mux_v I__1545 (
            .O(N__7976),
            .I(N__7946));
    Span4Mux_v I__1544 (
            .O(N__7971),
            .I(N__7946));
    Span4Mux_v I__1543 (
            .O(N__7964),
            .I(N__7946));
    InMux I__1542 (
            .O(N__7963),
            .I(N__7943));
    Span12Mux_v I__1541 (
            .O(N__7960),
            .I(N__7936));
    Sp12to4 I__1540 (
            .O(N__7953),
            .I(N__7936));
    Sp12to4 I__1539 (
            .O(N__7946),
            .I(N__7936));
    LocalMux I__1538 (
            .O(N__7943),
            .I(N__7933));
    Span12Mux_h I__1537 (
            .O(N__7936),
            .I(N__7930));
    Span12Mux_h I__1536 (
            .O(N__7933),
            .I(N__7927));
    Odrv12 I__1535 (
            .O(N__7930),
            .I(RESETn_c));
    Odrv12 I__1534 (
            .O(N__7927),
            .I(RESETn_c));
    IoInMux I__1533 (
            .O(N__7922),
            .I(N__7919));
    LocalMux I__1532 (
            .O(N__7919),
            .I(N__7916));
    Span12Mux_s7_v I__1531 (
            .O(N__7916),
            .I(N__7913));
    Odrv12 I__1530 (
            .O(N__7913),
            .I(RESETn_c_i));
    IoInMux I__1529 (
            .O(N__7910),
            .I(N__7907));
    LocalMux I__1528 (
            .O(N__7907),
            .I(N__7904));
    Span4Mux_s3_v I__1527 (
            .O(N__7904),
            .I(N__7901));
    Span4Mux_v I__1526 (
            .O(N__7901),
            .I(N__7898));
    Span4Mux_h I__1525 (
            .O(N__7898),
            .I(N__7895));
    Odrv4 I__1524 (
            .O(N__7895),
            .I(RASn_c));
    InMux I__1523 (
            .O(N__7892),
            .I(N__7889));
    LocalMux I__1522 (
            .O(N__7889),
            .I(\U712_CHIP_RAM.d_N_7 ));
    InMux I__1521 (
            .O(N__7886),
            .I(N__7883));
    LocalMux I__1520 (
            .O(N__7883),
            .I(\U712_CHIP_RAM.m185_0 ));
    InMux I__1519 (
            .O(N__7880),
            .I(N__7877));
    LocalMux I__1518 (
            .O(N__7877),
            .I(N__7874));
    Sp12to4 I__1517 (
            .O(N__7874),
            .I(N__7871));
    Span12Mux_v I__1516 (
            .O(N__7871),
            .I(N__7868));
    Span12Mux_h I__1515 (
            .O(N__7868),
            .I(N__7865));
    Odrv12 I__1514 (
            .O(N__7865),
            .I(A_c_16));
    InMux I__1513 (
            .O(N__7862),
            .I(N__7858));
    InMux I__1512 (
            .O(N__7861),
            .I(N__7855));
    LocalMux I__1511 (
            .O(N__7858),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ));
    LocalMux I__1510 (
            .O(N__7855),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ));
    InMux I__1509 (
            .O(N__7850),
            .I(N__7844));
    InMux I__1508 (
            .O(N__7849),
            .I(N__7844));
    LocalMux I__1507 (
            .O(N__7844),
            .I(N__7841));
    Span4Mux_v I__1506 (
            .O(N__7841),
            .I(N__7837));
    InMux I__1505 (
            .O(N__7840),
            .I(N__7834));
    Sp12to4 I__1504 (
            .O(N__7837),
            .I(N__7829));
    LocalMux I__1503 (
            .O(N__7834),
            .I(N__7829));
    Span12Mux_h I__1502 (
            .O(N__7829),
            .I(N__7826));
    Odrv12 I__1501 (
            .O(N__7826),
            .I(AWEn_c));
    CascadeMux I__1500 (
            .O(N__7823),
            .I(N__7820));
    InMux I__1499 (
            .O(N__7820),
            .I(N__7817));
    LocalMux I__1498 (
            .O(N__7817),
            .I(N__7813));
    CascadeMux I__1497 (
            .O(N__7816),
            .I(N__7810));
    Span4Mux_v I__1496 (
            .O(N__7813),
            .I(N__7806));
    InMux I__1495 (
            .O(N__7810),
            .I(N__7803));
    InMux I__1494 (
            .O(N__7809),
            .I(N__7796));
    Sp12to4 I__1493 (
            .O(N__7806),
            .I(N__7791));
    LocalMux I__1492 (
            .O(N__7803),
            .I(N__7791));
    InMux I__1491 (
            .O(N__7802),
            .I(N__7786));
    InMux I__1490 (
            .O(N__7801),
            .I(N__7786));
    InMux I__1489 (
            .O(N__7800),
            .I(N__7781));
    InMux I__1488 (
            .O(N__7799),
            .I(N__7781));
    LocalMux I__1487 (
            .O(N__7796),
            .I(\U712_CHIP_RAM.N_26_0 ));
    Odrv12 I__1486 (
            .O(N__7791),
            .I(\U712_CHIP_RAM.N_26_0 ));
    LocalMux I__1485 (
            .O(N__7786),
            .I(\U712_CHIP_RAM.N_26_0 ));
    LocalMux I__1484 (
            .O(N__7781),
            .I(\U712_CHIP_RAM.N_26_0 ));
    CascadeMux I__1483 (
            .O(N__7772),
            .I(N__7767));
    InMux I__1482 (
            .O(N__7771),
            .I(N__7763));
    InMux I__1481 (
            .O(N__7770),
            .I(N__7760));
    InMux I__1480 (
            .O(N__7767),
            .I(N__7757));
    CascadeMux I__1479 (
            .O(N__7766),
            .I(N__7753));
    LocalMux I__1478 (
            .O(N__7763),
            .I(N__7741));
    LocalMux I__1477 (
            .O(N__7760),
            .I(N__7741));
    LocalMux I__1476 (
            .O(N__7757),
            .I(N__7738));
    InMux I__1475 (
            .O(N__7756),
            .I(N__7727));
    InMux I__1474 (
            .O(N__7753),
            .I(N__7727));
    InMux I__1473 (
            .O(N__7752),
            .I(N__7727));
    InMux I__1472 (
            .O(N__7751),
            .I(N__7727));
    InMux I__1471 (
            .O(N__7750),
            .I(N__7727));
    InMux I__1470 (
            .O(N__7749),
            .I(N__7721));
    InMux I__1469 (
            .O(N__7748),
            .I(N__7718));
    InMux I__1468 (
            .O(N__7747),
            .I(N__7713));
    InMux I__1467 (
            .O(N__7746),
            .I(N__7713));
    Span4Mux_h I__1466 (
            .O(N__7741),
            .I(N__7710));
    Span4Mux_h I__1465 (
            .O(N__7738),
            .I(N__7705));
    LocalMux I__1464 (
            .O(N__7727),
            .I(N__7705));
    InMux I__1463 (
            .O(N__7726),
            .I(N__7698));
    InMux I__1462 (
            .O(N__7725),
            .I(N__7698));
    InMux I__1461 (
            .O(N__7724),
            .I(N__7698));
    LocalMux I__1460 (
            .O(N__7721),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1459 (
            .O(N__7718),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1458 (
            .O(N__7713),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1457 (
            .O(N__7710),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1456 (
            .O(N__7705),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1455 (
            .O(N__7698),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    CascadeMux I__1454 (
            .O(N__7685),
            .I(N__7682));
    InMux I__1453 (
            .O(N__7682),
            .I(N__7676));
    InMux I__1452 (
            .O(N__7681),
            .I(N__7673));
    InMux I__1451 (
            .O(N__7680),
            .I(N__7670));
    InMux I__1450 (
            .O(N__7679),
            .I(N__7667));
    LocalMux I__1449 (
            .O(N__7676),
            .I(N__7663));
    LocalMux I__1448 (
            .O(N__7673),
            .I(N__7660));
    LocalMux I__1447 (
            .O(N__7670),
            .I(N__7655));
    LocalMux I__1446 (
            .O(N__7667),
            .I(N__7655));
    InMux I__1445 (
            .O(N__7666),
            .I(N__7652));
    Odrv12 I__1444 (
            .O(N__7663),
            .I(\U712_CHIP_RAM.N_30_0 ));
    Odrv4 I__1443 (
            .O(N__7660),
            .I(\U712_CHIP_RAM.N_30_0 ));
    Odrv4 I__1442 (
            .O(N__7655),
            .I(\U712_CHIP_RAM.N_30_0 ));
    LocalMux I__1441 (
            .O(N__7652),
            .I(\U712_CHIP_RAM.N_30_0 ));
    CascadeMux I__1440 (
            .O(N__7643),
            .I(\U712_CHIP_RAM.N_62_0_cascade_ ));
    InMux I__1439 (
            .O(N__7640),
            .I(N__7637));
    LocalMux I__1438 (
            .O(N__7637),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_RNI9THUZ0Z5 ));
    CascadeMux I__1437 (
            .O(N__7634),
            .I(\U712_CHIP_RAM.CLK_EN_RNOZ0Z_2_cascade_ ));
    InMux I__1436 (
            .O(N__7631),
            .I(N__7628));
    LocalMux I__1435 (
            .O(N__7628),
            .I(N__7625));
    Odrv4 I__1434 (
            .O(N__7625),
            .I(\U712_CHIP_RAM.CLK_EN_RNOZ0Z_3 ));
    CascadeMux I__1433 (
            .O(N__7622),
            .I(\U712_CHIP_RAM.N_174_0_cascade_ ));
    InMux I__1432 (
            .O(N__7619),
            .I(N__7616));
    LocalMux I__1431 (
            .O(N__7616),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER43 ));
    IoInMux I__1430 (
            .O(N__7613),
            .I(N__7610));
    LocalMux I__1429 (
            .O(N__7610),
            .I(N__7607));
    Span4Mux_s1_h I__1428 (
            .O(N__7607),
            .I(N__7604));
    Sp12to4 I__1427 (
            .O(N__7604),
            .I(N__7601));
    Span12Mux_v I__1426 (
            .O(N__7601),
            .I(N__7598));
    Span12Mux_h I__1425 (
            .O(N__7598),
            .I(N__7594));
    InMux I__1424 (
            .O(N__7597),
            .I(N__7591));
    Odrv12 I__1423 (
            .O(N__7594),
            .I(CLK_EN_c));
    LocalMux I__1422 (
            .O(N__7591),
            .I(CLK_EN_c));
    CascadeMux I__1421 (
            .O(N__7586),
            .I(N__7583));
    InMux I__1420 (
            .O(N__7583),
            .I(N__7575));
    InMux I__1419 (
            .O(N__7582),
            .I(N__7568));
    InMux I__1418 (
            .O(N__7581),
            .I(N__7568));
    InMux I__1417 (
            .O(N__7580),
            .I(N__7568));
    CascadeMux I__1416 (
            .O(N__7579),
            .I(N__7565));
    CascadeMux I__1415 (
            .O(N__7578),
            .I(N__7561));
    LocalMux I__1414 (
            .O(N__7575),
            .I(N__7558));
    LocalMux I__1413 (
            .O(N__7568),
            .I(N__7555));
    InMux I__1412 (
            .O(N__7565),
            .I(N__7552));
    InMux I__1411 (
            .O(N__7564),
            .I(N__7549));
    InMux I__1410 (
            .O(N__7561),
            .I(N__7546));
    Span4Mux_v I__1409 (
            .O(N__7558),
            .I(N__7543));
    Span4Mux_v I__1408 (
            .O(N__7555),
            .I(N__7538));
    LocalMux I__1407 (
            .O(N__7552),
            .I(N__7538));
    LocalMux I__1406 (
            .O(N__7549),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    LocalMux I__1405 (
            .O(N__7546),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    Odrv4 I__1404 (
            .O(N__7543),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    Odrv4 I__1403 (
            .O(N__7538),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    CascadeMux I__1402 (
            .O(N__7529),
            .I(N__7525));
    CascadeMux I__1401 (
            .O(N__7528),
            .I(N__7521));
    InMux I__1400 (
            .O(N__7525),
            .I(N__7518));
    InMux I__1399 (
            .O(N__7524),
            .I(N__7515));
    InMux I__1398 (
            .O(N__7521),
            .I(N__7512));
    LocalMux I__1397 (
            .O(N__7518),
            .I(\U712_CHIP_RAM.N_62_0 ));
    LocalMux I__1396 (
            .O(N__7515),
            .I(\U712_CHIP_RAM.N_62_0 ));
    LocalMux I__1395 (
            .O(N__7512),
            .I(\U712_CHIP_RAM.N_62_0 ));
    InMux I__1394 (
            .O(N__7505),
            .I(N__7500));
    InMux I__1393 (
            .O(N__7504),
            .I(N__7494));
    InMux I__1392 (
            .O(N__7503),
            .I(N__7494));
    LocalMux I__1391 (
            .O(N__7500),
            .I(N__7491));
    InMux I__1390 (
            .O(N__7499),
            .I(N__7488));
    LocalMux I__1389 (
            .O(N__7494),
            .I(\U712_CHIP_RAM.N_52_0 ));
    Odrv4 I__1388 (
            .O(N__7491),
            .I(\U712_CHIP_RAM.N_52_0 ));
    LocalMux I__1387 (
            .O(N__7488),
            .I(\U712_CHIP_RAM.N_52_0 ));
    InMux I__1386 (
            .O(N__7481),
            .I(N__7478));
    LocalMux I__1385 (
            .O(N__7478),
            .I(N__7475));
    Span4Mux_v I__1384 (
            .O(N__7475),
            .I(N__7472));
    Sp12to4 I__1383 (
            .O(N__7472),
            .I(N__7469));
    Span12Mux_h I__1382 (
            .O(N__7469),
            .I(N__7466));
    Odrv12 I__1381 (
            .O(N__7466),
            .I(A_c_4));
    CascadeMux I__1380 (
            .O(N__7463),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_ ));
    InMux I__1379 (
            .O(N__7460),
            .I(N__7456));
    InMux I__1378 (
            .O(N__7459),
            .I(N__7453));
    LocalMux I__1377 (
            .O(N__7456),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ));
    LocalMux I__1376 (
            .O(N__7453),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ));
    InMux I__1375 (
            .O(N__7448),
            .I(N__7445));
    LocalMux I__1374 (
            .O(N__7445),
            .I(N__7442));
    Span4Mux_v I__1373 (
            .O(N__7442),
            .I(N__7439));
    Sp12to4 I__1372 (
            .O(N__7439),
            .I(N__7436));
    Span12Mux_h I__1371 (
            .O(N__7436),
            .I(N__7433));
    Odrv12 I__1370 (
            .O(N__7433),
            .I(A_c_5));
    InMux I__1369 (
            .O(N__7430),
            .I(N__7426));
    InMux I__1368 (
            .O(N__7429),
            .I(N__7423));
    LocalMux I__1367 (
            .O(N__7426),
            .I(N__7420));
    LocalMux I__1366 (
            .O(N__7423),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ));
    Odrv12 I__1365 (
            .O(N__7420),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ));
    InMux I__1364 (
            .O(N__7415),
            .I(N__7412));
    LocalMux I__1363 (
            .O(N__7412),
            .I(N__7409));
    Span4Mux_v I__1362 (
            .O(N__7409),
            .I(N__7406));
    Sp12to4 I__1361 (
            .O(N__7406),
            .I(N__7403));
    Span12Mux_h I__1360 (
            .O(N__7403),
            .I(N__7400));
    Odrv12 I__1359 (
            .O(N__7400),
            .I(A_c_6));
    InMux I__1358 (
            .O(N__7397),
            .I(N__7394));
    LocalMux I__1357 (
            .O(N__7394),
            .I(N__7390));
    InMux I__1356 (
            .O(N__7393),
            .I(N__7387));
    Span4Mux_v I__1355 (
            .O(N__7390),
            .I(N__7384));
    LocalMux I__1354 (
            .O(N__7387),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ));
    Odrv4 I__1353 (
            .O(N__7384),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ));
    InMux I__1352 (
            .O(N__7379),
            .I(N__7376));
    LocalMux I__1351 (
            .O(N__7376),
            .I(N__7373));
    Span12Mux_v I__1350 (
            .O(N__7373),
            .I(N__7370));
    Span12Mux_h I__1349 (
            .O(N__7370),
            .I(N__7367));
    Odrv12 I__1348 (
            .O(N__7367),
            .I(A_c_7));
    InMux I__1347 (
            .O(N__7364),
            .I(N__7361));
    LocalMux I__1346 (
            .O(N__7361),
            .I(N__7357));
    InMux I__1345 (
            .O(N__7360),
            .I(N__7354));
    Span4Mux_v I__1344 (
            .O(N__7357),
            .I(N__7351));
    LocalMux I__1343 (
            .O(N__7354),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ));
    Odrv4 I__1342 (
            .O(N__7351),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ));
    CascadeMux I__1341 (
            .O(N__7346),
            .I(\U712_CHIP_RAM.DMA_CYCLE_START_RNIJD6OZ0Z3_cascade_ ));
    CascadeMux I__1340 (
            .O(N__7343),
            .I(\U712_CHIP_RAM.N_204_cascade_ ));
    InMux I__1339 (
            .O(N__7340),
            .I(N__7337));
    LocalMux I__1338 (
            .O(N__7337),
            .I(N__7332));
    InMux I__1337 (
            .O(N__7336),
            .I(N__7329));
    InMux I__1336 (
            .O(N__7335),
            .I(N__7326));
    Span4Mux_v I__1335 (
            .O(N__7332),
            .I(N__7320));
    LocalMux I__1334 (
            .O(N__7329),
            .I(N__7320));
    LocalMux I__1333 (
            .O(N__7326),
            .I(N__7317));
    InMux I__1332 (
            .O(N__7325),
            .I(N__7314));
    Span4Mux_h I__1331 (
            .O(N__7320),
            .I(N__7311));
    Odrv4 I__1330 (
            .O(N__7317),
            .I(\U712_CHIP_RAM.N_364 ));
    LocalMux I__1329 (
            .O(N__7314),
            .I(\U712_CHIP_RAM.N_364 ));
    Odrv4 I__1328 (
            .O(N__7311),
            .I(\U712_CHIP_RAM.N_364 ));
    InMux I__1327 (
            .O(N__7304),
            .I(N__7300));
    InMux I__1326 (
            .O(N__7303),
            .I(N__7294));
    LocalMux I__1325 (
            .O(N__7300),
            .I(N__7291));
    InMux I__1324 (
            .O(N__7299),
            .I(N__7286));
    InMux I__1323 (
            .O(N__7298),
            .I(N__7286));
    InMux I__1322 (
            .O(N__7297),
            .I(N__7283));
    LocalMux I__1321 (
            .O(N__7294),
            .I(N__7276));
    Span4Mux_v I__1320 (
            .O(N__7291),
            .I(N__7273));
    LocalMux I__1319 (
            .O(N__7286),
            .I(N__7268));
    LocalMux I__1318 (
            .O(N__7283),
            .I(N__7268));
    InMux I__1317 (
            .O(N__7282),
            .I(N__7265));
    InMux I__1316 (
            .O(N__7281),
            .I(N__7262));
    InMux I__1315 (
            .O(N__7280),
            .I(N__7257));
    InMux I__1314 (
            .O(N__7279),
            .I(N__7257));
    Span4Mux_h I__1313 (
            .O(N__7276),
            .I(N__7254));
    Span4Mux_h I__1312 (
            .O(N__7273),
            .I(N__7249));
    Span4Mux_h I__1311 (
            .O(N__7268),
            .I(N__7249));
    LocalMux I__1310 (
            .O(N__7265),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1309 (
            .O(N__7262),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1308 (
            .O(N__7257),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1307 (
            .O(N__7254),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1306 (
            .O(N__7249),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    CascadeMux I__1305 (
            .O(N__7238),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_ ));
    IoInMux I__1304 (
            .O(N__7235),
            .I(N__7232));
    LocalMux I__1303 (
            .O(N__7232),
            .I(N__7229));
    Span4Mux_s2_v I__1302 (
            .O(N__7229),
            .I(N__7226));
    Span4Mux_v I__1301 (
            .O(N__7226),
            .I(N__7223));
    Span4Mux_h I__1300 (
            .O(N__7223),
            .I(N__7220));
    Sp12to4 I__1299 (
            .O(N__7220),
            .I(N__7217));
    Span12Mux_v I__1298 (
            .O(N__7217),
            .I(N__7213));
    InMux I__1297 (
            .O(N__7216),
            .I(N__7210));
    Odrv12 I__1296 (
            .O(N__7213),
            .I(DBDIR_c));
    LocalMux I__1295 (
            .O(N__7210),
            .I(DBDIR_c));
    IoInMux I__1294 (
            .O(N__7205),
            .I(N__7202));
    LocalMux I__1293 (
            .O(N__7202),
            .I(N__7199));
    IoSpan4Mux I__1292 (
            .O(N__7199),
            .I(N__7196));
    Span4Mux_s2_v I__1291 (
            .O(N__7196),
            .I(N__7193));
    Sp12to4 I__1290 (
            .O(N__7193),
            .I(N__7189));
    InMux I__1289 (
            .O(N__7192),
            .I(N__7186));
    Span12Mux_s8_v I__1288 (
            .O(N__7189),
            .I(N__7183));
    LocalMux I__1287 (
            .O(N__7186),
            .I(N__7180));
    Span12Mux_v I__1286 (
            .O(N__7183),
            .I(N__7177));
    Span12Mux_v I__1285 (
            .O(N__7180),
            .I(N__7174));
    Span12Mux_h I__1284 (
            .O(N__7177),
            .I(N__7171));
    Span12Mux_h I__1283 (
            .O(N__7174),
            .I(N__7168));
    Odrv12 I__1282 (
            .O(N__7171),
            .I(A_c_11));
    Odrv12 I__1281 (
            .O(N__7168),
            .I(A_c_11));
    CascadeMux I__1280 (
            .O(N__7163),
            .I(\U712_CHIP_RAM.N_3_0_cascade_ ));
    InMux I__1279 (
            .O(N__7160),
            .I(N__7157));
    LocalMux I__1278 (
            .O(N__7157),
            .I(\U712_CHIP_RAM.m187_0 ));
    InMux I__1277 (
            .O(N__7154),
            .I(N__7151));
    LocalMux I__1276 (
            .O(N__7151),
            .I(N__7148));
    Span4Mux_h I__1275 (
            .O(N__7148),
            .I(N__7145));
    Odrv4 I__1274 (
            .O(N__7145),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_1 ));
    CascadeMux I__1273 (
            .O(N__7142),
            .I(\U712_CHIP_RAM.N_163_0_cascade_ ));
    InMux I__1272 (
            .O(N__7139),
            .I(N__7133));
    InMux I__1271 (
            .O(N__7138),
            .I(N__7130));
    InMux I__1270 (
            .O(N__7137),
            .I(N__7125));
    InMux I__1269 (
            .O(N__7136),
            .I(N__7125));
    LocalMux I__1268 (
            .O(N__7133),
            .I(\U712_CHIP_RAM.N_67_0 ));
    LocalMux I__1267 (
            .O(N__7130),
            .I(\U712_CHIP_RAM.N_67_0 ));
    LocalMux I__1266 (
            .O(N__7125),
            .I(\U712_CHIP_RAM.N_67_0 ));
    SRMux I__1265 (
            .O(N__7118),
            .I(N__7115));
    LocalMux I__1264 (
            .O(N__7115),
            .I(N__7112));
    Span4Mux_v I__1263 (
            .O(N__7112),
            .I(N__7109));
    Span4Mux_h I__1262 (
            .O(N__7109),
            .I(N__7106));
    Odrv4 I__1261 (
            .O(N__7106),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    InMux I__1260 (
            .O(N__7103),
            .I(N__7100));
    LocalMux I__1259 (
            .O(N__7100),
            .I(N__7097));
    Span4Mux_h I__1258 (
            .O(N__7097),
            .I(N__7090));
    InMux I__1257 (
            .O(N__7096),
            .I(N__7087));
    InMux I__1256 (
            .O(N__7095),
            .I(N__7084));
    InMux I__1255 (
            .O(N__7094),
            .I(N__7079));
    InMux I__1254 (
            .O(N__7093),
            .I(N__7079));
    Odrv4 I__1253 (
            .O(N__7090),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__1252 (
            .O(N__7087),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__1251 (
            .O(N__7084),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__1250 (
            .O(N__7079),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    InMux I__1249 (
            .O(N__7070),
            .I(N__7064));
    InMux I__1248 (
            .O(N__7069),
            .I(N__7061));
    InMux I__1247 (
            .O(N__7068),
            .I(N__7056));
    InMux I__1246 (
            .O(N__7067),
            .I(N__7056));
    LocalMux I__1245 (
            .O(N__7064),
            .I(N__7051));
    LocalMux I__1244 (
            .O(N__7061),
            .I(N__7051));
    LocalMux I__1243 (
            .O(N__7056),
            .I(\U712_CHIP_RAM.N_48_0 ));
    Odrv4 I__1242 (
            .O(N__7051),
            .I(\U712_CHIP_RAM.N_48_0 ));
    InMux I__1241 (
            .O(N__7046),
            .I(N__7043));
    LocalMux I__1240 (
            .O(N__7043),
            .I(N__7039));
    InMux I__1239 (
            .O(N__7042),
            .I(N__7036));
    Span4Mux_h I__1238 (
            .O(N__7039),
            .I(N__7033));
    LocalMux I__1237 (
            .O(N__7036),
            .I(\U712_CHIP_RAM.N_363 ));
    Odrv4 I__1236 (
            .O(N__7033),
            .I(\U712_CHIP_RAM.N_363 ));
    CascadeMux I__1235 (
            .O(N__7028),
            .I(\U712_CHIP_RAM.N_158_0_cascade_ ));
    InMux I__1234 (
            .O(N__7025),
            .I(N__7019));
    InMux I__1233 (
            .O(N__7024),
            .I(N__7010));
    InMux I__1232 (
            .O(N__7023),
            .I(N__7010));
    InMux I__1231 (
            .O(N__7022),
            .I(N__7010));
    LocalMux I__1230 (
            .O(N__7019),
            .I(N__7007));
    InMux I__1229 (
            .O(N__7018),
            .I(N__7002));
    InMux I__1228 (
            .O(N__7017),
            .I(N__7002));
    LocalMux I__1227 (
            .O(N__7010),
            .I(\U712_CHIP_RAM.N_58_0 ));
    Odrv4 I__1226 (
            .O(N__7007),
            .I(\U712_CHIP_RAM.N_58_0 ));
    LocalMux I__1225 (
            .O(N__7002),
            .I(\U712_CHIP_RAM.N_58_0 ));
    InMux I__1224 (
            .O(N__6995),
            .I(N__6992));
    LocalMux I__1223 (
            .O(N__6992),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_1 ));
    InMux I__1222 (
            .O(N__6989),
            .I(N__6986));
    LocalMux I__1221 (
            .O(N__6986),
            .I(N__6983));
    Odrv4 I__1220 (
            .O(N__6983),
            .I(\U712_CHIP_RAM.d_N_6_0 ));
    InMux I__1219 (
            .O(N__6980),
            .I(N__6977));
    LocalMux I__1218 (
            .O(N__6977),
            .I(N__6972));
    InMux I__1217 (
            .O(N__6976),
            .I(N__6969));
    InMux I__1216 (
            .O(N__6975),
            .I(N__6966));
    Odrv4 I__1215 (
            .O(N__6972),
            .I(\U712_CHIP_RAM.N_43_0 ));
    LocalMux I__1214 (
            .O(N__6969),
            .I(\U712_CHIP_RAM.N_43_0 ));
    LocalMux I__1213 (
            .O(N__6966),
            .I(\U712_CHIP_RAM.N_43_0 ));
    CascadeMux I__1212 (
            .O(N__6959),
            .I(N__6956));
    InMux I__1211 (
            .O(N__6956),
            .I(N__6953));
    LocalMux I__1210 (
            .O(N__6953),
            .I(\U712_CHIP_RAM.m189_0 ));
    InMux I__1209 (
            .O(N__6950),
            .I(N__6947));
    LocalMux I__1208 (
            .O(N__6947),
            .I(N__6944));
    Span4Mux_h I__1207 (
            .O(N__6944),
            .I(N__6941));
    Sp12to4 I__1206 (
            .O(N__6941),
            .I(N__6938));
    Span12Mux_v I__1205 (
            .O(N__6938),
            .I(N__6935));
    Span12Mux_h I__1204 (
            .O(N__6935),
            .I(N__6932));
    Odrv12 I__1203 (
            .O(N__6932),
            .I(A_c_14));
    IoInMux I__1202 (
            .O(N__6929),
            .I(N__6926));
    LocalMux I__1201 (
            .O(N__6926),
            .I(N__6923));
    IoSpan4Mux I__1200 (
            .O(N__6923),
            .I(N__6920));
    Span4Mux_s0_v I__1199 (
            .O(N__6920),
            .I(N__6917));
    Sp12to4 I__1198 (
            .O(N__6917),
            .I(N__6914));
    Odrv12 I__1197 (
            .O(N__6914),
            .I(CMA_c_2));
    InMux I__1196 (
            .O(N__6911),
            .I(N__6908));
    LocalMux I__1195 (
            .O(N__6908),
            .I(\U712_CHIP_RAM.m186_1 ));
    IoInMux I__1194 (
            .O(N__6905),
            .I(N__6902));
    LocalMux I__1193 (
            .O(N__6902),
            .I(N__6899));
    Span4Mux_s1_v I__1192 (
            .O(N__6899),
            .I(N__6896));
    Span4Mux_v I__1191 (
            .O(N__6896),
            .I(N__6893));
    Sp12to4 I__1190 (
            .O(N__6893),
            .I(N__6890));
    Span12Mux_h I__1189 (
            .O(N__6890),
            .I(N__6887));
    Odrv12 I__1188 (
            .O(N__6887),
            .I(CMA_c_0));
    IoInMux I__1187 (
            .O(N__6884),
            .I(N__6881));
    LocalMux I__1186 (
            .O(N__6881),
            .I(N__6878));
    Span12Mux_s7_v I__1185 (
            .O(N__6878),
            .I(N__6875));
    Odrv12 I__1184 (
            .O(N__6875),
            .I(CMA_c_1));
    CascadeMux I__1183 (
            .O(N__6872),
            .I(\U712_CHIP_RAM.N_198_cascade_ ));
    ClkMux I__1182 (
            .O(N__6869),
            .I(N__6864));
    InMux I__1181 (
            .O(N__6868),
            .I(N__6861));
    ClkMux I__1180 (
            .O(N__6867),
            .I(N__6858));
    LocalMux I__1179 (
            .O(N__6864),
            .I(N__6855));
    LocalMux I__1178 (
            .O(N__6861),
            .I(N__6852));
    LocalMux I__1177 (
            .O(N__6858),
            .I(N__6849));
    Span4Mux_h I__1176 (
            .O(N__6855),
            .I(N__6842));
    Span4Mux_v I__1175 (
            .O(N__6852),
            .I(N__6842));
    Span4Mux_h I__1174 (
            .O(N__6849),
            .I(N__6842));
    Span4Mux_v I__1173 (
            .O(N__6842),
            .I(N__6839));
    Span4Mux_v I__1172 (
            .O(N__6839),
            .I(N__6836));
    Odrv4 I__1171 (
            .O(N__6836),
            .I(CLK40_PLL));
    IoInMux I__1170 (
            .O(N__6833),
            .I(N__6828));
    IoInMux I__1169 (
            .O(N__6832),
            .I(N__6825));
    IoInMux I__1168 (
            .O(N__6831),
            .I(N__6822));
    LocalMux I__1167 (
            .O(N__6828),
            .I(N__6819));
    LocalMux I__1166 (
            .O(N__6825),
            .I(N__6816));
    LocalMux I__1165 (
            .O(N__6822),
            .I(N__6813));
    IoSpan4Mux I__1164 (
            .O(N__6819),
            .I(N__6810));
    IoSpan4Mux I__1163 (
            .O(N__6816),
            .I(N__6807));
    Span12Mux_s6_v I__1162 (
            .O(N__6813),
            .I(N__6804));
    Sp12to4 I__1161 (
            .O(N__6810),
            .I(N__6801));
    Span4Mux_s2_h I__1160 (
            .O(N__6807),
            .I(N__6798));
    Span12Mux_v I__1159 (
            .O(N__6804),
            .I(N__6795));
    Span12Mux_s6_v I__1158 (
            .O(N__6801),
            .I(N__6792));
    Sp12to4 I__1157 (
            .O(N__6798),
            .I(N__6789));
    Span12Mux_h I__1156 (
            .O(N__6795),
            .I(N__6786));
    Span12Mux_v I__1155 (
            .O(N__6792),
            .I(N__6781));
    Span12Mux_h I__1154 (
            .O(N__6789),
            .I(N__6781));
    Odrv12 I__1153 (
            .O(N__6786),
            .I(CLK40_PLL_iso_i));
    Odrv12 I__1152 (
            .O(N__6781),
            .I(CLK40_PLL_iso_i));
    InMux I__1151 (
            .O(N__6776),
            .I(N__6773));
    LocalMux I__1150 (
            .O(N__6773),
            .I(\U712_CHIP_RAM.m187_1 ));
    IoInMux I__1149 (
            .O(N__6770),
            .I(N__6767));
    LocalMux I__1148 (
            .O(N__6767),
            .I(N__6764));
    IoSpan4Mux I__1147 (
            .O(N__6764),
            .I(N__6761));
    Span4Mux_s3_h I__1146 (
            .O(N__6761),
            .I(N__6758));
    Span4Mux_v I__1145 (
            .O(N__6758),
            .I(N__6755));
    Span4Mux_h I__1144 (
            .O(N__6755),
            .I(N__6752));
    Sp12to4 I__1143 (
            .O(N__6752),
            .I(N__6749));
    Odrv12 I__1142 (
            .O(N__6749),
            .I(CMA_c_4));
    IoInMux I__1141 (
            .O(N__6746),
            .I(N__6743));
    LocalMux I__1140 (
            .O(N__6743),
            .I(N__6740));
    Span4Mux_s3_h I__1139 (
            .O(N__6740),
            .I(N__6737));
    Span4Mux_v I__1138 (
            .O(N__6737),
            .I(N__6734));
    Span4Mux_h I__1137 (
            .O(N__6734),
            .I(N__6731));
    Span4Mux_h I__1136 (
            .O(N__6731),
            .I(N__6728));
    Span4Mux_h I__1135 (
            .O(N__6728),
            .I(N__6725));
    Odrv4 I__1134 (
            .O(N__6725),
            .I(CMA_c_3));
    IoInMux I__1133 (
            .O(N__6722),
            .I(N__6719));
    LocalMux I__1132 (
            .O(N__6719),
            .I(N__6716));
    Span4Mux_s2_v I__1131 (
            .O(N__6716),
            .I(N__6713));
    Sp12to4 I__1130 (
            .O(N__6713),
            .I(N__6710));
    Span12Mux_h I__1129 (
            .O(N__6710),
            .I(N__6707));
    Odrv12 I__1128 (
            .O(N__6707),
            .I(CMA_c_10));
    InMux I__1127 (
            .O(N__6704),
            .I(N__6701));
    LocalMux I__1126 (
            .O(N__6701),
            .I(\U712_CHIP_RAM.m189_1 ));
    InMux I__1125 (
            .O(N__6698),
            .I(N__6695));
    LocalMux I__1124 (
            .O(N__6695),
            .I(\U712_CHIP_RAM.m188_1 ));
    InMux I__1123 (
            .O(N__6692),
            .I(N__6689));
    LocalMux I__1122 (
            .O(N__6689),
            .I(\U712_CHIP_RAM.d_N_6_2 ));
    InMux I__1121 (
            .O(N__6686),
            .I(N__6683));
    LocalMux I__1120 (
            .O(N__6683),
            .I(N__6680));
    Span4Mux_v I__1119 (
            .O(N__6680),
            .I(N__6677));
    Sp12to4 I__1118 (
            .O(N__6677),
            .I(N__6674));
    Span12Mux_h I__1117 (
            .O(N__6674),
            .I(N__6671));
    Odrv12 I__1116 (
            .O(N__6671),
            .I(A_c_12));
    InMux I__1115 (
            .O(N__6668),
            .I(N__6665));
    LocalMux I__1114 (
            .O(N__6665),
            .I(\U712_CHIP_RAM.m188_0 ));
    InMux I__1113 (
            .O(N__6662),
            .I(N__6659));
    LocalMux I__1112 (
            .O(N__6659),
            .I(\U712_CHIP_RAM.d_N_6 ));
    InMux I__1111 (
            .O(N__6656),
            .I(N__6653));
    LocalMux I__1110 (
            .O(N__6653),
            .I(N__6650));
    Span12Mux_v I__1109 (
            .O(N__6650),
            .I(N__6647));
    Span12Mux_h I__1108 (
            .O(N__6647),
            .I(N__6644));
    Odrv12 I__1107 (
            .O(N__6644),
            .I(A_c_13));
    InMux I__1106 (
            .O(N__6641),
            .I(N__6638));
    LocalMux I__1105 (
            .O(N__6638),
            .I(\U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0 ));
    InMux I__1104 (
            .O(N__6635),
            .I(N__6632));
    LocalMux I__1103 (
            .O(N__6632),
            .I(\U712_CHIP_RAM.N_213 ));
    InMux I__1102 (
            .O(N__6629),
            .I(N__6626));
    LocalMux I__1101 (
            .O(N__6626),
            .I(N__6623));
    Span4Mux_v I__1100 (
            .O(N__6623),
            .I(N__6619));
    InMux I__1099 (
            .O(N__6622),
            .I(N__6616));
    Odrv4 I__1098 (
            .O(N__6619),
            .I(CPU_TACKm));
    LocalMux I__1097 (
            .O(N__6616),
            .I(CPU_TACKm));
    InMux I__1096 (
            .O(N__6611),
            .I(N__6607));
    InMux I__1095 (
            .O(N__6610),
            .I(N__6604));
    LocalMux I__1094 (
            .O(N__6607),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__1093 (
            .O(N__6604),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__1092 (
            .O(N__6599),
            .I(N__6595));
    InMux I__1091 (
            .O(N__6598),
            .I(N__6592));
    LocalMux I__1090 (
            .O(N__6595),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__1089 (
            .O(N__6592),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__1088 (
            .O(N__6587),
            .I(N__6583));
    InMux I__1087 (
            .O(N__6586),
            .I(N__6580));
    InMux I__1086 (
            .O(N__6583),
            .I(N__6577));
    LocalMux I__1085 (
            .O(N__6580),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1084 (
            .O(N__6577),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__1083 (
            .O(N__6572),
            .I(N__6568));
    InMux I__1082 (
            .O(N__6571),
            .I(N__6565));
    LocalMux I__1081 (
            .O(N__6568),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__1080 (
            .O(N__6565),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    CascadeMux I__1079 (
            .O(N__6560),
            .I(\U712_CHIP_RAM.N_333_mux_cascade_ ));
    InMux I__1078 (
            .O(N__6557),
            .I(N__6551));
    InMux I__1077 (
            .O(N__6556),
            .I(N__6546));
    InMux I__1076 (
            .O(N__6555),
            .I(N__6546));
    InMux I__1075 (
            .O(N__6554),
            .I(N__6541));
    LocalMux I__1074 (
            .O(N__6551),
            .I(N__6538));
    LocalMux I__1073 (
            .O(N__6546),
            .I(N__6535));
    InMux I__1072 (
            .O(N__6545),
            .I(N__6530));
    InMux I__1071 (
            .O(N__6544),
            .I(N__6530));
    LocalMux I__1070 (
            .O(N__6541),
            .I(N__6527));
    Odrv12 I__1069 (
            .O(N__6538),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1068 (
            .O(N__6535),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1067 (
            .O(N__6530),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1066 (
            .O(N__6527),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__1065 (
            .O(N__6518),
            .I(N__6514));
    InMux I__1064 (
            .O(N__6517),
            .I(N__6511));
    LocalMux I__1063 (
            .O(N__6514),
            .I(N__6508));
    LocalMux I__1062 (
            .O(N__6511),
            .I(\U712_CHIP_RAM.N_51_0 ));
    Odrv4 I__1061 (
            .O(N__6508),
            .I(\U712_CHIP_RAM.N_51_0 ));
    CascadeMux I__1060 (
            .O(N__6503),
            .I(\U712_CHIP_RAM.N_51_0_cascade_ ));
    InMux I__1059 (
            .O(N__6500),
            .I(N__6497));
    LocalMux I__1058 (
            .O(N__6497),
            .I(\U712_CHIP_RAM.N_54_0 ));
    InMux I__1057 (
            .O(N__6494),
            .I(N__6491));
    LocalMux I__1056 (
            .O(N__6491),
            .I(\U712_CHIP_RAM.m53_ns_1 ));
    InMux I__1055 (
            .O(N__6488),
            .I(N__6478));
    InMux I__1054 (
            .O(N__6487),
            .I(N__6471));
    InMux I__1053 (
            .O(N__6486),
            .I(N__6471));
    InMux I__1052 (
            .O(N__6485),
            .I(N__6471));
    InMux I__1051 (
            .O(N__6484),
            .I(N__6464));
    InMux I__1050 (
            .O(N__6483),
            .I(N__6464));
    InMux I__1049 (
            .O(N__6482),
            .I(N__6464));
    InMux I__1048 (
            .O(N__6481),
            .I(N__6461));
    LocalMux I__1047 (
            .O(N__6478),
            .I(\U712_CHIP_RAM.N_333_mux ));
    LocalMux I__1046 (
            .O(N__6471),
            .I(\U712_CHIP_RAM.N_333_mux ));
    LocalMux I__1045 (
            .O(N__6464),
            .I(\U712_CHIP_RAM.N_333_mux ));
    LocalMux I__1044 (
            .O(N__6461),
            .I(\U712_CHIP_RAM.N_333_mux ));
    InMux I__1043 (
            .O(N__6452),
            .I(N__6449));
    LocalMux I__1042 (
            .O(N__6449),
            .I(N__6446));
    Odrv4 I__1041 (
            .O(N__6446),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0 ));
    InMux I__1040 (
            .O(N__6443),
            .I(N__6434));
    InMux I__1039 (
            .O(N__6442),
            .I(N__6431));
    InMux I__1038 (
            .O(N__6441),
            .I(N__6428));
    CascadeMux I__1037 (
            .O(N__6440),
            .I(N__6425));
    InMux I__1036 (
            .O(N__6439),
            .I(N__6418));
    InMux I__1035 (
            .O(N__6438),
            .I(N__6418));
    InMux I__1034 (
            .O(N__6437),
            .I(N__6418));
    LocalMux I__1033 (
            .O(N__6434),
            .I(N__6415));
    LocalMux I__1032 (
            .O(N__6431),
            .I(N__6410));
    LocalMux I__1031 (
            .O(N__6428),
            .I(N__6410));
    InMux I__1030 (
            .O(N__6425),
            .I(N__6407));
    LocalMux I__1029 (
            .O(N__6418),
            .I(N__6399));
    Span4Mux_h I__1028 (
            .O(N__6415),
            .I(N__6399));
    Span4Mux_v I__1027 (
            .O(N__6410),
            .I(N__6399));
    LocalMux I__1026 (
            .O(N__6407),
            .I(N__6396));
    InMux I__1025 (
            .O(N__6406),
            .I(N__6393));
    Odrv4 I__1024 (
            .O(N__6399),
            .I(DBR_SYNCZ0Z_1));
    Odrv4 I__1023 (
            .O(N__6396),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__1022 (
            .O(N__6393),
            .I(DBR_SYNCZ0Z_1));
    InMux I__1021 (
            .O(N__6386),
            .I(N__6380));
    InMux I__1020 (
            .O(N__6385),
            .I(N__6380));
    LocalMux I__1019 (
            .O(N__6380),
            .I(N__6377));
    Odrv4 I__1018 (
            .O(N__6377),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ));
    CascadeMux I__1017 (
            .O(N__6374),
            .I(N__6371));
    InMux I__1016 (
            .O(N__6371),
            .I(N__6368));
    LocalMux I__1015 (
            .O(N__6368),
            .I(N__6364));
    InMux I__1014 (
            .O(N__6367),
            .I(N__6361));
    Odrv4 I__1013 (
            .O(N__6364),
            .I(\U712_CHIP_RAM.m41_1 ));
    LocalMux I__1012 (
            .O(N__6361),
            .I(\U712_CHIP_RAM.m41_1 ));
    CascadeMux I__1011 (
            .O(N__6356),
            .I(\U712_CHIP_RAM.N_31_0_cascade_ ));
    CascadeMux I__1010 (
            .O(N__6353),
            .I(\U712_CHIP_RAM.m217_ns_1_cascade_ ));
    InMux I__1009 (
            .O(N__6350),
            .I(N__6347));
    LocalMux I__1008 (
            .O(N__6347),
            .I(\U712_CHIP_RAM.N_218 ));
    CascadeMux I__1007 (
            .O(N__6344),
            .I(\U712_CHIP_RAM.m212_ns_1_cascade_ ));
    CascadeMux I__1006 (
            .O(N__6341),
            .I(\U712_CHIP_RAM.N_30_0_cascade_ ));
    InMux I__1005 (
            .O(N__6338),
            .I(N__6335));
    LocalMux I__1004 (
            .O(N__6335),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_2 ));
    InMux I__1003 (
            .O(N__6332),
            .I(N__6329));
    LocalMux I__1002 (
            .O(N__6329),
            .I(N__6326));
    Sp12to4 I__1001 (
            .O(N__6326),
            .I(N__6323));
    Span12Mux_v I__1000 (
            .O(N__6323),
            .I(N__6320));
    Span12Mux_h I__999 (
            .O(N__6320),
            .I(N__6317));
    Odrv12 I__998 (
            .O(N__6317),
            .I(A_c_2));
    InMux I__997 (
            .O(N__6314),
            .I(N__6310));
    InMux I__996 (
            .O(N__6313),
            .I(N__6307));
    LocalMux I__995 (
            .O(N__6310),
            .I(N__6304));
    LocalMux I__994 (
            .O(N__6307),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ));
    Odrv4 I__993 (
            .O(N__6304),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ));
    InMux I__992 (
            .O(N__6299),
            .I(N__6296));
    LocalMux I__991 (
            .O(N__6296),
            .I(N__6293));
    Span4Mux_v I__990 (
            .O(N__6293),
            .I(N__6290));
    Span4Mux_v I__989 (
            .O(N__6290),
            .I(N__6287));
    Sp12to4 I__988 (
            .O(N__6287),
            .I(N__6284));
    Span12Mux_h I__987 (
            .O(N__6284),
            .I(N__6281));
    Odrv12 I__986 (
            .O(N__6281),
            .I(A_c_20));
    InMux I__985 (
            .O(N__6278),
            .I(N__6274));
    InMux I__984 (
            .O(N__6277),
            .I(N__6271));
    LocalMux I__983 (
            .O(N__6274),
            .I(N__6268));
    LocalMux I__982 (
            .O(N__6271),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ));
    Odrv4 I__981 (
            .O(N__6268),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ));
    InMux I__980 (
            .O(N__6263),
            .I(N__6259));
    InMux I__979 (
            .O(N__6262),
            .I(N__6256));
    LocalMux I__978 (
            .O(N__6259),
            .I(N__6251));
    LocalMux I__977 (
            .O(N__6256),
            .I(N__6251));
    Odrv4 I__976 (
            .O(N__6251),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__975 (
            .O(N__6248),
            .I(N__6244));
    InMux I__974 (
            .O(N__6247),
            .I(N__6241));
    LocalMux I__973 (
            .O(N__6244),
            .I(N__6238));
    LocalMux I__972 (
            .O(N__6241),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    Odrv4 I__971 (
            .O(N__6238),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    CascadeMux I__970 (
            .O(N__6233),
            .I(N__6229));
    InMux I__969 (
            .O(N__6232),
            .I(N__6226));
    InMux I__968 (
            .O(N__6229),
            .I(N__6223));
    LocalMux I__967 (
            .O(N__6226),
            .I(N__6218));
    LocalMux I__966 (
            .O(N__6223),
            .I(N__6218));
    Odrv4 I__965 (
            .O(N__6218),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__964 (
            .O(N__6215),
            .I(N__6212));
    LocalMux I__963 (
            .O(N__6212),
            .I(N__6209));
    Odrv4 I__962 (
            .O(N__6209),
            .I(\U712_CHIP_RAM.REFRESH5lt7 ));
    InMux I__961 (
            .O(N__6206),
            .I(N__6203));
    LocalMux I__960 (
            .O(N__6203),
            .I(N__6198));
    InMux I__959 (
            .O(N__6202),
            .I(N__6195));
    InMux I__958 (
            .O(N__6201),
            .I(N__6192));
    Odrv4 I__957 (
            .O(N__6198),
            .I(\U712_CHIP_RAM.N_28_0 ));
    LocalMux I__956 (
            .O(N__6195),
            .I(\U712_CHIP_RAM.N_28_0 ));
    LocalMux I__955 (
            .O(N__6192),
            .I(\U712_CHIP_RAM.N_28_0 ));
    InMux I__954 (
            .O(N__6185),
            .I(N__6182));
    LocalMux I__953 (
            .O(N__6182),
            .I(\U712_CHIP_RAM.N_219 ));
    InMux I__952 (
            .O(N__6179),
            .I(N__6176));
    LocalMux I__951 (
            .O(N__6176),
            .I(\U712_CHIP_RAM.d_N_6_5 ));
    InMux I__950 (
            .O(N__6173),
            .I(N__6170));
    LocalMux I__949 (
            .O(N__6170),
            .I(\U712_CHIP_RAM.d_N_6_1 ));
    InMux I__948 (
            .O(N__6167),
            .I(N__6164));
    LocalMux I__947 (
            .O(N__6164),
            .I(N__6161));
    Odrv4 I__946 (
            .O(N__6161),
            .I(\U712_CHIP_RAM.N_353_mux ));
    CascadeMux I__945 (
            .O(N__6158),
            .I(\U712_CHIP_RAM.N_168_0_cascade_ ));
    InMux I__944 (
            .O(N__6155),
            .I(N__6152));
    LocalMux I__943 (
            .O(N__6152),
            .I(\U712_CHIP_RAM.m64_ns_1 ));
    CascadeMux I__942 (
            .O(N__6149),
            .I(\U712_CHIP_RAM.i67_mux_cascade_ ));
    InMux I__941 (
            .O(N__6146),
            .I(N__6143));
    LocalMux I__940 (
            .O(N__6143),
            .I(N__6140));
    Odrv4 I__939 (
            .O(N__6140),
            .I(\U712_CHIP_RAM.m66_ns_1 ));
    InMux I__938 (
            .O(N__6137),
            .I(N__6134));
    LocalMux I__937 (
            .O(N__6134),
            .I(\U712_CHIP_RAM.N_146_0 ));
    CascadeMux I__936 (
            .O(N__6131),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_2_cascade_ ));
    CascadeMux I__935 (
            .O(N__6128),
            .I(\U712_CHIP_RAM.N_151_0_cascade_ ));
    CascadeMux I__934 (
            .O(N__6125),
            .I(N__6122));
    InMux I__933 (
            .O(N__6122),
            .I(N__6117));
    InMux I__932 (
            .O(N__6121),
            .I(N__6112));
    InMux I__931 (
            .O(N__6120),
            .I(N__6112));
    LocalMux I__930 (
            .O(N__6117),
            .I(N__6107));
    LocalMux I__929 (
            .O(N__6112),
            .I(N__6107));
    Odrv4 I__928 (
            .O(N__6107),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ));
    InMux I__927 (
            .O(N__6104),
            .I(N__6101));
    LocalMux I__926 (
            .O(N__6101),
            .I(U712_REG_SM_UDSn_6_0));
    IoInMux I__925 (
            .O(N__6098),
            .I(N__6095));
    LocalMux I__924 (
            .O(N__6095),
            .I(N__6092));
    Span4Mux_s3_v I__923 (
            .O(N__6092),
            .I(N__6089));
    Span4Mux_v I__922 (
            .O(N__6089),
            .I(N__6086));
    Span4Mux_v I__921 (
            .O(N__6086),
            .I(N__6083));
    Sp12to4 I__920 (
            .O(N__6083),
            .I(N__6079));
    InMux I__919 (
            .O(N__6082),
            .I(N__6076));
    Odrv12 I__918 (
            .O(N__6079),
            .I(UDSn_c));
    LocalMux I__917 (
            .O(N__6076),
            .I(UDSn_c));
    InMux I__916 (
            .O(N__6071),
            .I(N__6068));
    LocalMux I__915 (
            .O(N__6068),
            .I(N__6065));
    Span4Mux_v I__914 (
            .O(N__6065),
            .I(N__6061));
    InMux I__913 (
            .O(N__6064),
            .I(N__6058));
    Span4Mux_v I__912 (
            .O(N__6061),
            .I(N__6055));
    LocalMux I__911 (
            .O(N__6058),
            .I(N__6052));
    Sp12to4 I__910 (
            .O(N__6055),
            .I(N__6049));
    Span4Mux_h I__909 (
            .O(N__6052),
            .I(N__6046));
    Odrv12 I__908 (
            .O(N__6049),
            .I(DBRn_c_i));
    Odrv4 I__907 (
            .O(N__6046),
            .I(DBRn_c_i));
    IoInMux I__906 (
            .O(N__6041),
            .I(N__6038));
    LocalMux I__905 (
            .O(N__6038),
            .I(N__6035));
    IoSpan4Mux I__904 (
            .O(N__6035),
            .I(N__6032));
    Span4Mux_s3_h I__903 (
            .O(N__6032),
            .I(N__6029));
    Sp12to4 I__902 (
            .O(N__6029),
            .I(N__6026));
    Span12Mux_h I__901 (
            .O(N__6026),
            .I(N__6023));
    Odrv12 I__900 (
            .O(N__6023),
            .I(CMA_c_8));
    IoInMux I__899 (
            .O(N__6020),
            .I(N__6016));
    InMux I__898 (
            .O(N__6019),
            .I(N__6013));
    LocalMux I__897 (
            .O(N__6016),
            .I(N__6010));
    LocalMux I__896 (
            .O(N__6013),
            .I(N__6007));
    Span12Mux_s4_v I__895 (
            .O(N__6010),
            .I(N__6004));
    Span4Mux_v I__894 (
            .O(N__6007),
            .I(N__6001));
    Span12Mux_v I__893 (
            .O(N__6004),
            .I(N__5998));
    Span4Mux_h I__892 (
            .O(N__6001),
            .I(N__5995));
    Span12Mux_h I__891 (
            .O(N__5998),
            .I(N__5992));
    Sp12to4 I__890 (
            .O(N__5995),
            .I(N__5989));
    Odrv12 I__889 (
            .O(N__5992),
            .I(A_c_9));
    Odrv12 I__888 (
            .O(N__5989),
            .I(A_c_9));
    CascadeMux I__887 (
            .O(N__5984),
            .I(\U712_CHIP_RAM.m186_0_cascade_ ));
    InMux I__886 (
            .O(N__5981),
            .I(N__5978));
    LocalMux I__885 (
            .O(N__5978),
            .I(N__5975));
    Sp12to4 I__884 (
            .O(N__5975),
            .I(N__5972));
    Span12Mux_v I__883 (
            .O(N__5972),
            .I(N__5969));
    Span12Mux_h I__882 (
            .O(N__5969),
            .I(N__5966));
    Odrv12 I__881 (
            .O(N__5966),
            .I(A_c_17));
    CascadeMux I__880 (
            .O(N__5963),
            .I(\U712_CHIP_RAM.m192_0_cascade_ ));
    InMux I__879 (
            .O(N__5960),
            .I(N__5956));
    InMux I__878 (
            .O(N__5959),
            .I(N__5953));
    LocalMux I__877 (
            .O(N__5956),
            .I(N__5950));
    LocalMux I__876 (
            .O(N__5953),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    Odrv4 I__875 (
            .O(N__5950),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    InMux I__874 (
            .O(N__5945),
            .I(N__5942));
    LocalMux I__873 (
            .O(N__5942),
            .I(\U712_CHIP_RAM.m192_1 ));
    CascadeMux I__872 (
            .O(N__5939),
            .I(N__5936));
    InMux I__871 (
            .O(N__5936),
            .I(N__5933));
    LocalMux I__870 (
            .O(N__5933),
            .I(N__5930));
    Odrv4 I__869 (
            .O(N__5930),
            .I(\U712_CHIP_RAM.N_215 ));
    InMux I__868 (
            .O(N__5927),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__867 (
            .O(N__5924),
            .I(N__5921));
    LocalMux I__866 (
            .O(N__5921),
            .I(N__5918));
    Odrv4 I__865 (
            .O(N__5918),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    InMux I__864 (
            .O(N__5915),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    InMux I__863 (
            .O(N__5912),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    InMux I__862 (
            .O(N__5909),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__861 (
            .O(N__5906),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__860 (
            .O(N__5903),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    CascadeMux I__859 (
            .O(N__5900),
            .I(N__5897));
    InMux I__858 (
            .O(N__5897),
            .I(N__5894));
    LocalMux I__857 (
            .O(N__5894),
            .I(N__5884));
    InMux I__856 (
            .O(N__5893),
            .I(N__5881));
    InMux I__855 (
            .O(N__5892),
            .I(N__5872));
    InMux I__854 (
            .O(N__5891),
            .I(N__5872));
    InMux I__853 (
            .O(N__5890),
            .I(N__5872));
    InMux I__852 (
            .O(N__5889),
            .I(N__5872));
    InMux I__851 (
            .O(N__5888),
            .I(N__5867));
    InMux I__850 (
            .O(N__5887),
            .I(N__5867));
    Odrv4 I__849 (
            .O(N__5884),
            .I(\U712_CHIP_RAM.N_56_0_i ));
    LocalMux I__848 (
            .O(N__5881),
            .I(\U712_CHIP_RAM.N_56_0_i ));
    LocalMux I__847 (
            .O(N__5872),
            .I(\U712_CHIP_RAM.N_56_0_i ));
    LocalMux I__846 (
            .O(N__5867),
            .I(\U712_CHIP_RAM.N_56_0_i ));
    InMux I__845 (
            .O(N__5858),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    CEMux I__844 (
            .O(N__5855),
            .I(N__5851));
    CEMux I__843 (
            .O(N__5854),
            .I(N__5847));
    LocalMux I__842 (
            .O(N__5851),
            .I(N__5844));
    CEMux I__841 (
            .O(N__5850),
            .I(N__5841));
    LocalMux I__840 (
            .O(N__5847),
            .I(N__5838));
    Span4Mux_v I__839 (
            .O(N__5844),
            .I(N__5835));
    LocalMux I__838 (
            .O(N__5841),
            .I(N__5832));
    Odrv4 I__837 (
            .O(N__5838),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    Odrv4 I__836 (
            .O(N__5835),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    Odrv4 I__835 (
            .O(N__5832),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    InMux I__834 (
            .O(N__5825),
            .I(N__5822));
    LocalMux I__833 (
            .O(N__5822),
            .I(\U712_CHIP_RAM.N_330 ));
    InMux I__832 (
            .O(N__5819),
            .I(N__5816));
    LocalMux I__831 (
            .O(N__5816),
            .I(N__5813));
    Odrv4 I__830 (
            .O(N__5813),
            .I(\U712_CHIP_RAM.m38_1 ));
    CascadeMux I__829 (
            .O(N__5810),
            .I(\U712_CHIP_RAM.N_34_0_cascade_ ));
    CascadeMux I__828 (
            .O(N__5807),
            .I(N__5804));
    InMux I__827 (
            .O(N__5804),
            .I(N__5801));
    LocalMux I__826 (
            .O(N__5801),
            .I(\U712_CHIP_RAM.N_359 ));
    InMux I__825 (
            .O(N__5798),
            .I(N__5792));
    InMux I__824 (
            .O(N__5797),
            .I(N__5785));
    InMux I__823 (
            .O(N__5796),
            .I(N__5785));
    InMux I__822 (
            .O(N__5795),
            .I(N__5785));
    LocalMux I__821 (
            .O(N__5792),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__820 (
            .O(N__5785),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    InMux I__819 (
            .O(N__5780),
            .I(N__5776));
    InMux I__818 (
            .O(N__5779),
            .I(N__5773));
    LocalMux I__817 (
            .O(N__5776),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ));
    LocalMux I__816 (
            .O(N__5773),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ));
    CascadeMux I__815 (
            .O(N__5768),
            .I(\U712_CHIP_RAM.N_28_0_cascade_ ));
    CascadeMux I__814 (
            .O(N__5765),
            .I(\U712_CHIP_RAM.N_47_0_cascade_ ));
    CascadeMux I__813 (
            .O(N__5762),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_cascade_ ));
    CEMux I__812 (
            .O(N__5759),
            .I(N__5756));
    LocalMux I__811 (
            .O(N__5756),
            .I(N__5753));
    Span4Mux_v I__810 (
            .O(N__5753),
            .I(N__5750));
    Odrv4 I__809 (
            .O(N__5750),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0 ));
    CascadeMux I__808 (
            .O(N__5747),
            .I(\U712_CHIP_RAM.N_146_0_cascade_ ));
    CascadeMux I__807 (
            .O(N__5744),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_3_cascade_ ));
    InMux I__806 (
            .O(N__5741),
            .I(N__5738));
    LocalMux I__805 (
            .O(N__5738),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_3 ));
    CascadeMux I__804 (
            .O(N__5735),
            .I(\U712_CHIP_RAM.N_154_0_cascade_ ));
    InMux I__803 (
            .O(N__5732),
            .I(N__5729));
    LocalMux I__802 (
            .O(N__5729),
            .I(N__5726));
    Odrv4 I__801 (
            .O(N__5726),
            .I(\U712_CHIP_RAM.N_7_0 ));
    InMux I__800 (
            .O(N__5723),
            .I(N__5719));
    InMux I__799 (
            .O(N__5722),
            .I(N__5716));
    LocalMux I__798 (
            .O(N__5719),
            .I(N_86_0));
    LocalMux I__797 (
            .O(N__5716),
            .I(N_86_0));
    CascadeMux I__796 (
            .O(N__5711),
            .I(N__5706));
    CascadeMux I__795 (
            .O(N__5710),
            .I(N__5702));
    InMux I__794 (
            .O(N__5709),
            .I(N__5696));
    InMux I__793 (
            .O(N__5706),
            .I(N__5693));
    InMux I__792 (
            .O(N__5705),
            .I(N__5690));
    InMux I__791 (
            .O(N__5702),
            .I(N__5687));
    CascadeMux I__790 (
            .O(N__5701),
            .I(N__5684));
    InMux I__789 (
            .O(N__5700),
            .I(N__5678));
    InMux I__788 (
            .O(N__5699),
            .I(N__5675));
    LocalMux I__787 (
            .O(N__5696),
            .I(N__5668));
    LocalMux I__786 (
            .O(N__5693),
            .I(N__5668));
    LocalMux I__785 (
            .O(N__5690),
            .I(N__5668));
    LocalMux I__784 (
            .O(N__5687),
            .I(N__5662));
    InMux I__783 (
            .O(N__5684),
            .I(N__5659));
    InMux I__782 (
            .O(N__5683),
            .I(N__5656));
    InMux I__781 (
            .O(N__5682),
            .I(N__5651));
    InMux I__780 (
            .O(N__5681),
            .I(N__5651));
    LocalMux I__779 (
            .O(N__5678),
            .I(N__5646));
    LocalMux I__778 (
            .O(N__5675),
            .I(N__5646));
    Span4Mux_v I__777 (
            .O(N__5668),
            .I(N__5643));
    InMux I__776 (
            .O(N__5667),
            .I(N__5636));
    InMux I__775 (
            .O(N__5666),
            .I(N__5636));
    InMux I__774 (
            .O(N__5665),
            .I(N__5636));
    Span4Mux_h I__773 (
            .O(N__5662),
            .I(N__5633));
    LocalMux I__772 (
            .O(N__5659),
            .I(U712_REG_SM_C3_SYNC_1));
    LocalMux I__771 (
            .O(N__5656),
            .I(U712_REG_SM_C3_SYNC_1));
    LocalMux I__770 (
            .O(N__5651),
            .I(U712_REG_SM_C3_SYNC_1));
    Odrv4 I__769 (
            .O(N__5646),
            .I(U712_REG_SM_C3_SYNC_1));
    Odrv4 I__768 (
            .O(N__5643),
            .I(U712_REG_SM_C3_SYNC_1));
    LocalMux I__767 (
            .O(N__5636),
            .I(U712_REG_SM_C3_SYNC_1));
    Odrv4 I__766 (
            .O(N__5633),
            .I(U712_REG_SM_C3_SYNC_1));
    IoInMux I__765 (
            .O(N__5618),
            .I(N__5615));
    LocalMux I__764 (
            .O(N__5615),
            .I(N__5611));
    IoInMux I__763 (
            .O(N__5614),
            .I(N__5608));
    IoSpan4Mux I__762 (
            .O(N__5611),
            .I(N__5605));
    LocalMux I__761 (
            .O(N__5608),
            .I(N__5602));
    Sp12to4 I__760 (
            .O(N__5605),
            .I(N__5599));
    Span4Mux_s1_v I__759 (
            .O(N__5602),
            .I(N__5596));
    Span12Mux_s7_h I__758 (
            .O(N__5599),
            .I(N__5593));
    Sp12to4 I__757 (
            .O(N__5596),
            .I(N__5590));
    Span12Mux_h I__756 (
            .O(N__5593),
            .I(N__5585));
    Span12Mux_h I__755 (
            .O(N__5590),
            .I(N__5585));
    Odrv12 I__754 (
            .O(N__5585),
            .I(BLSn_c));
    CEMux I__753 (
            .O(N__5582),
            .I(N__5579));
    LocalMux I__752 (
            .O(N__5579),
            .I(N__5576));
    Span4Mux_v I__751 (
            .O(N__5576),
            .I(N__5573));
    Span4Mux_h I__750 (
            .O(N__5573),
            .I(N__5570));
    Odrv4 I__749 (
            .O(N__5570),
            .I(\U712_REG_SM.N_86_0_0 ));
    CascadeMux I__748 (
            .O(N__5567),
            .I(\U712_CYCLE_TERM.N_36_0_cascade_ ));
    IoInMux I__747 (
            .O(N__5564),
            .I(N__5559));
    IoInMux I__746 (
            .O(N__5563),
            .I(N__5556));
    IoInMux I__745 (
            .O(N__5562),
            .I(N__5553));
    LocalMux I__744 (
            .O(N__5559),
            .I(N__5550));
    LocalMux I__743 (
            .O(N__5556),
            .I(N__5547));
    LocalMux I__742 (
            .O(N__5553),
            .I(N__5544));
    Span4Mux_s1_h I__741 (
            .O(N__5550),
            .I(N__5541));
    Span4Mux_s0_v I__740 (
            .O(N__5547),
            .I(N__5538));
    Span4Mux_s3_v I__739 (
            .O(N__5544),
            .I(N__5535));
    Sp12to4 I__738 (
            .O(N__5541),
            .I(N__5532));
    Span4Mux_h I__737 (
            .O(N__5538),
            .I(N__5529));
    Span4Mux_v I__736 (
            .O(N__5535),
            .I(N__5526));
    Span12Mux_s11_v I__735 (
            .O(N__5532),
            .I(N__5523));
    Sp12to4 I__734 (
            .O(N__5529),
            .I(N__5520));
    Span4Mux_h I__733 (
            .O(N__5526),
            .I(N__5517));
    Span12Mux_h I__732 (
            .O(N__5523),
            .I(N__5513));
    Span12Mux_h I__731 (
            .O(N__5520),
            .I(N__5510));
    Span4Mux_h I__730 (
            .O(N__5517),
            .I(N__5507));
    InMux I__729 (
            .O(N__5516),
            .I(N__5504));
    Odrv12 I__728 (
            .O(N__5513),
            .I(TACK_OUT));
    Odrv12 I__727 (
            .O(N__5510),
            .I(TACK_OUT));
    Odrv4 I__726 (
            .O(N__5507),
            .I(TACK_OUT));
    LocalMux I__725 (
            .O(N__5504),
            .I(TACK_OUT));
    InMux I__724 (
            .O(N__5495),
            .I(N__5490));
    InMux I__723 (
            .O(N__5494),
            .I(N__5485));
    InMux I__722 (
            .O(N__5493),
            .I(N__5485));
    LocalMux I__721 (
            .O(N__5490),
            .I(N__5480));
    LocalMux I__720 (
            .O(N__5485),
            .I(N__5480));
    Span4Mux_h I__719 (
            .O(N__5480),
            .I(N__5476));
    InMux I__718 (
            .O(N__5479),
            .I(N__5473));
    Span4Mux_v I__717 (
            .O(N__5476),
            .I(N__5470));
    LocalMux I__716 (
            .O(N__5473),
            .I(\U712_CYCLE_TERM.TACK_STARTZ0 ));
    Odrv4 I__715 (
            .O(N__5470),
            .I(\U712_CYCLE_TERM.TACK_STARTZ0 ));
    InMux I__714 (
            .O(N__5465),
            .I(N__5458));
    InMux I__713 (
            .O(N__5464),
            .I(N__5449));
    InMux I__712 (
            .O(N__5463),
            .I(N__5449));
    InMux I__711 (
            .O(N__5462),
            .I(N__5449));
    InMux I__710 (
            .O(N__5461),
            .I(N__5449));
    LocalMux I__709 (
            .O(N__5458),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__708 (
            .O(N__5449),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    CascadeMux I__707 (
            .O(N__5444),
            .I(N__5441));
    InMux I__706 (
            .O(N__5441),
            .I(N__5436));
    InMux I__705 (
            .O(N__5440),
            .I(N__5431));
    InMux I__704 (
            .O(N__5439),
            .I(N__5431));
    LocalMux I__703 (
            .O(N__5436),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__702 (
            .O(N__5431),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    InMux I__701 (
            .O(N__5426),
            .I(N__5423));
    LocalMux I__700 (
            .O(N__5423),
            .I(\U712_CHIP_RAM.N_83_0 ));
    CascadeMux I__699 (
            .O(N__5420),
            .I(\U712_CHIP_RAM.N_94_0_cascade_ ));
    InMux I__698 (
            .O(N__5417),
            .I(N__5412));
    InMux I__697 (
            .O(N__5416),
            .I(N__5405));
    InMux I__696 (
            .O(N__5415),
            .I(N__5405));
    LocalMux I__695 (
            .O(N__5412),
            .I(N__5402));
    InMux I__694 (
            .O(N__5411),
            .I(N__5399));
    InMux I__693 (
            .O(N__5410),
            .I(N__5396));
    LocalMux I__692 (
            .O(N__5405),
            .I(U712_REG_SM_STATE_COUNT_1));
    Odrv4 I__691 (
            .O(N__5402),
            .I(U712_REG_SM_STATE_COUNT_1));
    LocalMux I__690 (
            .O(N__5399),
            .I(U712_REG_SM_STATE_COUNT_1));
    LocalMux I__689 (
            .O(N__5396),
            .I(U712_REG_SM_STATE_COUNT_1));
    InMux I__688 (
            .O(N__5387),
            .I(N__5383));
    InMux I__687 (
            .O(N__5386),
            .I(N__5380));
    LocalMux I__686 (
            .O(N__5383),
            .I(U712_REG_SM_STATE_COUNT_2));
    LocalMux I__685 (
            .O(N__5380),
            .I(U712_REG_SM_STATE_COUNT_2));
    InMux I__684 (
            .O(N__5375),
            .I(N__5371));
    CascadeMux I__683 (
            .O(N__5374),
            .I(N__5368));
    LocalMux I__682 (
            .O(N__5371),
            .I(N__5365));
    InMux I__681 (
            .O(N__5368),
            .I(N__5362));
    Odrv4 I__680 (
            .O(N__5365),
            .I(DBR_SYNC_i_1));
    LocalMux I__679 (
            .O(N__5362),
            .I(DBR_SYNC_i_1));
    InMux I__678 (
            .O(N__5357),
            .I(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ));
    InMux I__677 (
            .O(N__5354),
            .I(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ));
    InMux I__676 (
            .O(N__5351),
            .I(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_2 ));
    InMux I__675 (
            .O(N__5348),
            .I(N__5345));
    LocalMux I__674 (
            .O(N__5345),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1 ));
    CascadeMux I__673 (
            .O(N__5342),
            .I(N__5339));
    InMux I__672 (
            .O(N__5339),
            .I(N__5336));
    LocalMux I__671 (
            .O(N__5336),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2 ));
    InMux I__670 (
            .O(N__5333),
            .I(N__5327));
    InMux I__669 (
            .O(N__5332),
            .I(N__5327));
    LocalMux I__668 (
            .O(N__5327),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ));
    CascadeMux I__667 (
            .O(N__5324),
            .I(N__5321));
    InMux I__666 (
            .O(N__5321),
            .I(N__5315));
    InMux I__665 (
            .O(N__5320),
            .I(N__5315));
    LocalMux I__664 (
            .O(N__5315),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_1 ));
    CascadeMux I__663 (
            .O(N__5312),
            .I(N__5309));
    InMux I__662 (
            .O(N__5309),
            .I(N__5306));
    LocalMux I__661 (
            .O(N__5306),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3 ));
    InMux I__660 (
            .O(N__5303),
            .I(N__5297));
    InMux I__659 (
            .O(N__5302),
            .I(N__5297));
    LocalMux I__658 (
            .O(N__5297),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ));
    InMux I__657 (
            .O(N__5294),
            .I(N__5290));
    IoInMux I__656 (
            .O(N__5293),
            .I(N__5287));
    LocalMux I__655 (
            .O(N__5290),
            .I(N__5284));
    LocalMux I__654 (
            .O(N__5287),
            .I(N__5281));
    Span4Mux_v I__653 (
            .O(N__5284),
            .I(N__5278));
    IoSpan4Mux I__652 (
            .O(N__5281),
            .I(N__5275));
    Sp12to4 I__651 (
            .O(N__5278),
            .I(N__5272));
    IoSpan4Mux I__650 (
            .O(N__5275),
            .I(N__5269));
    Span12Mux_h I__649 (
            .O(N__5272),
            .I(N__5266));
    IoSpan4Mux I__648 (
            .O(N__5269),
            .I(N__5263));
    Odrv12 I__647 (
            .O(N__5266),
            .I(C1_c));
    Odrv4 I__646 (
            .O(N__5263),
            .I(C1_c));
    InMux I__645 (
            .O(N__5258),
            .I(N__5255));
    LocalMux I__644 (
            .O(N__5255),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    InMux I__643 (
            .O(N__5252),
            .I(N__5249));
    LocalMux I__642 (
            .O(N__5249),
            .I(\U712_CHIP_RAM.m231_0 ));
    InMux I__641 (
            .O(N__5246),
            .I(N__5243));
    LocalMux I__640 (
            .O(N__5243),
            .I(\U712_CHIP_RAM.N_236 ));
    InMux I__639 (
            .O(N__5240),
            .I(N__5235));
    InMux I__638 (
            .O(N__5239),
            .I(N__5232));
    InMux I__637 (
            .O(N__5238),
            .I(N__5229));
    LocalMux I__636 (
            .O(N__5235),
            .I(N__5224));
    LocalMux I__635 (
            .O(N__5232),
            .I(N__5224));
    LocalMux I__634 (
            .O(N__5229),
            .I(U712_REG_SM_STATE_COUNT_0_sqmuxa_1));
    Odrv4 I__633 (
            .O(N__5224),
            .I(U712_REG_SM_STATE_COUNT_0_sqmuxa_1));
    CascadeMux I__632 (
            .O(N__5219),
            .I(\U712_CHIP_RAM.N_83_0_cascade_ ));
    CascadeMux I__631 (
            .O(N__5216),
            .I(N__5212));
    CascadeMux I__630 (
            .O(N__5215),
            .I(N__5209));
    InMux I__629 (
            .O(N__5212),
            .I(N__5204));
    InMux I__628 (
            .O(N__5209),
            .I(N__5201));
    InMux I__627 (
            .O(N__5208),
            .I(N__5196));
    InMux I__626 (
            .O(N__5207),
            .I(N__5196));
    LocalMux I__625 (
            .O(N__5204),
            .I(U712_REG_SM_REG_CYCLE_START));
    LocalMux I__624 (
            .O(N__5201),
            .I(U712_REG_SM_REG_CYCLE_START));
    LocalMux I__623 (
            .O(N__5196),
            .I(U712_REG_SM_REG_CYCLE_START));
    InMux I__622 (
            .O(N__5189),
            .I(N__5183));
    InMux I__621 (
            .O(N__5188),
            .I(N__5183));
    LocalMux I__620 (
            .O(N__5183),
            .I(U712_REG_SM_START_RST));
    InMux I__619 (
            .O(N__5180),
            .I(N__5177));
    LocalMux I__618 (
            .O(N__5177),
            .I(N__5174));
    Odrv4 I__617 (
            .O(N__5174),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_3 ));
    InMux I__616 (
            .O(N__5171),
            .I(N__5168));
    LocalMux I__615 (
            .O(N__5168),
            .I(N__5165));
    Span4Mux_h I__614 (
            .O(N__5165),
            .I(N__5162));
    Span4Mux_v I__613 (
            .O(N__5162),
            .I(N__5158));
    IoInMux I__612 (
            .O(N__5161),
            .I(N__5155));
    Span4Mux_v I__611 (
            .O(N__5158),
            .I(N__5152));
    LocalMux I__610 (
            .O(N__5155),
            .I(N__5149));
    Span4Mux_v I__609 (
            .O(N__5152),
            .I(N__5146));
    IoSpan4Mux I__608 (
            .O(N__5149),
            .I(N__5143));
    Odrv4 I__607 (
            .O(N__5146),
            .I(RAMENn_c));
    Odrv4 I__606 (
            .O(N__5143),
            .I(RAMENn_c));
    CascadeMux I__605 (
            .O(N__5138),
            .I(N__5134));
    InMux I__604 (
            .O(N__5137),
            .I(N__5129));
    InMux I__603 (
            .O(N__5134),
            .I(N__5129));
    LocalMux I__602 (
            .O(N__5129),
            .I(N__5126));
    Span4Mux_v I__601 (
            .O(N__5126),
            .I(N__5123));
    Sp12to4 I__600 (
            .O(N__5123),
            .I(N__5120));
    Span12Mux_h I__599 (
            .O(N__5120),
            .I(N__5117));
    Span12Mux_v I__598 (
            .O(N__5117),
            .I(N__5114));
    Odrv12 I__597 (
            .O(N__5114),
            .I(TSn_c));
    CascadeMux I__596 (
            .O(N__5111),
            .I(\U712_CHIP_RAM.m223_ns_1_cascade_ ));
    InMux I__595 (
            .O(N__5108),
            .I(N__5105));
    LocalMux I__594 (
            .O(N__5105),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_5 ));
    InMux I__593 (
            .O(N__5102),
            .I(N__5098));
    InMux I__592 (
            .O(N__5101),
            .I(N__5095));
    LocalMux I__591 (
            .O(N__5098),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_4 ));
    LocalMux I__590 (
            .O(N__5095),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_4 ));
    InMux I__589 (
            .O(N__5090),
            .I(N__5087));
    LocalMux I__588 (
            .O(N__5087),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__587 (
            .O(N__5084),
            .I(bfn_9_11_0_));
    InMux I__586 (
            .O(N__5081),
            .I(N__5077));
    InMux I__585 (
            .O(N__5080),
            .I(N__5074));
    LocalMux I__584 (
            .O(N__5077),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    LocalMux I__583 (
            .O(N__5074),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    InMux I__582 (
            .O(N__5069),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__581 (
            .O(N__5066),
            .I(N__5062));
    InMux I__580 (
            .O(N__5065),
            .I(N__5059));
    LocalMux I__579 (
            .O(N__5062),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    LocalMux I__578 (
            .O(N__5059),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    InMux I__577 (
            .O(N__5054),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__576 (
            .O(N__5051),
            .I(N__5047));
    InMux I__575 (
            .O(N__5050),
            .I(N__5044));
    LocalMux I__574 (
            .O(N__5047),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__573 (
            .O(N__5044),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__572 (
            .O(N__5039),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    CascadeMux I__571 (
            .O(N__5036),
            .I(N__5032));
    InMux I__570 (
            .O(N__5035),
            .I(N__5029));
    InMux I__569 (
            .O(N__5032),
            .I(N__5026));
    LocalMux I__568 (
            .O(N__5029),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__567 (
            .O(N__5026),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__566 (
            .O(N__5021),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__565 (
            .O(N__5018),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__564 (
            .O(N__5015),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__563 (
            .O(N__5012),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    ClkMux I__562 (
            .O(N__5009),
            .I(N__4982));
    ClkMux I__561 (
            .O(N__5008),
            .I(N__4982));
    ClkMux I__560 (
            .O(N__5007),
            .I(N__4982));
    ClkMux I__559 (
            .O(N__5006),
            .I(N__4982));
    ClkMux I__558 (
            .O(N__5005),
            .I(N__4982));
    ClkMux I__557 (
            .O(N__5004),
            .I(N__4982));
    ClkMux I__556 (
            .O(N__5003),
            .I(N__4982));
    ClkMux I__555 (
            .O(N__5002),
            .I(N__4982));
    ClkMux I__554 (
            .O(N__5001),
            .I(N__4982));
    GlobalMux I__553 (
            .O(N__4982),
            .I(N__4979));
    gio2CtrlBuf I__552 (
            .O(N__4979),
            .I(C1_c_g));
    InMux I__551 (
            .O(N__4976),
            .I(N__4973));
    LocalMux I__550 (
            .O(N__4973),
            .I(N__4970));
    Span4Mux_v I__549 (
            .O(N__4970),
            .I(N__4967));
    Span4Mux_v I__548 (
            .O(N__4967),
            .I(N__4964));
    Sp12to4 I__547 (
            .O(N__4964),
            .I(N__4961));
    Span12Mux_h I__546 (
            .O(N__4961),
            .I(N__4958));
    Odrv12 I__545 (
            .O(N__4958),
            .I(REGSPACEn_c));
    InMux I__544 (
            .O(N__4955),
            .I(N__4950));
    InMux I__543 (
            .O(N__4954),
            .I(N__4944));
    InMux I__542 (
            .O(N__4953),
            .I(N__4944));
    LocalMux I__541 (
            .O(N__4950),
            .I(N__4941));
    InMux I__540 (
            .O(N__4949),
            .I(N__4938));
    LocalMux I__539 (
            .O(N__4944),
            .I(U712_REG_SM_WRITE_CYCLE));
    Odrv4 I__538 (
            .O(N__4941),
            .I(U712_REG_SM_WRITE_CYCLE));
    LocalMux I__537 (
            .O(N__4938),
            .I(U712_REG_SM_WRITE_CYCLE));
    IoInMux I__536 (
            .O(N__4931),
            .I(N__4928));
    LocalMux I__535 (
            .O(N__4928),
            .I(N__4925));
    IoSpan4Mux I__534 (
            .O(N__4925),
            .I(N__4922));
    Span4Mux_s3_v I__533 (
            .O(N__4922),
            .I(N__4919));
    Sp12to4 I__532 (
            .O(N__4919),
            .I(N__4916));
    Span12Mux_s11_v I__531 (
            .O(N__4916),
            .I(N__4912));
    InMux I__530 (
            .O(N__4915),
            .I(N__4909));
    Odrv12 I__529 (
            .O(N__4912),
            .I(PRnW_c));
    LocalMux I__528 (
            .O(N__4909),
            .I(PRnW_c));
    InMux I__527 (
            .O(N__4904),
            .I(N__4901));
    LocalMux I__526 (
            .O(N__4901),
            .I(N__4898));
    Odrv4 I__525 (
            .O(N__4898),
            .I(\U712_CHIP_RAM.N_332 ));
    InMux I__524 (
            .O(N__4895),
            .I(N__4892));
    LocalMux I__523 (
            .O(N__4892),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ));
    InMux I__522 (
            .O(N__4889),
            .I(N__4886));
    LocalMux I__521 (
            .O(N__4886),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_2 ));
    IoInMux I__520 (
            .O(N__4883),
            .I(N__4879));
    IoInMux I__519 (
            .O(N__4882),
            .I(N__4875));
    LocalMux I__518 (
            .O(N__4879),
            .I(N__4872));
    IoInMux I__517 (
            .O(N__4878),
            .I(N__4869));
    LocalMux I__516 (
            .O(N__4875),
            .I(N__4866));
    IoSpan4Mux I__515 (
            .O(N__4872),
            .I(N__4863));
    LocalMux I__514 (
            .O(N__4869),
            .I(N__4860));
    Span4Mux_s0_h I__513 (
            .O(N__4866),
            .I(N__4857));
    Span4Mux_s0_v I__512 (
            .O(N__4863),
            .I(N__4854));
    IoSpan4Mux I__511 (
            .O(N__4860),
            .I(N__4851));
    Sp12to4 I__510 (
            .O(N__4857),
            .I(N__4848));
    Span4Mux_v I__509 (
            .O(N__4854),
            .I(N__4845));
    IoSpan4Mux I__508 (
            .O(N__4851),
            .I(N__4842));
    Span12Mux_v I__507 (
            .O(N__4848),
            .I(N__4837));
    Sp12to4 I__506 (
            .O(N__4845),
            .I(N__4834));
    Span4Mux_s2_v I__505 (
            .O(N__4842),
            .I(N__4831));
    InMux I__504 (
            .O(N__4841),
            .I(N__4828));
    InMux I__503 (
            .O(N__4840),
            .I(N__4825));
    Span12Mux_h I__502 (
            .O(N__4837),
            .I(N__4816));
    Span12Mux_h I__501 (
            .O(N__4834),
            .I(N__4816));
    Sp12to4 I__500 (
            .O(N__4831),
            .I(N__4816));
    LocalMux I__499 (
            .O(N__4828),
            .I(N__4816));
    LocalMux I__498 (
            .O(N__4825),
            .I(TACK_EN));
    Odrv12 I__497 (
            .O(N__4816),
            .I(TACK_EN));
    SRMux I__496 (
            .O(N__4811),
            .I(N__4808));
    LocalMux I__495 (
            .O(N__4808),
            .I(\U712_CYCLE_TERM.TACK_RST_0_i ));
    InMux I__494 (
            .O(N__4805),
            .I(N__4802));
    LocalMux I__493 (
            .O(N__4802),
            .I(U712_REG_SM_STATE_COUNT_7));
    InMux I__492 (
            .O(N__4799),
            .I(N__4791));
    InMux I__491 (
            .O(N__4798),
            .I(N__4791));
    InMux I__490 (
            .O(N__4797),
            .I(N__4786));
    InMux I__489 (
            .O(N__4796),
            .I(N__4786));
    LocalMux I__488 (
            .O(N__4791),
            .I(U712_REG_SM_STATE_COUNT_0));
    LocalMux I__487 (
            .O(N__4786),
            .I(U712_REG_SM_STATE_COUNT_0));
    InMux I__486 (
            .O(N__4781),
            .I(N__4778));
    LocalMux I__485 (
            .O(N__4778),
            .I(\U712_CHIP_RAM.N_79_0 ));
    InMux I__484 (
            .O(N__4775),
            .I(N__4771));
    InMux I__483 (
            .O(N__4774),
            .I(N__4768));
    LocalMux I__482 (
            .O(N__4771),
            .I(U712_REG_SM_STATE_COUNT_5));
    LocalMux I__481 (
            .O(N__4768),
            .I(U712_REG_SM_STATE_COUNT_5));
    InMux I__480 (
            .O(N__4763),
            .I(N__4760));
    LocalMux I__479 (
            .O(N__4760),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_6 ));
    InMux I__478 (
            .O(N__4757),
            .I(N__4754));
    LocalMux I__477 (
            .O(N__4754),
            .I(\U712_CHIP_RAM.N_103_0 ));
    InMux I__476 (
            .O(N__4751),
            .I(N__4741));
    InMux I__475 (
            .O(N__4750),
            .I(N__4741));
    InMux I__474 (
            .O(N__4749),
            .I(N__4736));
    InMux I__473 (
            .O(N__4748),
            .I(N__4736));
    InMux I__472 (
            .O(N__4747),
            .I(N__4731));
    InMux I__471 (
            .O(N__4746),
            .I(N__4731));
    LocalMux I__470 (
            .O(N__4741),
            .I(U712_REG_SM_STATE_COUNT_8));
    LocalMux I__469 (
            .O(N__4736),
            .I(U712_REG_SM_STATE_COUNT_8));
    LocalMux I__468 (
            .O(N__4731),
            .I(U712_REG_SM_STATE_COUNT_8));
    CascadeMux I__467 (
            .O(N__4724),
            .I(\U712_CHIP_RAM.N_103_0_cascade_ ));
    InMux I__466 (
            .O(N__4721),
            .I(N__4718));
    LocalMux I__465 (
            .O(N__4718),
            .I(\U712_CHIP_RAM.m106_nsZ0Z_1 ));
    InMux I__464 (
            .O(N__4715),
            .I(N__4712));
    LocalMux I__463 (
            .O(N__4712),
            .I(i62_mux));
    InMux I__462 (
            .O(N__4709),
            .I(N__4706));
    LocalMux I__461 (
            .O(N__4706),
            .I(N__4702));
    InMux I__460 (
            .O(N__4705),
            .I(N__4699));
    Span12Mux_h I__459 (
            .O(N__4702),
            .I(N__4696));
    LocalMux I__458 (
            .O(N__4699),
            .I(N__4693));
    Span12Mux_v I__457 (
            .O(N__4696),
            .I(N__4690));
    Span12Mux_h I__456 (
            .O(N__4693),
            .I(N__4687));
    Odrv12 I__455 (
            .O(N__4690),
            .I(DBRn_c));
    Odrv12 I__454 (
            .O(N__4687),
            .I(DBRn_c));
    InMux I__453 (
            .O(N__4682),
            .I(N__4679));
    LocalMux I__452 (
            .O(N__4679),
            .I(DBR_SYNCZ0Z_0));
    IoInMux I__451 (
            .O(N__4676),
            .I(N__4673));
    LocalMux I__450 (
            .O(N__4673),
            .I(N__4670));
    Odrv12 I__449 (
            .O(N__4670),
            .I(VBENn_c));
    InMux I__448 (
            .O(N__4667),
            .I(N__4663));
    InMux I__447 (
            .O(N__4666),
            .I(N__4660));
    LocalMux I__446 (
            .O(N__4663),
            .I(REG_TACK));
    LocalMux I__445 (
            .O(N__4660),
            .I(REG_TACK));
    InMux I__444 (
            .O(N__4655),
            .I(N__4652));
    LocalMux I__443 (
            .O(N__4652),
            .I(U712_CHIP_RAM_m113_0));
    CascadeMux I__442 (
            .O(N__4649),
            .I(N__4646));
    InMux I__441 (
            .O(N__4646),
            .I(N__4643));
    LocalMux I__440 (
            .O(N__4643),
            .I(\U712_CHIP_RAM.N_87_0 ));
    CascadeMux I__439 (
            .O(N__4640),
            .I(\U712_CHIP_RAM.N_87_0_cascade_ ));
    CascadeMux I__438 (
            .O(N__4637),
            .I(\U712_CHIP_RAM.N_97_0_cascade_ ));
    CascadeMux I__437 (
            .O(N__4634),
            .I(N__4631));
    InMux I__436 (
            .O(N__4631),
            .I(N__4628));
    LocalMux I__435 (
            .O(N__4628),
            .I(N_112_0));
    InMux I__434 (
            .O(N__4625),
            .I(N__4622));
    LocalMux I__433 (
            .O(N__4622),
            .I(U712_REG_SM_REG_TACK_7_0));
    CascadeMux I__432 (
            .O(N__4619),
            .I(N_19_0_cascade_));
    InMux I__431 (
            .O(N__4616),
            .I(N__4608));
    InMux I__430 (
            .O(N__4615),
            .I(N__4608));
    InMux I__429 (
            .O(N__4614),
            .I(N__4603));
    InMux I__428 (
            .O(N__4613),
            .I(N__4603));
    LocalMux I__427 (
            .O(N__4608),
            .I(U712_REG_SM_STATE_COUNT_3));
    LocalMux I__426 (
            .O(N__4603),
            .I(U712_REG_SM_STATE_COUNT_3));
    InMux I__425 (
            .O(N__4598),
            .I(N__4595));
    LocalMux I__424 (
            .O(N__4595),
            .I(N_19_0));
    InMux I__423 (
            .O(N__4592),
            .I(N__4589));
    LocalMux I__422 (
            .O(N__4589),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    IoInMux I__421 (
            .O(N__4586),
            .I(N__4583));
    LocalMux I__420 (
            .O(N__4583),
            .I(N__4580));
    IoSpan4Mux I__419 (
            .O(N__4580),
            .I(N__4577));
    Span4Mux_s3_h I__418 (
            .O(N__4577),
            .I(N__4574));
    Span4Mux_v I__417 (
            .O(N__4574),
            .I(N__4570));
    InMux I__416 (
            .O(N__4573),
            .I(N__4567));
    Span4Mux_h I__415 (
            .O(N__4570),
            .I(N__4564));
    LocalMux I__414 (
            .O(N__4567),
            .I(N__4561));
    Sp12to4 I__413 (
            .O(N__4564),
            .I(N__4558));
    Span4Mux_v I__412 (
            .O(N__4561),
            .I(N__4555));
    Span12Mux_h I__411 (
            .O(N__4558),
            .I(N__4550));
    Sp12to4 I__410 (
            .O(N__4555),
            .I(N__4550));
    Span12Mux_h I__409 (
            .O(N__4550),
            .I(N__4547));
    Odrv12 I__408 (
            .O(N__4547),
            .I(C3_c));
    InMux I__407 (
            .O(N__4544),
            .I(N__4541));
    LocalMux I__406 (
            .O(N__4541),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    IoInMux I__405 (
            .O(N__4538),
            .I(N__4535));
    LocalMux I__404 (
            .O(N__4535),
            .I(N__4532));
    Span4Mux_s3_h I__403 (
            .O(N__4532),
            .I(N__4529));
    Odrv4 I__402 (
            .O(N__4529),
            .I(DBRn_c_i_0));
    IoInMux I__401 (
            .O(N__4526),
            .I(N__4523));
    LocalMux I__400 (
            .O(N__4523),
            .I(N__4520));
    Span4Mux_s2_v I__399 (
            .O(N__4520),
            .I(N__4517));
    Span4Mux_v I__398 (
            .O(N__4517),
            .I(N__4514));
    Odrv4 I__397 (
            .O(N__4514),
            .I(CLK80_PLL_i_i));
    IoInMux I__396 (
            .O(N__4511),
            .I(N__4508));
    LocalMux I__395 (
            .O(N__4508),
            .I(N__4505));
    IoSpan4Mux I__394 (
            .O(N__4505),
            .I(N__4502));
    Span4Mux_s2_v I__393 (
            .O(N__4502),
            .I(N__4499));
    Sp12to4 I__392 (
            .O(N__4499),
            .I(N__4496));
    Span12Mux_v I__391 (
            .O(N__4496),
            .I(N__4493));
    Odrv12 I__390 (
            .O(N__4493),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_A1_nesrC  (
            .O(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .I(N__5001));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .I(N__5004));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .I(N__5006));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .I(N__5008));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .I(N__5009));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .I(N__5003));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .I(N__5005));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ),
            .I(N__5007));
    INV \INVU712_CYCLE_TERM.TACK_OUTC  (
            .O(\INVU712_CYCLE_TERM.TACK_OUTC_net ),
            .I(N__6867));
    INV \INVU712_CYCLE_TERM.TACK_ENC  (
            .O(\INVU712_CYCLE_TERM.TACK_ENC_net ),
            .I(N__6869));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_10_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_14_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_16_0_));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__5293),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__7922),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB DBRn_c_i_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__4538),
            .GLOBALBUFFEROUTPUT(DBRn_c_i_0_g));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__4586),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_2_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_2_11_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_2_11_1  (
            .in0(_gnd_net_),
            .in1(N__6064),
            .in2(_gnd_net_),
            .in3(N__11327),
            .lcout(DBRn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_3_1_5.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_3_1_5.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_3_1_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 CLKRAM_obuf_RNO_LC_3_1_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11474),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBRn_ibuf_RNIBAB_LC_6_13_6.C_ON=1'b0;
    defparam DBRn_ibuf_RNIBAB_LC_6_13_6.SEQ_MODE=4'b0000;
    defparam DBRn_ibuf_RNIBAB_LC_6_13_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 DBRn_ibuf_RNIBAB_LC_6_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4709),
            .lcout(DBRn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_LC_7_11_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_7_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_7_11_0 .LUT_INIT=16'b0101110101010001;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_7_11_0  (
            .in0(N__4625),
            .in1(N__4655),
            .in2(N__4634),
            .in3(N__4666),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11454),
            .ce(),
            .sr(N__11281));
    defparam \U712_CHIP_RAM.m111_LC_7_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m111_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m111_LC_7_12_3 .LUT_INIT=16'b0010110000100000;
    LogicCell40 \U712_CHIP_RAM.m111_LC_7_12_3  (
            .in0(N__4748),
            .in1(N__5700),
            .in2(N__9458),
            .in3(N__4613),
            .lcout(N_112_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m101_LC_7_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m101_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m101_LC_7_12_5 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \U712_CHIP_RAM.m101_LC_7_12_5  (
            .in0(N__4749),
            .in1(N__4614),
            .in2(_gnd_net_),
            .in3(N__4955),
            .lcout(U712_REG_SM_REG_TACK_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m18_LC_7_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m18_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m18_LC_7_13_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.m18_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__5683),
            .in2(_gnd_net_),
            .in3(N__9452),
            .lcout(N_19_0),
            .ltout(N_19_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_7_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_7_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_7_13_1 .LUT_INIT=16'b0100110000001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_7_13_1  (
            .in0(N__4616),
            .in1(N__8109),
            .in2(N__4619),
            .in3(N__4757),
            .lcout(U712_REG_SM_STATE_COUNT_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11461),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_7_13_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_7_13_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_7_13_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_7_13_2  (
            .in0(N__8110),
            .in1(N__4615),
            .in2(_gnd_net_),
            .in3(N__4598),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11461),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_5_LC_7_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_7_13_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_7_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_5_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(N__8111),
            .in2(_gnd_net_),
            .in3(N__4592),
            .lcout(U712_REG_SM_STATE_COUNT_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11461),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_0_LC_7_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_7_14_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_7_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_7_14_1  (
            .in0(N__4573),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11464),
            .ce(),
            .sr(N__11267));
    defparam \U712_REG_SM.C3_SYNC_1_LC_7_14_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_7_14_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_7_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_7_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4544),
            .lcout(U712_REG_SM_C3_SYNC_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11464),
            .ce(),
            .sr(N__11267));
    defparam DBR_SYNC_1_LC_7_16_1.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_7_16_1.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_7_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_7_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4682),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11468),
            .ce(),
            .sr(N__11262));
    defparam DBR_SYNC_0_LC_7_17_3.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_7_17_3.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_7_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_0_LC_7_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4705),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11470),
            .ce(),
            .sr(N__11258));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNI59L8_LC_8_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNI59L8_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNI59L8_LC_8_5_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNI59L8_LC_8_5_1  (
            .in0(N__11076),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11122),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_START_LC_8_10_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_START_LC_8_10_4 .SEQ_MODE=4'b1010;
    defparam \U712_CYCLE_TERM.TACK_START_LC_8_10_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_CYCLE_TERM.TACK_START_LC_8_10_4  (
            .in0(N__4667),
            .in1(N__6629),
            .in2(_gnd_net_),
            .in3(N__5479),
            .lcout(\U712_CYCLE_TERM.TACK_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11446),
            .ce(),
            .sr(N__4811));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_8_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_8_11_3 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_8_11_3  (
            .in0(N__5050),
            .in1(N__5065),
            .in2(N__5036),
            .in3(N__5080),
            .lcout(\U712_CHIP_RAM.REFRESH5lt7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m113_0_LC_8_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m113_0_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m113_0_LC_8_12_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.m113_0_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(N__4774),
            .in2(_gnd_net_),
            .in3(N__4799),
            .lcout(U712_CHIP_RAM_m113_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m79_LC_8_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m79_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m79_LC_8_12_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.m79_LC_8_12_7  (
            .in0(N__9440),
            .in1(N__4798),
            .in2(N__5215),
            .in3(N__5699),
            .lcout(U712_REG_SM_STATE_COUNT_0_sqmuxa_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_8_LC_8_13_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_8_LC_8_13_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_8_LC_8_13_0 .LUT_INIT=16'b1000110010001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_8_LC_8_13_0  (
            .in0(N__4805),
            .in1(N__8099),
            .in2(N__4649),
            .in3(N__4751),
            .lcout(U712_REG_SM_STATE_COUNT_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11457),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m86_LC_8_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m86_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m86_LC_8_13_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_CHIP_RAM.m86_LC_8_13_1  (
            .in0(N__5682),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9425),
            .lcout(\U712_CHIP_RAM.N_87_0 ),
            .ltout(\U712_CHIP_RAM.N_87_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m96_LC_8_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m96_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m96_LC_8_13_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U712_CHIP_RAM.m96_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4640),
            .in3(N__4750),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_97_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_8_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_8_13_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_8_13_3 .LUT_INIT=16'b0111011111110101;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_8_13_3  (
            .in0(N__8096),
            .in1(N__4781),
            .in2(N__4637),
            .in3(N__4797),
            .lcout(U712_REG_SM_STATE_COUNT_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11457),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_7_LC_8_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_7_LC_8_13_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_7_LC_8_13_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_7_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__8098),
            .in2(_gnd_net_),
            .in3(N__4763),
            .lcout(U712_REG_SM_STATE_COUNT_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11457),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m20_e_LC_8_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m20_e_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m20_e_LC_8_13_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.m20_e_LC_8_13_5  (
            .in0(_gnd_net_),
            .in1(N__4796),
            .in2(_gnd_net_),
            .in3(N__5207),
            .lcout(\U712_CHIP_RAM.N_332 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m78_LC_8_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m78_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m78_LC_8_13_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.m78_LC_8_13_6  (
            .in0(N__5208),
            .in1(N__5681),
            .in2(_gnd_net_),
            .in3(N__9431),
            .lcout(\U712_CHIP_RAM.N_79_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_6_LC_8_13_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_8_13_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_6_LC_8_13_7  (
            .in0(N__8097),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4775),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11457),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m106_ns_1_LC_8_14_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m106_ns_1_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m106_ns_1_LC_8_14_0 .LUT_INIT=16'b0111011100110011;
    LogicCell40 \U712_CHIP_RAM.m106_ns_1_LC_8_14_0  (
            .in0(N__5666),
            .in1(N__4949),
            .in2(_gnd_net_),
            .in3(N__9414),
            .lcout(\U712_CHIP_RAM.m106_nsZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_8_14_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_8_14_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_8_14_3 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_8_14_3  (
            .in0(N__11109),
            .in1(N__8100),
            .in2(_gnd_net_),
            .in3(N__4715),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11462),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m98_LC_8_14_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m98_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m98_LC_8_14_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \U712_CHIP_RAM.m98_LC_8_14_4  (
            .in0(N__5665),
            .in1(N__5410),
            .in2(N__9439),
            .in3(N__4746),
            .lcout(N_99_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m102_LC_8_14_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m102_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m102_LC_8_14_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.m102_LC_8_14_6  (
            .in0(N__5667),
            .in1(N__9415),
            .in2(N__6440),
            .in3(N__5386),
            .lcout(\U712_CHIP_RAM.N_103_0 ),
            .ltout(\U712_CHIP_RAM.N_103_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m106_ns_LC_8_14_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m106_ns_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m106_ns_LC_8_14_7 .LUT_INIT=16'b1010101100000001;
    LogicCell40 \U712_CHIP_RAM.m106_ns_LC_8_14_7  (
            .in0(N__4747),
            .in1(N__11108),
            .in2(N__4724),
            .in3(N__4721),
            .lcout(i62_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.WRITE_CYCLE_LC_8_15_3 .C_ON=1'b0;
    defparam \U712_REG_SM.WRITE_CYCLE_LC_8_15_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.WRITE_CYCLE_LC_8_15_3 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \U712_REG_SM.WRITE_CYCLE_LC_8_15_3  (
            .in0(N__10792),
            .in1(N__5239),
            .in2(_gnd_net_),
            .in3(N__4953),
            .lcout(U712_REG_SM_WRITE_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11465),
            .ce(),
            .sr(N__11263));
    defparam \U712_REG_SM.PRnW_LC_8_15_4 .C_ON=1'b0;
    defparam \U712_REG_SM.PRnW_LC_8_15_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.PRnW_LC_8_15_4 .LUT_INIT=16'b1111010111001100;
    LogicCell40 \U712_REG_SM.PRnW_LC_8_15_4  (
            .in0(N__4954),
            .in1(N__4915),
            .in2(N__5701),
            .in3(N__5723),
            .lcout(PRnW_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11465),
            .ce(),
            .sr(N__11263));
    defparam DBR_SYNC_RNITKK4_1_LC_8_16_1.C_ON=1'b0;
    defparam DBR_SYNC_RNITKK4_1_LC_8_16_1.SEQ_MODE=4'b0000;
    defparam DBR_SYNC_RNITKK4_1_LC_8_16_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 DBR_SYNC_RNITKK4_1_LC_8_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6406),
            .lcout(DBR_SYNC_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m85_LC_8_16_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m85_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m85_LC_8_16_2 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \U712_CHIP_RAM.m85_LC_8_16_2  (
            .in0(N__9435),
            .in1(N__5411),
            .in2(N__5710),
            .in3(N__4904),
            .lcout(N_86_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_LC_9_5_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_9_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_9_5_6 .LUT_INIT=16'b0000110100001100;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_LC_9_5_6  (
            .in0(N__5465),
            .in1(N__4840),
            .in2(N__5444),
            .in3(N__5495),
            .lcout(TACK_EN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CYCLE_TERM.TACK_ENC_net ),
            .ce(),
            .sr(N__11297));
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_9_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_9_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_1_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11486),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11439),
            .ce(),
            .sr(N__11282));
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_9_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_9_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_2_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4895),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11439),
            .ce(),
            .sr(N__11282));
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_9_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_9_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_3_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4889),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11439),
            .ce(),
            .sr(N__11282));
    defparam \U712_CYCLE_TERM.TACK_START_RNO_0_LC_9_10_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_START_RNO_0_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_START_RNO_0_LC_9_10_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_START_RNO_0_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(N__8095),
            .in2(_gnd_net_),
            .in3(N__4841),
            .lcout(\U712_CYCLE_TERM.TACK_RST_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_11_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_11_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__5090),
            .in2(_gnd_net_),
            .in3(N__5084),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__5002),
            .ce(),
            .sr(N__7118));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_11_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_11_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(N__5081),
            .in2(_gnd_net_),
            .in3(N__5069),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__5002),
            .ce(),
            .sr(N__7118));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_11_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_11_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(N__5066),
            .in2(_gnd_net_),
            .in3(N__5054),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__5002),
            .ce(),
            .sr(N__7118));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_11_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_11_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__5051),
            .in2(_gnd_net_),
            .in3(N__5039),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__5002),
            .ce(),
            .sr(N__7118));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_11_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_11_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(N__5035),
            .in2(_gnd_net_),
            .in3(N__5021),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__5002),
            .ce(),
            .sr(N__7118));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_11_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_11_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_11_5  (
            .in0(_gnd_net_),
            .in1(N__6247),
            .in2(_gnd_net_),
            .in3(N__5018),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__5002),
            .ce(),
            .sr(N__7118));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_11_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_11_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(N__6263),
            .in2(_gnd_net_),
            .in3(N__5015),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__5002),
            .ce(),
            .sr(N__7118));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_11_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_11_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_11_7  (
            .in0(_gnd_net_),
            .in1(N__6232),
            .in2(_gnd_net_),
            .in3(N__5012),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5002),
            .ce(),
            .sr(N__7118));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_12_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_12_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_12_2 .LUT_INIT=16'b0101000001110011;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_9_12_2  (
            .in0(N__5189),
            .in1(N__4976),
            .in2(N__5216),
            .in3(N__5137),
            .lcout(U712_REG_SM_REG_CYCLE_START),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11450),
            .ce(),
            .sr(N__11268));
    defparam \U712_REG_SM.START_RST_LC_9_12_3 .C_ON=1'b0;
    defparam \U712_REG_SM.START_RST_LC_9_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.START_RST_LC_9_12_3 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \U712_REG_SM.START_RST_LC_9_12_3  (
            .in0(N__5238),
            .in1(N__5188),
            .in2(_gnd_net_),
            .in3(N__5417),
            .lcout(U712_REG_SM_START_RST),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11450),
            .ce(),
            .sr(N__11268));
    defparam \U712_CHIP_RAM.RAS_SYNC_5_LC_9_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_5_LC_9_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_5_LC_9_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_5_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5102),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11450),
            .ce(),
            .sr(N__11268));
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_9_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_9_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_9_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_4_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5180),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11450),
            .ce(),
            .sr(N__11268));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_12_7 .LUT_INIT=16'b0011011100000101;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_12_7  (
            .in0(N__5171),
            .in1(N__10992),
            .in2(N__5138),
            .in3(N__5798),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11450),
            .ce(),
            .sr(N__11268));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIBFJU_LC_9_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIBFJU_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIBFJU_LC_9_13_0 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIBFJU_LC_9_13_0  (
            .in0(N__7279),
            .in1(_gnd_net_),
            .in2(N__8882),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_363 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIPMTA2_LC_9_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIPMTA2_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIPMTA2_LC_9_13_1 .LUT_INIT=16'b0100010001110100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIPMTA2_LC_9_13_1  (
            .in0(N__8664),
            .in1(N__7280),
            .in2(N__6374),
            .in3(N__7103),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m223_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRTQU5_3_LC_9_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRTQU5_3_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRTQU5_3_LC_9_13_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIRTQU5_3_LC_9_13_2  (
            .in0(N__7325),
            .in1(N__7748),
            .in2(N__5111),
            .in3(N__7681),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_9_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_9_13_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_9_13_3  (
            .in0(N__5108),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5101),
            .lcout(\U712_CHIP_RAM.m231_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_9_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_9_13_4 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_9_13_4  (
            .in0(N__8841),
            .in1(N__9124),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_364 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_14_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5258),
            .lcout(U712_REG_SM_C1_SYNC_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11458),
            .ce(),
            .sr(N__11264));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_14_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_14_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_14_4 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_9_14_4  (
            .in0(N__5246),
            .in1(N__5779),
            .in2(_gnd_net_),
            .in3(N__7564),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11458),
            .ce(),
            .sr(N__11264));
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_14_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_14_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5294),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11458),
            .ce(),
            .sr(N__11264));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_14_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_14_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_14_6 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_14_6  (
            .in0(N__8155),
            .in1(N__7282),
            .in2(N__10352),
            .in3(N__5252),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11458),
            .ce(),
            .sr(N__11264));
    defparam \U712_CHIP_RAM.m77_LC_9_15_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m77_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m77_LC_9_15_0 .LUT_INIT=16'b0000111100001101;
    LogicCell40 \U712_CHIP_RAM.m77_LC_9_15_0  (
            .in0(N__10155),
            .in1(N__10794),
            .in2(N__9450),
            .in3(N__5732),
            .lcout(U712_REG_SM_UDSn_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_15_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_15_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_15_2  (
            .in0(N__7840),
            .in1(N__10793),
            .in2(_gnd_net_),
            .in3(N__7281),
            .lcout(\U712_CHIP_RAM.N_236 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m82_LC_9_15_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m82_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m82_LC_9_15_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.m82_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__5705),
            .in2(_gnd_net_),
            .in3(N__9426),
            .lcout(\U712_CHIP_RAM.N_83_0 ),
            .ltout(\U712_CHIP_RAM.N_83_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_9_15_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_9_15_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_9_15_4 .LUT_INIT=16'b0000101010001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_9_15_4  (
            .in0(N__8085),
            .in1(N__5240),
            .in2(N__5219),
            .in3(N__5415),
            .lcout(U712_REG_SM_STATE_COUNT_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11463),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m93_LC_9_15_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m93_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m93_LC_9_15_5 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \U712_CHIP_RAM.m93_LC_9_15_5  (
            .in0(N__5387),
            .in1(N__9430),
            .in2(N__5711),
            .in3(N__6441),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_94_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_9_15_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_9_15_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_9_15_6 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_9_15_6  (
            .in0(N__8086),
            .in1(N__5426),
            .in2(N__5420),
            .in3(N__5416),
            .lcout(U712_REG_SM_STATE_COUNT_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11463),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_9_16_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_9_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(N__6385),
            .in2(N__5374),
            .in3(N__5375),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_9_16_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_9_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__5320),
            .in2(_gnd_net_),
            .in3(N__5357),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_9_16_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_9_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__5332),
            .in2(_gnd_net_),
            .in3(N__5354),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_9_16_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_9_16_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(N__5302),
            .in2(_gnd_net_),
            .in3(N__5351),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_1_LC_9_16_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_1_LC_9_16_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_1_LC_9_16_4 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_1_LC_9_16_4  (
            .in0(N__8112),
            .in1(N__5348),
            .in2(N__8156),
            .in3(N__6439),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11466),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_2_LC_9_16_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_2_LC_9_16_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_2_LC_9_16_5 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_2_LC_9_16_5  (
            .in0(N__6437),
            .in1(N__8113),
            .in2(N__5342),
            .in3(N__8152),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11466),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_9_16_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_9_16_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_9_16_6  (
            .in0(N__5303),
            .in1(N__5333),
            .in2(N__5324),
            .in3(N__6386),
            .lcout(\U712_CHIP_RAM.N_330 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_3_LC_9_16_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_3_LC_9_16_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_3_LC_9_16_7 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_3_LC_9_16_7  (
            .in0(N__6438),
            .in1(N__8114),
            .in2(N__5312),
            .in3(N__8153),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11466),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m6_LC_9_17_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m6_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m6_LC_9_17_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \U712_CHIP_RAM.m6_LC_9_17_3  (
            .in0(N__10077),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9987),
            .lcout(\U712_CHIP_RAM.N_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REGENn_ess_RNO_LC_9_17_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_ess_RNO_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REGENn_ess_RNO_LC_9_17_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.REGENn_ess_RNO_LC_9_17_4  (
            .in0(_gnd_net_),
            .in1(N__11324),
            .in2(_gnd_net_),
            .in3(N__5722),
            .lcout(\U712_REG_SM.N_86_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REGENn_ess_LC_9_18_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_ess_LC_9_18_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_ess_LC_9_18_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_REG_SM.REGENn_ess_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(N__5709),
            .in2(_gnd_net_),
            .in3(N__9451),
            .lcout(BLSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11469),
            .ce(N__5582),
            .sr(N__11246));
    defparam \U712_CYCLE_TERM.TACK_OUT_RNO_0_LC_10_5_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUT_RNO_0_LC_10_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_OUT_RNO_0_LC_10_5_1 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUT_RNO_0_LC_10_5_1  (
            .in0(N__5439),
            .in1(N__5461),
            .in2(_gnd_net_),
            .in3(N__5493),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_36_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_OUT_LC_10_5_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUT_LC_10_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_OUT_LC_10_5_2 .LUT_INIT=16'b1011111110110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUT_LC_10_5_2  (
            .in0(N__5464),
            .in1(N__8080),
            .in2(N__5567),
            .in3(N__5516),
            .lcout(TACK_OUT),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CYCLE_TERM.TACK_OUTC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_10_5_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_10_5_3 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_10_5_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_10_5_3  (
            .in0(N__5440),
            .in1(N__5463),
            .in2(N__8108),
            .in3(N__5494),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CYCLE_TERM.TACK_OUTC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_10_5_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_10_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_10_5_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_10_5_6  (
            .in0(N__5462),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8084),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CYCLE_TERM.TACK_OUTC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIEG6A1_LC_10_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIEG6A1_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIEG6A1_LC_10_9_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIEG6A1_LC_10_9_2  (
            .in0(N__8039),
            .in1(N__9130),
            .in2(_gnd_net_),
            .in3(N__8640),
            .lcout(\U712_CHIP_RAM.m38_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_10_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_10_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_10_10_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_LC_10_10_0  (
            .in0(_gnd_net_),
            .in1(N__7335),
            .in2(_gnd_net_),
            .in3(N__6980),
            .lcout(\U712_CHIP_RAM.CPU_CYCLEm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11440),
            .ce(N__5759),
            .sr(N__11275));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_11_0 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_11_0  (
            .in0(N__8886),
            .in1(N__6975),
            .in2(N__5939),
            .in3(N__9086),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_11_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_11_1  (
            .in0(N__11325),
            .in1(_gnd_net_),
            .in2(N__5762),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIIHAH6_LC_10_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIIHAH6_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIIHAH6_LC_10_11_2 .LUT_INIT=16'b0000000111111011;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIIHAH6_LC_10_11_2  (
            .in0(N__7303),
            .in1(N__7067),
            .in2(N__5807),
            .in3(N__7018),
            .lcout(\U712_CHIP_RAM.m64_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_10_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_10_11_3 .LUT_INIT=16'b1100000011100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_10_11_3  (
            .in0(N__7068),
            .in1(N__8887),
            .in2(N__7823),
            .in3(N__8666),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFK326_0_LC_10_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFK326_0_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFK326_0_LC_10_11_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIFK326_0_LC_10_11_4  (
            .in0(N__8665),
            .in1(N__8772),
            .in2(_gnd_net_),
            .in3(N__7017),
            .lcout(\U712_CHIP_RAM.N_146_0 ),
            .ltout(\U712_CHIP_RAM.N_146_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_11_5 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_11_5  (
            .in0(N__7680),
            .in1(N__8888),
            .in2(N__5747),
            .in3(N__8667),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_11_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_11_6  (
            .in0(_gnd_net_),
            .in1(N__9087),
            .in2(N__5744),
            .in3(N__5741),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_154_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_11_7 .LUT_INIT=16'b1101111101010111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_11_7  (
            .in0(N__7963),
            .in1(N__7139),
            .in2(N__5735),
            .in3(N__11984),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11444),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIRHVM3_LC_10_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIRHVM3_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIRHVM3_LC_10_12_0 .LUT_INIT=16'b1111000100000000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIRHVM3_LC_10_12_0  (
            .in0(N__7094),
            .in1(N__5797),
            .in2(N__6125),
            .in3(N__8771),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_34_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIKHPV5_LC_10_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIKHPV5_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIKHPV5_LC_10_12_1 .LUT_INIT=16'b0101111111111111;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIKHPV5_LC_10_12_1  (
            .in0(N__5819),
            .in1(_gnd_net_),
            .in2(N__5810),
            .in3(N__7042),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_10_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_10_12_2 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_10_12_2  (
            .in0(N__7093),
            .in1(N__6121),
            .in2(_gnd_net_),
            .in3(N__5795),
            .lcout(\U712_CHIP_RAM.N_359 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNI1EAT_LC_10_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNI1EAT_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNI1EAT_LC_10_12_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNI1EAT_LC_10_12_4  (
            .in0(N__8585),
            .in1(N__6120),
            .in2(_gnd_net_),
            .in3(N__5796),
            .lcout(\U712_CHIP_RAM.m41_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_12_7 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_12_7  (
            .in0(N__5924),
            .in1(N__8047),
            .in2(N__5900),
            .in3(N__5780),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11447),
            .ce(N__5850),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_13_1 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_13_1  (
            .in0(N__8057),
            .in1(N__6185),
            .in2(N__8702),
            .in3(N__5893),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11451),
            .ce(N__5855),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_3_LC_10_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_3_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_3_LC_10_13_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_3_LC_10_13_2  (
            .in0(N__8593),
            .in1(N__7746),
            .in2(_gnd_net_),
            .in3(N__7799),
            .lcout(\U712_CHIP_RAM.N_28_0 ),
            .ltout(\U712_CHIP_RAM.N_28_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIBDIU5_3_LC_10_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIBDIU5_3_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIBDIU5_3_LC_10_13_3 .LUT_INIT=16'b0100011111001111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIBDIU5_3_LC_10_13_3  (
            .in0(N__7747),
            .in1(N__9125),
            .in2(N__5768),
            .in3(N__6488),
            .lcout(\U712_CHIP_RAM.m66_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_13_4 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_13_4  (
            .in0(N__8594),
            .in1(N__8873),
            .in2(N__7578),
            .in3(N__7800),
            .lcout(\U712_CHIP_RAM.N_353_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIA1VV6_1_LC_10_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIA1VV6_1_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIA1VV6_1_LC_10_13_6 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIA1VV6_1_LC_10_13_6  (
            .in0(N__8595),
            .in1(N__8874),
            .in2(N__8784),
            .in3(N__6201),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_47_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIAEA2H_LC_10_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIAEA2H_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIAEA2H_LC_10_13_7 .LUT_INIT=16'b1111110101110101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIAEA2H_LC_10_13_7  (
            .in0(N__8056),
            .in1(N__9126),
            .in2(N__5765),
            .in3(N__6500),
            .lcout(\U712_CHIP_RAM.N_56_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_14_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_14_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(N__8589),
            .in2(_gnd_net_),
            .in3(N__6517),
            .lcout(\U712_CHIP_RAM.N_215 ),
            .ltout(),
            .carryin(bfn_10_14_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_14_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_14_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_14_1  (
            .in0(N__5889),
            .in1(N__8872),
            .in2(_gnd_net_),
            .in3(N__5927),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(N__11455),
            .ce(N__5854),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_14_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(N__6557),
            .in2(_gnd_net_),
            .in3(N__5915),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_14_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_14_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_14_3  (
            .in0(N__5890),
            .in1(N__7749),
            .in2(_gnd_net_),
            .in3(N__5912),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__11455),
            .ce(N__5854),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_14_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_14_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_14_4  (
            .in0(N__5887),
            .in1(N__6586),
            .in2(_gnd_net_),
            .in3(N__5909),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__11455),
            .ce(N__5854),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_14_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_14_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_14_5  (
            .in0(N__5891),
            .in1(N__6599),
            .in2(_gnd_net_),
            .in3(N__5906),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__11455),
            .ce(N__5854),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_14_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_14_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_14_6  (
            .in0(N__5888),
            .in1(N__6611),
            .in2(_gnd_net_),
            .in3(N__5903),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__11455),
            .ce(N__5854),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_14_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_14_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_14_7  (
            .in0(N__5892),
            .in1(N__6572),
            .in2(_gnd_net_),
            .in3(N__5858),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11455),
            .ce(N__5854),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_10_15_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_10_15_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_10_15_0 .LUT_INIT=16'b1010101001110111;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_10_15_0  (
            .in0(N__8154),
            .in1(N__5825),
            .in2(_gnd_net_),
            .in3(N__6442),
            .lcout(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11459),
            .ce(),
            .sr(N__11255));
    defparam \U712_REG_SM.UDSn_LC_10_15_5 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_LC_10_15_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.UDSn_LC_10_15_5 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \U712_REG_SM.UDSn_LC_10_15_5  (
            .in0(N__6082),
            .in1(N__6104),
            .in2(_gnd_net_),
            .in3(N__8209),
            .lcout(UDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11459),
            .ce(),
            .sr(N__11255));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_11_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_11_6_2 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_11_6_2  (
            .in0(N__6071),
            .in1(N__11845),
            .in2(N__11789),
            .in3(N__5959),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ),
            .ce(),
            .sr(N__11286));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_11_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_11_7_1 .LUT_INIT=16'b1111101100000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_11_7_1  (
            .in0(N__9617),
            .in1(N__12214),
            .in2(N__11044),
            .in3(N__5945),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11428),
            .ce(N__9646),
            .sr(N__11283));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_8_1 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_8_1  (
            .in0(N__6019),
            .in1(N__12123),
            .in2(N__8369),
            .in3(N__10939),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m186_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_11_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_11_8_2 .LUT_INIT=16'b1011000000010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_11_8_2  (
            .in0(N__8294),
            .in1(N__6173),
            .in2(N__5984),
            .in3(N__10478),
            .lcout(\U712_CHIP_RAM.m186_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_11_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_11_8_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(N__10937),
            .in2(_gnd_net_),
            .in3(N__12122),
            .lcout(\U712_CHIP_RAM.m186_m2_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_11_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_11_8_6 .LUT_INIT=16'b0000000011011111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_11_8_6  (
            .in0(N__10938),
            .in1(N__5981),
            .in2(N__12182),
            .in3(N__8354),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m192_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_11_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_11_8_7 .LUT_INIT=16'b1101000000010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_11_8_7  (
            .in0(N__6179),
            .in1(N__8295),
            .in2(N__5963),
            .in3(N__5960),
            .lcout(\U712_CHIP_RAM.m192_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_8_LC_11_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_8_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_8_LC_11_9_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_8_LC_11_9_0  (
            .in0(N__12120),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6278),
            .lcout(\U712_CHIP_RAM.d_N_6_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_0_LC_11_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_0_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_0_LC_11_9_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_0_LC_11_9_2  (
            .in0(N__12121),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6314),
            .lcout(\U712_CHIP_RAM.d_N_6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNILLSM_0_LC_11_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNILLSM_0_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNILLSM_0_LC_11_9_7 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNILLSM_0_LC_11_9_7  (
            .in0(N__9221),
            .in1(N__12119),
            .in2(N__9873),
            .in3(N__10915),
            .lcout(\U712_CHIP_RAM.m184_m2_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_11_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_11_10_0 .LUT_INIT=16'b1010001110100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_11_10_0  (
            .in0(N__6167),
            .in1(N__8671),
            .in2(N__9120),
            .in3(N__8786),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_168_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_10_1 .LUT_INIT=16'b1101111101010111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_10_1  (
            .in0(N__8037),
            .in1(N__7136),
            .in2(N__6158),
            .in3(N__9884),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11437),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIO6RP9_3_LC_11_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIO6RP9_3_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIO6RP9_3_LC_11_10_2 .LUT_INIT=16'b1011000100010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIO6RP9_3_LC_11_10_2  (
            .in0(N__8668),
            .in1(N__6155),
            .in2(N__7772),
            .in3(N__7679),
            .lcout(),
            .ltout(\U712_CHIP_RAM.i67_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNISRNIG_LC_11_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNISRNIG_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNISRNIG_LC_11_10_3 .LUT_INIT=16'b0100000011101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNISRNIG_LC_11_10_3  (
            .in0(N__8914),
            .in1(N__9088),
            .in2(N__6149),
            .in3(N__6146),
            .lcout(\U712_CHIP_RAM.N_67_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_11_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_11_10_4 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_11_10_4  (
            .in0(N__8670),
            .in1(N__6137),
            .in2(N__7685),
            .in3(N__8915),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_11_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_11_10_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(N__9089),
            .in2(N__6131),
            .in3(N__6338),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_151_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_10_6 .LUT_INIT=16'b1011111100110111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_10_6  (
            .in0(N__7137),
            .in1(N__8038),
            .in2(N__6128),
            .in3(N__9233),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11437),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_11_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_11_10_7 .LUT_INIT=16'b1010000001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_11_10_7  (
            .in0(N__8913),
            .in1(N__7070),
            .in2(N__7816),
            .in3(N__8669),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_0_LC_11_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_0_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_0_LC_11_11_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_0_LC_11_11_2  (
            .in0(N__6332),
            .in1(N__6313),
            .in2(_gnd_net_),
            .in3(N__8977),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11441),
            .ce(),
            .sr(N__11265));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_11_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_11_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_11_11_3 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_11_11_3  (
            .in0(N__8978),
            .in1(N__6299),
            .in2(N__11782),
            .in3(N__6277),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11441),
            .ce(),
            .sr(N__11265));
    defparam \U712_CHIP_RAM.REFRESH_LC_11_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_11_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_11_11_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_11_11_5  (
            .in0(N__6262),
            .in1(N__6248),
            .in2(N__6233),
            .in3(N__6215),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11441),
            .ce(),
            .sr(N__11265));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_11_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_11_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_11_11_7 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_11_11_7  (
            .in0(N__9102),
            .in1(N__8923),
            .in2(_gnd_net_),
            .in3(N__6206),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11441),
            .ce(),
            .sr(N__11265));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_12_0 .LUT_INIT=16'b1100101011000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_12_0  (
            .in0(N__8885),
            .in1(N__6350),
            .in2(N__9121),
            .in3(N__6202),
            .lcout(\U712_CHIP_RAM.N_219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIA7LA2_3_LC_11_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIA7LA2_3_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIA7LA2_3_LC_11_12_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIA7LA2_3_LC_11_12_1  (
            .in0(N__6483),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7750),
            .lcout(\U712_CHIP_RAM.N_48_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_2_LC_11_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_2_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_2_LC_11_12_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_2_LC_11_12_2  (
            .in0(N__7752),
            .in1(N__6556),
            .in2(_gnd_net_),
            .in3(N__6484),
            .lcout(\U712_CHIP_RAM.N_31_0 ),
            .ltout(\U712_CHIP_RAM.N_31_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNI50JL4_LC_11_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNI50JL4_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNI50JL4_LC_11_12_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNI50JL4_LC_11_12_3  (
            .in0(N__7297),
            .in1(N__6367),
            .in2(N__6356),
            .in3(N__7096),
            .lcout(\U712_CHIP_RAM.N_43_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_0_2_LC_11_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_0_2_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_0_2_LC_11_12_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_0_2_LC_11_12_4  (
            .in0(N__7751),
            .in1(N__6555),
            .in2(_gnd_net_),
            .in3(N__6482),
            .lcout(\U712_CHIP_RAM.N_58_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_3_LC_11_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_3_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_3_LC_11_12_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_3_LC_11_12_5  (
            .in0(N__7802),
            .in1(N__8639),
            .in2(_gnd_net_),
            .in3(N__7756),
            .lcout(\U712_CHIP_RAM.CLK_EN_RNOZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_3_0_LC_11_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_3_0_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_3_0_LC_11_12_6 .LUT_INIT=16'b0010011100100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_3_0_LC_11_12_6  (
            .in0(N__8883),
            .in1(N__6518),
            .in2(N__7766),
            .in3(N__7801),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m217_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_11_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_11_12_7 .LUT_INIT=16'b1001110000010100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_11_12_7  (
            .in0(N__8625),
            .in1(N__8884),
            .in2(N__6353),
            .in3(N__7505),
            .lcout(\U712_CHIP_RAM.N_218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_11_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_11_13_0 .LUT_INIT=16'b0010111100001111;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_11_13_0  (
            .in0(N__10994),
            .in1(N__8628),
            .in2(N__8899),
            .in3(N__7024),
            .lcout(\U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_11_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_11_13_1 .LUT_INIT=16'b0000011000000100;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_11_13_1  (
            .in0(N__8627),
            .in1(N__8867),
            .in2(N__7586),
            .in3(N__10993),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m212_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_13_2 .LUT_INIT=16'b1111100000001000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_13_2  (
            .in0(N__8871),
            .in1(N__7023),
            .in2(N__6344),
            .in3(N__7524),
            .lcout(\U712_CHIP_RAM.N_213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI96LA2_0_2_LC_11_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI96LA2_0_2_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI96LA2_0_2_LC_11_13_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI96LA2_0_2_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__6545),
            .in2(_gnd_net_),
            .in3(N__6481),
            .lcout(\U712_CHIP_RAM.N_30_0 ),
            .ltout(\U712_CHIP_RAM.N_30_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_13_4 .LUT_INIT=16'b0110010000100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_13_4  (
            .in0(N__8866),
            .in1(N__8626),
            .in2(N__6341),
            .in3(N__7022),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_11_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_11_13_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_11_13_5 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_11_13_5  (
            .in0(N__6622),
            .in1(N__6641),
            .in2(N__9131),
            .in3(N__6635),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11448),
            .ce(),
            .sr(N__11259));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_13_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_13_6  (
            .in0(N__6610),
            .in1(N__6598),
            .in2(N__6587),
            .in3(N__6571),
            .lcout(\U712_CHIP_RAM.N_333_mux ),
            .ltout(\U712_CHIP_RAM.N_333_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI96LA2_2_LC_11_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI96LA2_2_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI96LA2_2_LC_11_13_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI96LA2_2_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6560),
            .in3(N__6544),
            .lcout(\U712_CHIP_RAM.N_26_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNI2E2T2_LC_11_14_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNI2E2T2_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNI2E2T2_LC_11_14_0 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNI2E2T2_LC_11_14_0  (
            .in0(N__7724),
            .in1(N__6554),
            .in2(N__7579),
            .in3(N__6485),
            .lcout(\U712_CHIP_RAM.N_51_0 ),
            .ltout(\U712_CHIP_RAM.N_51_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFI279_1_LC_11_14_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFI279_1_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFI279_1_LC_11_14_1 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIFI279_1_LC_11_14_1  (
            .in0(N__8846),
            .in1(N__6494),
            .in2(N__6503),
            .in3(N__7499),
            .lcout(\U712_CHIP_RAM.N_54_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_11_14_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_11_14_2 .LUT_INIT=16'b0000110100001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_11_14_2  (
            .in0(N__7726),
            .in1(N__8845),
            .in2(N__8641),
            .in3(N__6487),
            .lcout(\U712_CHIP_RAM.m53_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_RNIAPHI2_LC_11_14_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_RNIAPHI2_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_RNIAPHI2_LC_11_14_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_RNIAPHI2_LC_11_14_5  (
            .in0(N__6486),
            .in1(N__10337),
            .in2(_gnd_net_),
            .in3(N__7725),
            .lcout(\U712_CHIP_RAM.N_52_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_0_LC_11_16_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_0_LC_11_16_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_0_LC_11_16_7 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_0_LC_11_16_7  (
            .in0(N__8094),
            .in1(N__6452),
            .in2(N__8148),
            .in3(N__6443),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11460),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_12_4_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_12_4_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_12_4_0 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_12_4_0  (
            .in0(N__11071),
            .in1(N__9803),
            .in2(N__12228),
            .in3(N__6704),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11424),
            .ce(N__9666),
            .sr(N__11291));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_4_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_4_2 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_12_4_2  (
            .in0(N__11070),
            .in1(N__9308),
            .in2(N__12227),
            .in3(N__6698),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11424),
            .ce(N__9666),
            .sr(N__11291));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_4_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_4_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_12_4_5  (
            .in0(N__8370),
            .in1(N__12014),
            .in2(_gnd_net_),
            .in3(N__12199),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11424),
            .ce(N__9666),
            .sr(N__11291));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_5_0 .LUT_INIT=16'b1101000000010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_5_0  (
            .in0(N__6662),
            .in1(N__8303),
            .in2(N__6959),
            .in3(N__9707),
            .lcout(\U712_CHIP_RAM.m189_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_5_5 .LUT_INIT=16'b1100010000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_5_5  (
            .in0(N__6692),
            .in1(N__6668),
            .in2(N__8306),
            .in3(N__9752),
            .lcout(\U712_CHIP_RAM.m188_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_6_0 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_6_0  (
            .in0(N__9242),
            .in1(N__12183),
            .in2(N__9892),
            .in3(N__7364),
            .lcout(\U712_CHIP_RAM.d_N_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_3_LC_12_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_3_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_3_LC_12_6_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_3_LC_12_6_1  (
            .in0(N__12185),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7430),
            .lcout(\U712_CHIP_RAM.d_N_6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_12_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_12_6_2 .LUT_INIT=16'b0000000011011111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_12_6_2  (
            .in0(N__11045),
            .in1(N__6686),
            .in2(N__12225),
            .in3(N__8360),
            .lcout(\U712_CHIP_RAM.m188_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_4_LC_12_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_4_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_4_LC_12_6_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_4_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(N__12184),
            .in2(_gnd_net_),
            .in3(N__7397),
            .lcout(\U712_CHIP_RAM.d_N_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_6_6 .LUT_INIT=16'b0000000010111111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_6_6  (
            .in0(N__6656),
            .in1(N__11060),
            .in2(N__12226),
            .in3(N__8361),
            .lcout(\U712_CHIP_RAM.m189_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_6_7 .LUT_INIT=16'b1100010011000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_6_7  (
            .in0(N__6950),
            .in1(N__12186),
            .in2(N__8371),
            .in3(N__11046),
            .lcout(\U712_CHIP_RAM.m185_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_7_1 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_12_7_1  (
            .in0(N__11000),
            .in1(N__9608),
            .in2(N__12242),
            .in3(N__6776),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11427),
            .ce(N__9645),
            .sr(N__11278));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_12_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_12_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_12_7_5 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_12_7_5  (
            .in0(N__10998),
            .in1(N__10463),
            .in2(N__12240),
            .in3(N__6911),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11427),
            .ce(N__9645),
            .sr(N__11278));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_7_7 .LUT_INIT=16'b0000000011101111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_12_7_7  (
            .in0(N__10999),
            .in1(N__10589),
            .in2(N__12241),
            .in3(N__8399),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11427),
            .ce(N__9645),
            .sr(N__11278));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_8_2 .LUT_INIT=16'b0000011000000111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_8_2  (
            .in0(N__9234),
            .in1(N__12148),
            .in2(N__12006),
            .in3(N__9880),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_198_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_8_3 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_8_3  (
            .in0(N__11326),
            .in1(_gnd_net_),
            .in2(N__6872),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_198_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLK40_PLL_derived_clock_RNIIOT_LC_12_8_5.C_ON=1'b0;
    defparam CLK40_PLL_derived_clock_RNIIOT_LC_12_8_5.SEQ_MODE=4'b0000;
    defparam CLK40_PLL_derived_clock_RNIIOT_LC_12_8_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLK40_PLL_derived_clock_RNIIOT_LC_12_8_5 (
            .in0(N__6868),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK40_PLL_iso_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_8_7 .LUT_INIT=16'b1100010000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_8_7  (
            .in0(N__6989),
            .in1(N__7160),
            .in2(N__8304),
            .in3(N__9599),
            .lcout(\U712_CHIP_RAM.m187_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_9_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__9220),
            .in2(_gnd_net_),
            .in3(N__9855),
            .lcout(\U712_CHIP_RAM.N_3_0 ),
            .ltout(\U712_CHIP_RAM.N_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_9_1 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_9_1  (
            .in0(N__11004),
            .in1(N__7192),
            .in2(N__7163),
            .in3(N__12163),
            .lcout(\U712_CHIP_RAM.m187_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_12_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_12_9_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_12_9_5  (
            .in0(N__9122),
            .in1(N__7154),
            .in2(_gnd_net_),
            .in3(N__6995),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_163_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_12_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_12_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_12_9_6 .LUT_INIT=16'b1011101100111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_12_9_6  (
            .in0(N__12164),
            .in1(N__8061),
            .in2(N__7142),
            .in3(N__7138),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11431),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_12_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_12_10_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_12_10_4  (
            .in0(N__9228),
            .in1(N__9854),
            .in2(N__12181),
            .in3(N__11996),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_12_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_12_10_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_12_10_5  (
            .in0(N__7304),
            .in1(N__7095),
            .in2(_gnd_net_),
            .in3(N__7069),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_158_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_12_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_12_10_6 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_12_10_6  (
            .in0(N__7046),
            .in1(N__8676),
            .in2(N__7028),
            .in3(N__7025),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_2_LC_12_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_2_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_2_LC_12_10_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_2_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(N__12118),
            .in2(_gnd_net_),
            .in3(N__7459),
            .lcout(\U712_CHIP_RAM.d_N_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIU7TF5_LC_12_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIU7TF5_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIU7TF5_LC_12_11_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIU7TF5_LC_12_11_3  (
            .in0(_gnd_net_),
            .in1(N__7336),
            .in2(_gnd_net_),
            .in3(N__6976),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_2_LC_12_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_2_LC_12_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_2_LC_12_11_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_2_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(N__7481),
            .in2(N__7463),
            .in3(N__7460),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11436),
            .ce(),
            .sr(N__11261));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_3_LC_12_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_3_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_3_LC_12_11_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_3_LC_12_11_5  (
            .in0(N__7448),
            .in1(N__7429),
            .in2(_gnd_net_),
            .in3(N__8974),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11436),
            .ce(),
            .sr(N__11261));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_4_LC_12_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_4_LC_12_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_4_LC_12_11_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_4_LC_12_11_6  (
            .in0(N__8975),
            .in1(N__7415),
            .in2(_gnd_net_),
            .in3(N__7393),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11436),
            .ce(),
            .sr(N__11261));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_5_LC_12_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_5_LC_12_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_5_LC_12_11_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_5_LC_12_11_7  (
            .in0(N__7379),
            .in1(N__7360),
            .in2(_gnd_net_),
            .in3(N__8976),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11436),
            .ce(),
            .sr(N__11261));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIJD6O3_LC_12_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIJD6O3_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIJD6O3_LC_12_12_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIJD6O3_LC_12_12_1  (
            .in0(N__7298),
            .in1(N__8681),
            .in2(_gnd_net_),
            .in3(N__8779),
            .lcout(),
            .ltout(\U712_CHIP_RAM.DMA_CYCLE_START_RNIJD6OZ0Z3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ1M5A_1_LC_12_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ1M5A_1_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ1M5A_1_LC_12_12_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ1M5A_1_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__8922),
            .in2(N__7346),
            .in3(N__7640),
            .lcout(\U712_CHIP_RAM.N_204 ),
            .ltout(\U712_CHIP_RAM.N_204_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_12_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_12_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_12_12_3 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_LC_12_12_3  (
            .in0(N__9103),
            .in1(N__7861),
            .in2(N__7343),
            .in3(N__10331),
            .lcout(\U712_CHIP_RAM.DMA_CYCLEm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11438),
            .ce(),
            .sr(N__11257));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_12_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_12_12_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_12_12_4  (
            .in0(N__8780),
            .in1(N__7340),
            .in2(N__8687),
            .in3(N__7299),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBDIR_LC_12_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_12_12_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_12_12_5 .LUT_INIT=16'b0011111100110000;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(N__7849),
            .in2(N__7238),
            .in3(N__7216),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11438),
            .ce(),
            .sr(N__11257));
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_12_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_12_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_12_12_7 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_12_12_7  (
            .in0(N__7862),
            .in1(N__10723),
            .in2(_gnd_net_),
            .in3(N__7850),
            .lcout(\U712_CHIP_RAM.DMA_WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11438),
            .ce(),
            .sr(N__11257));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_12_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_12_13_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_1_LC_12_13_0  (
            .in0(N__8920),
            .in1(N__7771),
            .in2(N__8680),
            .in3(N__7809),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_3_LC_12_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_3_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_3_LC_12_13_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_3_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(N__7770),
            .in2(_gnd_net_),
            .in3(N__7666),
            .lcout(\U712_CHIP_RAM.N_62_0 ),
            .ltout(\U712_CHIP_RAM.N_62_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNI9THU5_LC_12_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNI9THU5_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNI9THU5_LC_12_13_2 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNI9THU5_LC_12_13_2  (
            .in0(N__8653),
            .in1(N__7580),
            .in2(N__7643),
            .in3(N__7503),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_RNI9THUZ0Z5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_2_LC_12_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_2_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_2_LC_12_13_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_2_LC_12_13_3  (
            .in0(N__7582),
            .in1(N__11030),
            .in2(N__7529),
            .in3(N__8658),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CLK_EN_RNOZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_12_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_12_13_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_0_LC_12_13_4  (
            .in0(N__8921),
            .in1(_gnd_net_),
            .in2(N__7634),
            .in3(N__7631),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_174_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_LC_12_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_12_13_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_12_13_5 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_12_13_5  (
            .in0(N__7597),
            .in1(N__9119),
            .in2(N__7622),
            .in3(N__7619),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11443),
            .ce(),
            .sr(N__11254));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_12_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_12_13_6 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_12_13_6  (
            .in0(N__8654),
            .in1(N__7581),
            .in2(N__7528),
            .in3(N__7504),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_208_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_12_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_12_13_7 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(N__8919),
            .in2(N__8213),
            .in3(N__9118),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_ess_RNO_LC_12_14_4 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_12_14_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_REG_SM.ASn_ess_RNO_LC_12_14_4  (
            .in0(N__11323),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8202),
            .lcout(\U712_REG_SM.N_99_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDSn_LC_12_16_5 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_LC_12_16_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.LDSn_LC_12_16_5 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \U712_REG_SM.LDSn_LC_12_16_5  (
            .in0(N__8167),
            .in1(N__9341),
            .in2(_gnd_net_),
            .in3(N__8210),
            .lcout(LDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11453),
            .ce(),
            .sr(N__11245));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_12_17_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_12_17_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_12_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10289),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11456),
            .ce(),
            .sr(N__11244));
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_4.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_4.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8036),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RASn_LC_13_2_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_13_2_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_13_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_13_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9241),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11423),
            .ce(),
            .sr(N__11301));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_13_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_13_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_13_5_5 .LUT_INIT=16'b1100111011111110;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_13_5_5  (
            .in0(N__7892),
            .in1(N__7886),
            .in2(N__8429),
            .in3(N__10601),
            .lcout(\U712_CHIP_RAM.m185_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_13_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_13_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_13_5_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_13_5_7  (
            .in0(_gnd_net_),
            .in1(N__8372),
            .in2(_gnd_net_),
            .in3(N__12230),
            .lcout(\U712_CHIP_RAM.m194_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_6_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_6_3  (
            .in0(N__11846),
            .in1(N__11942),
            .in2(_gnd_net_),
            .in3(N__11746),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .ce(N__11564),
            .sr(N__11287));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_13_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_13_7_2 .LUT_INIT=16'b0011001100010011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_13_7_2  (
            .in0(N__11022),
            .in1(N__8368),
            .in2(N__12229),
            .in3(N__7880),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m191_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_7_3 .LUT_INIT=16'b1101000000010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_7_3  (
            .in0(N__8477),
            .in1(N__8305),
            .in2(N__8486),
            .in3(N__8483),
            .lcout(\U712_CHIP_RAM.m191_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_7_LC_13_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_7_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_7_LC_13_8_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_7_LC_13_8_3  (
            .in0(_gnd_net_),
            .in1(N__9146),
            .in2(_gnd_net_),
            .in3(N__12151),
            .lcout(\U712_CHIP_RAM.d_N_6_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_8_4 .LUT_INIT=16'b1010101000100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_8_4  (
            .in0(N__12152),
            .in1(N__8461),
            .in2(N__11061),
            .in3(N__8355),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m184_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_8_5 .LUT_INIT=16'b1111010011111110;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_8_5  (
            .in0(N__8425),
            .in1(N__9176),
            .in2(N__8402),
            .in3(N__10538),
            .lcout(\U712_CHIP_RAM.m184_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_13_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_13_8_6 .LUT_INIT=16'b0000000011011111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_13_8_6  (
            .in0(N__12153),
            .in1(N__8393),
            .in2(N__11062),
            .in3(N__8356),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m190_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_8_7 .LUT_INIT=16'b1011000000010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_8_7  (
            .in0(N__8299),
            .in1(N__8222),
            .in2(N__8252),
            .in3(N__9590),
            .lcout(\U712_CHIP_RAM.m190_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_13_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_13_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_13_9_5 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_13_9_5  (
            .in0(N__9584),
            .in1(N__11029),
            .in2(N__12224),
            .in3(N__8249),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11435),
            .ce(N__9647),
            .sr(N__11276));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_6_LC_13_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_6_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_6_LC_13_10_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_6_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(N__8935),
            .in2(_gnd_net_),
            .in3(N__12150),
            .lcout(\U712_CHIP_RAM.d_N_6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_10_2 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_10_2  (
            .in0(N__9232),
            .in1(N__12149),
            .in2(N__9891),
            .in3(N__8992),
            .lcout(\U712_CHIP_RAM.d_N_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_13_10_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_13_10_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_13_10_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_13_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_7_LC_13_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_7_LC_13_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_7_LC_13_11_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_7_LC_13_11_2  (
            .in0(N__8981),
            .in1(N__9167),
            .in2(_gnd_net_),
            .in3(N__9145),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11442),
            .ce(),
            .sr(N__11266));
    defparam \U712_CHIP_RAM.DBENn_LC_13_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_13_11_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_13_11_3 .LUT_INIT=16'b0010111010101010;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_13_11_3  (
            .in0(N__10235),
            .in1(N__9123),
            .in2(N__8738),
            .in3(N__9020),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11442),
            .ce(),
            .sr(N__11266));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_1_LC_13_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_1_LC_13_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_1_LC_13_11_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_1_LC_13_11_5  (
            .in0(N__9014),
            .in1(N__8993),
            .in2(_gnd_net_),
            .in3(N__8979),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11442),
            .ce(),
            .sr(N__11266));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_6_LC_13_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_6_LC_13_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_6_LC_13_11_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_6_LC_13_11_6  (
            .in0(N__8980),
            .in1(N__8948),
            .in2(_gnd_net_),
            .in3(N__8936),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11442),
            .ce(),
            .sr(N__11266));
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_13_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_13_12_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNO_0_LC_13_12_0  (
            .in0(N__8924),
            .in1(N__8785),
            .in2(N__8685),
            .in3(N__10364),
            .lcout(\U712_CHIP_RAM.DBENn_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_13_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_13_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_13_12_1  (
            .in0(N__8719),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8672),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_13_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_13_13_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_13_13_6 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_LC_13_13_6  (
            .in0(N__10330),
            .in1(N__8497),
            .in2(N__8686),
            .in3(N__8513),
            .lcout(LATCH_CLK_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11449),
            .ce(),
            .sr(N__11260));
    defparam \U712_REG_SM.ASn_ess_LC_13_14_5 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_LC_13_14_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_ess_LC_13_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.ASn_ess_LC_13_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9457),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11452),
            .ce(N__9470),
            .sr(N__11256));
    defparam \U712_CHIP_RAM.m74_LC_13_16_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m74_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m74_LC_13_16_3 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \U712_CHIP_RAM.m74_LC_13_16_3  (
            .in0(N__9938),
            .in1(N__10801),
            .in2(_gnd_net_),
            .in3(N__9453),
            .lcout(U712_REG_SM_LDSn_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m8_LC_13_17_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m8_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m8_LC_13_17_4 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \U712_CHIP_RAM.m8_LC_13_17_4  (
            .in0(N__9989),
            .in1(_gnd_net_),
            .in2(N__10097),
            .in3(N__10167),
            .lcout(\U712_CHIP_RAM.N_325_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m11_LC_13_17_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m11_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m11_LC_13_17_7 .LUT_INIT=16'b0011000111000100;
    LogicCell40 \U712_CHIP_RAM.m11_LC_13_17_7  (
            .in0(N__10034),
            .in1(N__10090),
            .in2(N__10169),
            .in3(N__9988),
            .lcout(LMBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_14_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_14_4_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_14_4_2 .LUT_INIT=16'b0000000011101111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_14_4_2  (
            .in0(N__9296),
            .in1(N__11043),
            .in2(N__12248),
            .in3(N__9335),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11426),
            .ce(N__9667),
            .sr(N__11298));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_5_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_5_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_5_4  (
            .in0(N__11779),
            .in1(N__10572),
            .in2(_gnd_net_),
            .in3(N__9793),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11602),
            .ce(N__11568),
            .sr(N__11294));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_5_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_5_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_5_5  (
            .in0(N__9743),
            .in1(N__11780),
            .in2(_gnd_net_),
            .in3(N__10630),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11602),
            .ce(N__11568),
            .sr(N__11294));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_6_2 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_14_6_2  (
            .in0(N__9290),
            .in1(N__9269),
            .in2(N__11080),
            .in3(N__11615),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11429),
            .ce(N__9671),
            .sr(N__11292));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_14_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_14_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_14_6_7 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_14_6_7  (
            .in0(N__11855),
            .in1(N__11072),
            .in2(N__12243),
            .in3(N__9698),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11429),
            .ce(N__9671),
            .sr(N__11292));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_7_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_7_4  (
            .in0(N__11828),
            .in1(N__11937),
            .in2(_gnd_net_),
            .in3(N__11706),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11601),
            .ce(N__11565),
            .sr(N__11288));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_7_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_7_6  (
            .in0(N__10529),
            .in1(N__10571),
            .in2(_gnd_net_),
            .in3(N__11705),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11601),
            .ce(N__11565),
            .sr(N__11288));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_8_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_8_3  (
            .in0(N__10580),
            .in1(N__9782),
            .in2(_gnd_net_),
            .in3(N__11751),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__11562),
            .sr(N__11284));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_8_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_8_7  (
            .in0(N__11886),
            .in1(N__11936),
            .in2(_gnd_net_),
            .in3(N__11752),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__11562),
            .sr(N__11284));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_9_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_9_6  (
            .in0(N__10629),
            .in1(N__11750),
            .in2(_gnd_net_),
            .in3(N__11885),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11597),
            .ce(N__11560),
            .sr(N__11279));
    defparam \U712_CHIP_RAM.DBENn_RNI6U6F1_0_LC_14_14_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNI6U6F1_0_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNI6U6F1_0_LC_14_14_1 .LUT_INIT=16'b0100110001011111;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNI6U6F1_0_LC_14_14_1  (
            .in0(N__10280),
            .in1(N__9910),
            .in2(N__10262),
            .in3(N__11063),
            .lcout(CUMBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_RNI8DDB1_LC_14_14_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNI8DDB1_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNI8DDB1_LC_14_14_3 .LUT_INIT=16'b1100010011110101;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNI8DDB1_LC_14_14_3  (
            .in0(N__10298),
            .in1(N__9547),
            .in2(N__10263),
            .in3(N__11066),
            .lcout(CLMBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_RNI8DDB1_0_LC_14_14_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNI8DDB1_0_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNI8DDB1_0_LC_14_14_4 .LUT_INIT=16'b0000110111011101;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNI8DDB1_0_LC_14_14_4  (
            .in0(N__11065),
            .in1(N__10114),
            .in2(N__10264),
            .in3(N__10297),
            .lcout(CUUBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_RNIMKV8_LC_14_14_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_RNIMKV8_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_RNIMKV8_LC_14_14_5 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_RNIMKV8_LC_14_14_5  (
            .in0(N__10856),
            .in1(N__10350),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_346 ),
            .ltout(\U712_CHIP_RAM.N_346_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_RNI6U6F1_LC_14_14_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNI6U6F1_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNI6U6F1_LC_14_14_6 .LUT_INIT=16'b1100111101000101;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNI6U6F1_LC_14_14_6  (
            .in0(N__11064),
            .in1(N__10252),
            .in2(N__10217),
            .in3(N__10186),
            .lcout(CLLBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m9_LC_14_17_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m9_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m9_LC_14_17_1 .LUT_INIT=16'b1101111000010010;
    LogicCell40 \U712_CHIP_RAM.m9_LC_14_17_1  (
            .in0(N__10096),
            .in1(N__10037),
            .in2(N__10000),
            .in3(N__9937),
            .lcout(LLBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m13_LC_14_17_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m13_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m13_LC_14_17_6 .LUT_INIT=16'b0000111011100000;
    LogicCell40 \U712_CHIP_RAM.m13_LC_14_17_6  (
            .in0(N__10036),
            .in1(N__10168),
            .in2(N__10001),
            .in3(N__10095),
            .lcout(UUBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m12_LC_14_17_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m12_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m12_LC_14_17_7 .LUT_INIT=16'b0111101101001000;
    LogicCell40 \U712_CHIP_RAM.m12_LC_14_17_7  (
            .in0(N__10094),
            .in1(N__10035),
            .in2(N__9999),
            .in3(N__9936),
            .lcout(UMBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WEn_LC_15_2_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_15_2_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_15_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_15_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9896),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11425),
            .ce(),
            .sr(N__11307));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_4_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_4_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_4_7  (
            .in0(N__9742),
            .in1(N__9794),
            .in2(_gnd_net_),
            .in3(N__11781),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11603),
            .ce(N__11573),
            .sr(N__11302));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_15_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_15_5_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_15_5_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_15_5_0  (
            .in0(N__9740),
            .in1(N__9792),
            .in2(_gnd_net_),
            .in3(N__11777),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .ce(N__11571),
            .sr(N__11299));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_5_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_5_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_5_7  (
            .in0(N__11778),
            .in1(N__10646),
            .in2(_gnd_net_),
            .in3(N__9741),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .ce(N__11571),
            .sr(N__11299));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_6_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_6_6  (
            .in0(N__11776),
            .in1(N__10642),
            .in2(_gnd_net_),
            .in3(N__11894),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__11569),
            .sr(N__11295));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_7_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_7_6  (
            .in0(N__11701),
            .in1(N__10418),
            .in2(_gnd_net_),
            .in3(N__10528),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11599),
            .ce(N__11567),
            .sr(N__11293));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_8_5  (
            .in0(N__10579),
            .in1(N__10527),
            .in2(_gnd_net_),
            .in3(N__11749),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__11566),
            .sr(N__11289));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_15_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_15_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_15_9_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_15_9_3  (
            .in0(N__10413),
            .in1(N__10517),
            .in2(_gnd_net_),
            .in3(N__11748),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__11563),
            .sr(N__11285));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_10_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_10_0  (
            .in0(N__11747),
            .in1(N__10450),
            .in2(_gnd_net_),
            .in3(N__10417),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11596),
            .ce(N__11561),
            .sr(N__11280));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_15_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_15_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_15_11_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_15_11_2  (
            .in0(N__10451),
            .in1(_gnd_net_),
            .in2(N__11710),
            .in3(N__10409),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__11559),
            .sr(N__11277));
    defparam \U712_CHIP_RAM.DMA_CYCLE_RNIVA8H_LC_15_14_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_RNIVA8H_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_RNIVA8H_LC_15_14_4 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_RNIVA8H_LC_15_14_4  (
            .in0(N__10351),
            .in1(N__10712),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_345 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_15_17_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_15_17_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_15_17_4 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_15_17_4  (
            .in0(N__10708),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10852),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11467),
            .ce(),
            .sr(N__11250));
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_RNIVHJN_LC_15_19_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_RNIVHJN_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_RNIVHJN_LC_15_19_0 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \U712_CHIP_RAM.DMA_WRITE_CYCLE_RNIVHJN_LC_15_19_0  (
            .in0(N__10735),
            .in1(N__10707),
            .in2(_gnd_net_),
            .in3(N__10845),
            .lcout(DMA_LATCH_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CASn_LC_16_4_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_16_4_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_16_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_16_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12247),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11430),
            .ce(),
            .sr(N__11306));
    defparam \U712_CHIP_RAM.CRCSn_LC_16_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_16_4_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_16_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_16_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12013),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11430),
            .ce(),
            .sr(N__11306));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_16_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_16_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_16_6_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_16_6_0  (
            .in0(N__11938),
            .in1(N__11893),
            .in2(_gnd_net_),
            .in3(N__11775),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11600),
            .ce(N__11572),
            .sr(N__11300));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_16_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_16_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_16_7_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_16_7_1  (
            .in0(N__11841),
            .in1(N__11521),
            .in2(_gnd_net_),
            .in3(N__11700),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11598),
            .ce(N__11570),
            .sr(N__11296));
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_16_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_16_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_16_9_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_0_LC_16_9_0  (
            .in0(_gnd_net_),
            .in1(N__11522),
            .in2(_gnd_net_),
            .in3(N__11498),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11445),
            .ce(),
            .sr(N__11290));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIQ44J_LC_24_19_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIQ44J_LC_24_19_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIQ44J_LC_24_19_1 .LUT_INIT=16'b0101010101000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNIQ44J_LC_24_19_1  (
            .in0(N__11129),
            .in1(N__10683),
            .in2(N__10836),
            .in3(N__11087),
            .lcout(N_338_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_RNIRVG61_LC_24_19_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_RNIRVG61_LC_24_19_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_RNIRVG61_LC_24_19_5 .LUT_INIT=16'b0010011100001111;
    LogicCell40 \U712_CHIP_RAM.DMA_WRITE_CYCLE_RNIRVG61_LC_24_19_5  (
            .in0(N__10830),
            .in1(N__10802),
            .in2(N__10742),
            .in3(N__10684),
            .lcout(N_328_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U712_TOP

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 19 2024 10:10:35

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U111_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U111_TOP
entity U111_TOP is
port (
    D_LL_AMIGA : inout std_logic_vector(7 downto 0);
    D_LM_AMIGA : inout std_logic_vector(7 downto 0);
    D_UU_AMIGA : inout std_logic_vector(7 downto 0);
    D_UM_AMIGA : inout std_logic_vector(7 downto 0);
    D_UU_040 : inout std_logic_vector(7 downto 0);
    D_LL_040 : inout std_logic_vector(7 downto 0);
    D_LM_040 : inout std_logic_vector(7 downto 0);
    D_UM_040 : inout std_logic_vector(7 downto 0);
    A_AMIGA : out std_logic_vector(1 downto 0);
    A_040 : in std_logic_vector(1 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    TSn : out std_logic;
    RESETn : in std_logic;
    CLKRAMA : out std_logic;
    PORTSIZE : in std_logic;
    CLK40B : out std_logic;
    TBI_CPUn : out std_logic;
    TAn : out std_logic;
    CPUBGn : out std_logic;
    BUFENn : out std_logic;
    RnW : in std_logic;
    CLK80_CPU : out std_logic;
    BUFDIR : out std_logic;
    TCI_CPUn : out std_logic;
    TS_CPUn : in std_logic;
    CLKRAMB : out std_logic;
    CLK40A : out std_logic;
    DMAn : out std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    TACKn : in std_logic;
    BGn : in std_logic);
end U111_TOP;

-- Architecture of U111_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U111_TOP is

signal \N__8230\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7827\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7275\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6996\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3997\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3959\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3938\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3779\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3622\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3587\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3548\ : std_logic;
signal \N__3545\ : std_logic;
signal \N__3542\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3521\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3482\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3476\ : std_logic;
signal \N__3473\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3382\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3353\ : std_logic;
signal \N__3350\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3338\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3329\ : std_logic;
signal \N__3326\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3263\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3254\ : std_logic;
signal \N__3251\ : std_logic;
signal \N__3248\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3176\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3157\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3121\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3067\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2987\ : std_logic;
signal \N__2984\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2932\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2920\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2870\ : std_logic;
signal \N__2867\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2854\ : std_logic;
signal \N__2851\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2845\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2836\ : std_logic;
signal \N__2833\ : std_logic;
signal \N__2830\ : std_logic;
signal \N__2827\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2767\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2752\ : std_logic;
signal \N__2749\ : std_logic;
signal \N__2746\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2737\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2705\ : std_logic;
signal \N__2702\ : std_logic;
signal \N__2699\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2689\ : std_logic;
signal \N__2686\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2669\ : std_logic;
signal \N__2668\ : std_logic;
signal \N__2661\ : std_logic;
signal \N__2658\ : std_logic;
signal \N__2655\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2647\ : std_logic;
signal \N__2646\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2644\ : std_logic;
signal \N__2643\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2639\ : std_logic;
signal \N__2636\ : std_logic;
signal \N__2635\ : std_logic;
signal \N__2634\ : std_logic;
signal \N__2633\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2631\ : std_logic;
signal \N__2630\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2617\ : std_logic;
signal \N__2614\ : std_logic;
signal \N__2609\ : std_logic;
signal \N__2606\ : std_logic;
signal \N__2603\ : std_logic;
signal \N__2600\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2596\ : std_logic;
signal \N__2595\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2593\ : std_logic;
signal \N__2590\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2574\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2569\ : std_logic;
signal \N__2568\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2556\ : std_logic;
signal \N__2553\ : std_logic;
signal \N__2550\ : std_logic;
signal \N__2547\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2535\ : std_logic;
signal \N__2532\ : std_logic;
signal \N__2529\ : std_logic;
signal \N__2526\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2515\ : std_logic;
signal \N__2508\ : std_logic;
signal \N__2497\ : std_logic;
signal \N__2494\ : std_logic;
signal \N__2491\ : std_logic;
signal \N__2490\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2484\ : std_logic;
signal \N__2481\ : std_logic;
signal \N__2478\ : std_logic;
signal \N__2473\ : std_logic;
signal \N__2468\ : std_logic;
signal \N__2465\ : std_logic;
signal \N__2462\ : std_logic;
signal \N__2459\ : std_logic;
signal \N__2456\ : std_logic;
signal \N__2453\ : std_logic;
signal \N__2450\ : std_logic;
signal \N__2447\ : std_logic;
signal \N__2442\ : std_logic;
signal \N__2439\ : std_logic;
signal \N__2434\ : std_logic;
signal \N__2429\ : std_logic;
signal \N__2426\ : std_logic;
signal \N__2417\ : std_logic;
signal \N__2414\ : std_logic;
signal \N__2411\ : std_logic;
signal \N__2408\ : std_logic;
signal \N__2405\ : std_logic;
signal \N__2402\ : std_logic;
signal \N__2399\ : std_logic;
signal \N__2396\ : std_logic;
signal \N__2393\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2384\ : std_logic;
signal \N__2381\ : std_logic;
signal \N__2378\ : std_logic;
signal \N__2375\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2369\ : std_logic;
signal \N__2366\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2360\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2354\ : std_logic;
signal \N__2351\ : std_logic;
signal \N__2348\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2342\ : std_logic;
signal \N__2339\ : std_logic;
signal \N__2336\ : std_logic;
signal \N__2333\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2324\ : std_logic;
signal \N__2321\ : std_logic;
signal \N__2318\ : std_logic;
signal \N__2315\ : std_logic;
signal \N__2312\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2306\ : std_logic;
signal \N__2303\ : std_logic;
signal \N__2300\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2294\ : std_logic;
signal \N__2291\ : std_logic;
signal \N__2288\ : std_logic;
signal \N__2285\ : std_logic;
signal \N__2282\ : std_logic;
signal \N__2279\ : std_logic;
signal \N__2276\ : std_logic;
signal \N__2275\ : std_logic;
signal \N__2272\ : std_logic;
signal \N__2269\ : std_logic;
signal \N__2266\ : std_logic;
signal \N__2263\ : std_logic;
signal \N__2260\ : std_logic;
signal \N__2257\ : std_logic;
signal \N__2254\ : std_logic;
signal \N__2251\ : std_logic;
signal \N__2248\ : std_logic;
signal \N__2245\ : std_logic;
signal \N__2242\ : std_logic;
signal \N__2239\ : std_logic;
signal \N__2236\ : std_logic;
signal \N__2233\ : std_logic;
signal \N__2228\ : std_logic;
signal \N__2225\ : std_logic;
signal \N__2222\ : std_logic;
signal \N__2219\ : std_logic;
signal \N__2216\ : std_logic;
signal \N__2213\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \A_040_c_0\ : std_logic;
signal \A_AMIGA_c_0\ : std_logic;
signal \A_040_c_1\ : std_logic;
signal \A_AMIGA_c_1_cascade_\ : std_logic;
signal \D_LL_AMIGA_in_3\ : std_logic;
signal \un1_D_LL_AMIGA_3\ : std_logic;
signal \D_LL_AMIGA_in_4\ : std_logic;
signal \un1_D_LL_AMIGA_4\ : std_logic;
signal \D_UM_040_in_0\ : std_logic;
signal \D_LL_040_in_0\ : std_logic;
signal \un1_D_UM_040_0\ : std_logic;
signal \D_UM_040_in_2\ : std_logic;
signal \D_LL_040_in_2\ : std_logic;
signal \un1_D_UM_040_2\ : std_logic;
signal \D_LL_040_in_1\ : std_logic;
signal \D_UM_040_in_1\ : std_logic;
signal \un1_D_UM_040_1\ : std_logic;
signal \D_LL_040_in_7\ : std_logic;
signal \D_UM_040_in_7\ : std_logic;
signal \un1_D_UM_040_7\ : std_logic;
signal \D_UU_040_in_1\ : std_logic;
signal \D_LM_040_in_1\ : std_logic;
signal \un1_D_UU_040_1\ : std_logic;
signal \D_LM_AMIGA_in_3\ : std_logic;
signal \un1_D_LM_AMIGA_3\ : std_logic;
signal \D_LM_040_in_7\ : std_logic;
signal \D_UU_040_in_7\ : std_logic;
signal \un1_D_UU_040_7\ : std_logic;
signal \D_LM_040_in_3\ : std_logic;
signal \D_UU_040_in_3\ : std_logic;
signal \un1_D_UU_040_3\ : std_logic;
signal \RnW_c_i_0\ : std_logic;
signal \D_LL_AMIGA_in_6\ : std_logic;
signal \un1_D_LL_AMIGA_6\ : std_logic;
signal \D_LM_AMIGA_in_5\ : std_logic;
signal \un1_D_LM_AMIGA_5\ : std_logic;
signal \D_LM_AMIGA_in_7\ : std_logic;
signal \un1_D_LM_AMIGA_7\ : std_logic;
signal \TSn_c\ : std_logic;
signal \INVU111_CYCLE_SM.TSnC_net\ : std_logic;
signal \D_LL_AMIGA_in_0\ : std_logic;
signal \un1_D_LL_AMIGA_0\ : std_logic;
signal \D_UU_040_in_4\ : std_logic;
signal \D_LM_040_in_4\ : std_logic;
signal \un1_D_UU_040_4\ : std_logic;
signal \D_LL_AMIGA_in_1\ : std_logic;
signal \un1_D_LL_AMIGA_1\ : std_logic;
signal \D_LL_AMIGA_in_2\ : std_logic;
signal \un1_D_LL_AMIGA_2\ : std_logic;
signal \D_LM_AMIGA_in_0\ : std_logic;
signal \un1_D_LM_AMIGA_0\ : std_logic;
signal \D_UU_040_in_2\ : std_logic;
signal \D_LM_040_in_2\ : std_logic;
signal \un1_D_UU_040_2\ : std_logic;
signal \D_UU_040_in_0\ : std_logic;
signal \D_LM_040_in_0\ : std_logic;
signal \un1_D_UU_040_0\ : std_logic;
signal \D_LL_040_in_4\ : std_logic;
signal \D_UM_040_in_4\ : std_logic;
signal \un1_D_UM_040_4\ : std_logic;
signal \D_LM_AMIGA_in_2\ : std_logic;
signal \un1_D_LM_AMIGA_2\ : std_logic;
signal \D_LM_AMIGA_in_6\ : std_logic;
signal \un1_D_LM_AMIGA_6\ : std_logic;
signal \D_UM_040_in_3\ : std_logic;
signal \D_LL_040_in_3\ : std_logic;
signal \un1_D_UM_040_3\ : std_logic;
signal \D_UU_040_in_5\ : std_logic;
signal \D_LM_040_in_5\ : std_logic;
signal \un1_D_UU_040_5\ : std_logic;
signal \D_UM_040_in_5\ : std_logic;
signal \D_LL_040_in_5\ : std_logic;
signal \un1_D_UM_040_5\ : std_logic;
signal \D_LL_AMIGA_in_5\ : std_logic;
signal \un1_D_LL_AMIGA_5\ : std_logic;
signal \D_LL_AMIGA_in_7\ : std_logic;
signal \un1_D_LL_AMIGA_7\ : std_logic;
signal \un1_D_UM_AMIGA_2\ : std_logic;
signal \INVU111_CYCLE_SM.TA_ENC_net\ : std_logic;
signal \U111_CYCLE_SM.RESETn_c_i\ : std_logic;
signal \D_UM_AMIGA_in_2\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\ : std_logic;
signal \INVU111_CYCLE_SM.UM_LATCHED_nesr_2C_net\ : std_logic;
signal \U111_CYCLE_SM.un3_LW_CYCLE_START_cascade_\ : std_logic;
signal \TS_CPUn_c\ : std_logic;
signal \U111_CYCLE_SM.N_69_0_cascade_\ : std_logic;
signal \U111_CYCLE_SM.TS_EN_5\ : std_logic;
signal \U111_CYCLE_SM.TS_ENZ0\ : std_logic;
signal \INVU111_CYCLE_SM.LW_CYCLE_STARTC_net\ : std_logic;
signal \INVU111_CYCLE_SM.UU_LATCHED_nesr_6C_net\ : std_logic;
signal \PORTSIZE_c\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\ : std_logic;
signal \D_UU_AMIGA_in_3\ : std_logic;
signal \un1_D_UU_AMIGA_3\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\ : std_logic;
signal \D_UU_AMIGA_in_6\ : std_logic;
signal \un1_D_UU_AMIGA_6\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\ : std_logic;
signal \D_UU_AMIGA_in_2\ : std_logic;
signal \un1_D_UU_AMIGA_2\ : std_logic;
signal \GB_BUFFER_CLK40_THRU_CO\ : std_logic;
signal \D_LM_AMIGA_in_1\ : std_logic;
signal \un1_D_LM_AMIGA_1\ : std_logic;
signal \D_UM_040_in_6\ : std_logic;
signal \D_LL_040_in_6\ : std_logic;
signal \un1_D_UM_040_6\ : std_logic;
signal \U111_CYCLE_SM.TA_ENZ0\ : std_logic;
signal \U111_CYCLE_SM_TAn_0_i\ : std_logic;
signal \D_LM_AMIGA_in_4\ : std_logic;
signal \un1_D_LM_AMIGA_4\ : std_logic;
signal \INVU111_CYCLE_SM.LW_CYCLEC_net\ : std_logic;
signal \U111_CYCLE_SM.LW_CYCLE_0\ : std_logic;
signal \U111_CYCLE_SM.A_OUT_0_sqmuxa_0_a3_0\ : std_logic;
signal \CLK40\ : std_logic;
signal \U111_CYCLE_SM.N_91_cascade_\ : std_logic;
signal \U111_CYCLE_SM.LW_CYCLE_STARTZ0\ : std_logic;
signal \U111_CYCLE_SM.A_OUT_0_cascade_\ : std_logic;
signal \U111_CYCLE_SM.A_OUTZ0\ : std_logic;
signal \INVU111_CYCLE_SM.CYCLE_STATE_0C_net\ : std_logic;
signal \TACKn_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0_cascade_\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa\ : std_logic;
signal \INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\ : std_logic;
signal \D_UU_AMIGA_in_0\ : std_logic;
signal \un1_D_UU_AMIGA_0\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\ : std_logic;
signal \D_UM_AMIGA_in_5\ : std_logic;
signal \un1_D_UM_AMIGA_5\ : std_logic;
signal \U111_CYCLE_SM.un1_LW_TRANS_1_0\ : std_logic;
signal \D_UU_040_in_6\ : std_logic;
signal \D_LM_040_in_6\ : std_logic;
signal \A_AMIGA_c_1\ : std_logic;
signal \un1_D_UU_040_6\ : std_logic;
signal \D_UU_AMIGA_in_4\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\ : std_logic;
signal \un1_D_UU_AMIGA_4\ : std_logic;
signal \CLK80\ : std_logic;
signal \GB_BUFFER_CLK80_THRU_CO\ : std_logic;
signal \un1_D_UM_AMIGA_0\ : std_logic;
signal \un1_D_UM_AMIGA_6\ : std_logic;
signal \D_UM_AMIGA_in_6\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\ : std_logic;
signal \D_UM_AMIGA_in_0\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\ : std_logic;
signal \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net\ : std_logic;
signal \INVU111_CYCLE_SM.UM_LATCHED_nesr_1C_net\ : std_logic;
signal \INVU111_CYCLE_SM.UU_LATCHED_nesr_5C_net\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\ : std_logic;
signal \D_UM_AMIGA_in_3\ : std_logic;
signal \un1_D_UM_AMIGA_3\ : std_logic;
signal \D_UM_AMIGA_in_1\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\ : std_logic;
signal \un1_D_UM_AMIGA_1\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\ : std_logic;
signal \D_UU_AMIGA_in_1\ : std_logic;
signal \un1_D_UU_AMIGA_1\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\ : std_logic;
signal \D_UM_AMIGA_in_4\ : std_logic;
signal \un1_D_UM_AMIGA_4\ : std_logic;
signal \D_UM_AMIGA_in_7\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\ : std_logic;
signal \un1_D_UM_AMIGA_7\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\ : std_logic;
signal \D_UU_AMIGA_in_7\ : std_logic;
signal \un1_D_UU_AMIGA_7\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\ : std_logic;
signal \D_UU_AMIGA_in_5\ : std_logic;
signal \U111_CYCLE_SM.LW_CYCLEZ0\ : std_logic;
signal \un1_D_UU_AMIGA_5\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK40_IN_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \CPUBGn_wire\ : std_logic;
signal \A_040_wire\ : std_logic_vector(1 downto 0);
signal \A_AMIGA_wire\ : std_logic_vector(1 downto 0);
signal \CLK40B_wire\ : std_logic;
signal \TBI_CPUn_wire\ : std_logic;
signal \CLK40A_wire\ : std_logic;
signal \BUFDIR_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \TS_CPUn_wire\ : std_logic;
signal \CLKRAMA_wire\ : std_logic;
signal \TCI_CPUn_wire\ : std_logic;
signal \CLKRAMB_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \TAn_wire\ : std_logic;
signal \DMAn_wire\ : std_logic;
signal \CLK80_CPU_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \pll_pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK40_IN_wire\ <= CLK40_IN;
    \TACKn_wire\ <= TACKn;
    CPUBGn <= \CPUBGn_wire\;
    \A_040_wire\ <= A_040;
    A_AMIGA <= \A_AMIGA_wire\;
    CLK40B <= \CLK40B_wire\;
    TBI_CPUn <= \TBI_CPUn_wire\;
    CLK40A <= \CLK40A_wire\;
    BUFDIR <= \BUFDIR_wire\;
    \SIZ_wire\ <= SIZ;
    \TS_CPUn_wire\ <= TS_CPUn;
    CLKRAMA <= \CLKRAMA_wire\;
    TCI_CPUn <= \TCI_CPUn_wire\;
    CLKRAMB <= \CLKRAMB_wire\;
    BUFENn <= \BUFENn_wire\;
    \RnW_wire\ <= RnW;
    TAn <= \TAn_wire\;
    DMAn <= \DMAn_wire\;
    CLK80_CPU <= \CLK80_CPU_wire\;
    TSn <= \TSn_wire\;
    \PORTSIZE_wire\ <= PORTSIZE;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    \pll_pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll_pll\ : PLL40_2F
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            SCLK => '0',
            PLLOUTGLOBALA => \CLK80\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALB => \CLK40\,
            SDI => '0',
            PLLOUTCOREA => OPEN,
            BYPASS => '0',
            RESETB => \N__4458\,
            PLLOUTCOREB => OPEN,
            LOCK => OPEN,
            SDO => OPEN,
            EXTFEEDBACK => '0',
            DYNAMICDELAY => \pll_pll_DYNAMICDELAY_wire\,
            PLLIN => \N__8230\
        );

    \pll_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \VCCG0\,
            DIN => '0',
            DOUT => \N__8230\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \D_UM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8214\,
            DIN => \N__8213\,
            DOUT => \N__8212\,
            PACKAGEPIN => D_UM_040(3)
        );

    \D_UM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8214\,
            PADOUT => \N__8213\,
            PADIN => \N__8212\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5114\,
            DIN0 => \D_UM_040_in_3\,
            DOUT0 => \N__7022\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8205\,
            DIN => \N__8204\,
            DOUT => \N__8203\,
            PACKAGEPIN => D_LL_AMIGA(1)
        );

    \D_LL_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8205\,
            PADOUT => \N__8204\,
            PADIN => \N__8203\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2682\,
            DIN0 => \D_LL_AMIGA_in_1\,
            DOUT0 => \N__3163\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8196\,
            DIN => \N__8195\,
            DOUT => \N__8194\,
            PACKAGEPIN => D_UU_AMIGA(5)
        );

    \D_UU_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8196\,
            PADOUT => \N__8195\,
            PADIN => \N__8194\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2630\,
            DIN0 => \D_UU_AMIGA_in_5\,
            DOUT0 => \N__3707\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8187\,
            DIN => \N__8186\,
            DOUT => \N__8185\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8187\,
            PADOUT => \N__8186\,
            PADIN => \N__8185\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TACKn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8178\,
            DIN => \N__8177\,
            DOUT => \N__8176\,
            PACKAGEPIN => D_UU_040(6)
        );

    \D_UU_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8178\,
            PADOUT => \N__8177\,
            PADIN => \N__8176\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5158\,
            DIN0 => \D_UU_040_in_6\,
            DOUT0 => \N__4904\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CPUBGn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8169\,
            DIN => \N__8168\,
            DOUT => \N__8167\,
            PACKAGEPIN => \CPUBGn_wire\
        );

    \CPUBGn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8169\,
            PADOUT => \N__8168\,
            PADIN => \N__8167\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8160\,
            DIN => \N__8159\,
            DOUT => \N__8158\,
            PACKAGEPIN => D_LL_040(7)
        );

    \D_LL_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8160\,
            PADOUT => \N__8159\,
            PADIN => \N__8158\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5220\,
            DIN0 => \D_LL_040_in_7\,
            DOUT0 => \N__4283\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8151\,
            DIN => \N__8150\,
            DOUT => \N__8149\,
            PACKAGEPIN => D_LL_AMIGA(4)
        );

    \D_LL_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8151\,
            PADOUT => \N__8150\,
            PADIN => \N__8149\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2681\,
            DIN0 => \D_LL_AMIGA_in_4\,
            DOUT0 => \N__4004\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8142\,
            DIN => \N__8141\,
            DOUT => \N__8140\,
            PACKAGEPIN => D_UM_AMIGA(3)
        );

    \D_UM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8142\,
            PADOUT => \N__8141\,
            PADIN => \N__8140\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2574\,
            DIN0 => \D_UM_AMIGA_in_3\,
            DOUT0 => \N__3788\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8133\,
            DIN => \N__8132\,
            DOUT => \N__8131\,
            PACKAGEPIN => D_UU_040(3)
        );

    \D_UU_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8133\,
            PADOUT => \N__8132\,
            PADIN => \N__8131\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5153\,
            DIN0 => \D_UU_040_in_3\,
            DOUT0 => \N__4361\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8124\,
            DIN => \N__8123\,
            DOUT => \N__8122\,
            PACKAGEPIN => \A_040_wire\(1)
        );

    \A_040_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8124\,
            PADOUT => \N__8123\,
            PADIN => \N__8122\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8115\,
            DIN => \N__8114\,
            DOUT => \N__8113\,
            PACKAGEPIN => D_LM_AMIGA(3)
        );

    \D_LM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8115\,
            PADOUT => \N__8114\,
            PADIN => \N__8113\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2647\,
            DIN0 => \D_LM_AMIGA_in_3\,
            DOUT0 => \N__2780\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8106\,
            DIN => \N__8105\,
            DOUT => \N__8104\,
            PACKAGEPIN => D_LM_040(0)
        );

    \D_LM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8106\,
            PADOUT => \N__8105\,
            PADIN => \N__8104\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5221\,
            DIN0 => \D_LM_040_in_0\,
            DOUT0 => \N__3260\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8097\,
            DIN => \N__8096\,
            DOUT => \N__8095\,
            PACKAGEPIN => D_UM_AMIGA(6)
        );

    \D_UM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8097\,
            PADOUT => \N__8096\,
            PADIN => \N__8095\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2629\,
            DIN0 => \D_UM_AMIGA_in_6\,
            DOUT0 => \N__4685\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8088\,
            DIN => \N__8087\,
            DOUT => \N__8086\,
            PACKAGEPIN => D_LM_AMIGA(4)
        );

    \D_LM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8088\,
            PADOUT => \N__8087\,
            PADIN => \N__8086\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2632\,
            DIN0 => \D_LM_AMIGA_in_4\,
            DOUT0 => \N__3419\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8079\,
            DIN => \N__8078\,
            DOUT => \N__8077\,
            PACKAGEPIN => \A_AMIGA_wire\(1)
        );

    \A_AMIGA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8079\,
            PADOUT => \N__8078\,
            PADIN => \N__8077\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5833\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8070\,
            DIN => \N__8069\,
            DOUT => \N__8068\,
            PACKAGEPIN => D_LM_040(7)
        );

    \D_LM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8070\,
            PADOUT => \N__8069\,
            PADIN => \N__8068\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5039\,
            DIN0 => \D_LM_040_in_7\,
            DOUT0 => \N__3500\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8061\,
            DIN => \N__8060\,
            DOUT => \N__8059\,
            PACKAGEPIN => D_UM_040(4)
        );

    \D_UM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8061\,
            PADOUT => \N__8060\,
            PADIN => \N__8059\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5154\,
            DIN0 => \D_UM_040_in_4\,
            DOUT0 => \N__6794\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8052\,
            DIN => \N__8051\,
            DOUT => \N__8050\,
            PACKAGEPIN => \CLK40B_wire\
        );

    \CLK40B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8052\,
            PADOUT => \N__8051\,
            PADIN => \N__8050\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4823\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8043\,
            DIN => \N__8042\,
            DOUT => \N__8041\,
            PACKAGEPIN => D_UU_AMIGA(0)
        );

    \D_UU_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8043\,
            PADOUT => \N__8042\,
            PADIN => \N__8041\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2644\,
            DIN0 => \D_UU_AMIGA_in_0\,
            DOUT0 => \N__4022\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8034\,
            DIN => \N__8033\,
            DOUT => \N__8032\,
            PACKAGEPIN => \A_040_wire\(0)
        );

    \A_040_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8034\,
            PADOUT => \N__8033\,
            PADIN => \N__8032\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8025\,
            DIN => \N__8024\,
            DOUT => \N__8023\,
            PACKAGEPIN => D_LM_AMIGA(0)
        );

    \D_LM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8025\,
            PADOUT => \N__8024\,
            PADIN => \N__8023\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2569\,
            DIN0 => \D_LM_AMIGA_in_0\,
            DOUT0 => \N__4070\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8016\,
            DIN => \N__8015\,
            DOUT => \N__8014\,
            PACKAGEPIN => D_UM_040(1)
        );

    \D_UM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8016\,
            PADOUT => \N__8015\,
            PADIN => \N__8014\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5112\,
            DIN0 => \D_UM_040_in_1\,
            DOUT0 => \N__6944\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8007\,
            DIN => \N__8006\,
            DOUT => \N__8005\,
            PACKAGEPIN => \TBI_CPUn_wire\
        );

    \TBI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8007\,
            PADOUT => \N__8006\,
            PADIN => \N__8005\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7998\,
            DIN => \N__7997\,
            DOUT => \N__7996\,
            PACKAGEPIN => \CLK40A_wire\
        );

    \CLK40A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7998\,
            PADOUT => \N__7997\,
            PADIN => \N__7996\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4822\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7989\,
            DIN => \N__7988\,
            DOUT => \N__7987\,
            PACKAGEPIN => D_LM_040(3)
        );

    \D_LM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7989\,
            PADOUT => \N__7988\,
            PADIN => \N__7987\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5145\,
            DIN0 => \D_LM_040_in_3\,
            DOUT0 => \N__2885\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7980\,
            DIN => \N__7979\,
            DOUT => \N__7978\,
            PACKAGEPIN => D_LL_040(4)
        );

    \D_LL_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7980\,
            PADOUT => \N__7979\,
            PADIN => \N__7978\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5238\,
            DIN0 => \D_LL_040_in_4\,
            DOUT0 => \N__2318\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7971\,
            DIN => \N__7970\,
            DOUT => \N__7969\,
            PACKAGEPIN => D_LL_AMIGA(7)
        );

    \D_LL_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7971\,
            PADOUT => \N__7970\,
            PADIN => \N__7969\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2568\,
            DIN0 => \D_LL_AMIGA_in_7\,
            DOUT0 => \N__3077\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7962\,
            DIN => \N__7961\,
            DOUT => \N__7960\,
            PACKAGEPIN => D_UU_AMIGA(7)
        );

    \D_UU_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7962\,
            PADOUT => \N__7961\,
            PADIN => \N__7960\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2642\,
            DIN0 => \D_UU_AMIGA_in_7\,
            DOUT0 => \N__2798\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7953\,
            DIN => \N__7952\,
            DOUT => \N__7951\,
            PACKAGEPIN => \BUFDIR_wire\
        );

    \BUFDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7953\,
            PADOUT => \N__7952\,
            PADIN => \N__7951\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5236\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7944\,
            DIN => \N__7943\,
            DOUT => \N__7942\,
            PACKAGEPIN => D_LM_AMIGA(5)
        );

    \D_LM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7944\,
            PADOUT => \N__7943\,
            PADIN => \N__7942\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2595\,
            DIN0 => \D_LM_AMIGA_in_5\,
            DOUT0 => \N__3743\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7935\,
            DIN => \N__7934\,
            DOUT => \N__7933\,
            PACKAGEPIN => D_UU_040(4)
        );

    \D_UU_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7935\,
            PADOUT => \N__7934\,
            PADIN => \N__7933\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5189\,
            DIN0 => \D_UU_040_in_4\,
            DOUT0 => \N__5660\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7926\,
            DIN => \N__7925\,
            DOUT => \N__7924\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7926\,
            PADOUT => \N__7925\,
            PADIN => \N__7924\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7917\,
            DIN => \N__7916\,
            DOUT => \N__7915\,
            PACKAGEPIN => D_LM_040(6)
        );

    \D_LM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7917\,
            PADOUT => \N__7916\,
            PADIN => \N__7915\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5022\,
            DIN0 => \D_LM_040_in_6\,
            DOUT0 => \N__3872\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7908\,
            DIN => \N__7907\,
            DOUT => \N__7906\,
            PACKAGEPIN => D_UM_040(5)
        );

    \D_UM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7908\,
            PADOUT => \N__7907\,
            PADIN => \N__7906\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5155\,
            DIN0 => \D_UM_040_in_5\,
            DOUT0 => \N__6347\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TS_CPUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7899\,
            DIN => \N__7898\,
            DOUT => \N__7897\,
            PACKAGEPIN => \TS_CPUn_wire\
        );

    \TS_CPUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7899\,
            PADOUT => \N__7898\,
            PADIN => \N__7897\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TS_CPUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7890\,
            DIN => \N__7889\,
            DOUT => \N__7888\,
            PACKAGEPIN => D_LL_040(1)
        );

    \D_LL_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7890\,
            PADOUT => \N__7889\,
            PADIN => \N__7888\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5237\,
            DIN0 => \D_LL_040_in_1\,
            DOUT0 => \N__3341\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7881\,
            DIN => \N__7880\,
            DOUT => \N__7879\,
            PACKAGEPIN => D_LL_AMIGA(3)
        );

    \D_LL_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7881\,
            PADOUT => \N__7880\,
            PADIN => \N__7879\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2689\,
            DIN0 => \D_LL_AMIGA_in_3\,
            DOUT0 => \N__3830\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7872\,
            DIN => \N__7871\,
            DOUT => \N__7870\,
            PACKAGEPIN => D_UM_AMIGA(5)
        );

    \D_UM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7872\,
            PADOUT => \N__7871\,
            PADIN => \N__7870\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2645\,
            DIN0 => \D_UM_AMIGA_in_5\,
            DOUT0 => \N__3614\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7863\,
            DIN => \N__7862\,
            DOUT => \N__7861\,
            PACKAGEPIN => D_UU_040(1)
        );

    \D_UU_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7863\,
            PADOUT => \N__7862\,
            PADIN => \N__7861\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5115\,
            DIN0 => \D_UU_040_in_1\,
            DOUT0 => \N__6872\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7854\,
            DIN => \N__7853\,
            DOUT => \N__7852\,
            PACKAGEPIN => D_UU_AMIGA(3)
        );

    \D_UU_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7854\,
            PADOUT => \N__7853\,
            PADIN => \N__7852\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2631\,
            DIN0 => \D_UU_AMIGA_in_3\,
            DOUT0 => \N__2708\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7845\,
            DIN => \N__7844\,
            DOUT => \N__7843\,
            PACKAGEPIN => D_LM_AMIGA(1)
        );

    \D_LM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7845\,
            PADOUT => \N__7844\,
            PADIN => \N__7843\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2515\,
            DIN0 => \D_LM_AMIGA_in_1\,
            DOUT0 => \N__2956\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7836\,
            DIN => \N__7835\,
            DOUT => \N__7834\,
            PACKAGEPIN => D_LM_040(2)
        );

    \D_LM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7836\,
            PADOUT => \N__7835\,
            PADIN => \N__7834\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5194\,
            DIN0 => \D_LM_040_in_2\,
            DOUT0 => \N__3905\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7827\,
            DIN => \N__7826\,
            DOUT => \N__7825\,
            PACKAGEPIN => D_LL_040(5)
        );

    \D_LL_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7827\,
            PADOUT => \N__7826\,
            PADIN => \N__7825\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5222\,
            DIN0 => \D_LL_040_in_5\,
            DOUT0 => \N__4319\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7818\,
            DIN => \N__7817\,
            DOUT => \N__7816\,
            PACKAGEPIN => D_LL_AMIGA(6)
        );

    \D_LL_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7818\,
            PADOUT => \N__7817\,
            PADIN => \N__7816\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2668\,
            DIN0 => \D_LL_AMIGA_in_6\,
            DOUT0 => \N__4736\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7809\,
            DIN => \N__7808\,
            DOUT => \N__7807\,
            PACKAGEPIN => D_UU_AMIGA(6)
        );

    \D_UU_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7809\,
            PADOUT => \N__7808\,
            PADIN => \N__7807\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2646\,
            DIN0 => \D_UU_AMIGA_in_6\,
            DOUT0 => \N__5723\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7800\,
            DIN => \N__7799\,
            DOUT => \N__7798\,
            PACKAGEPIN => D_UM_AMIGA(1)
        );

    \D_UM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7800\,
            PADOUT => \N__7799\,
            PADIN => \N__7798\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2596\,
            DIN0 => \D_UM_AMIGA_in_1\,
            DOUT0 => \N__3092\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7791\,
            DIN => \N__7790\,
            DOUT => \N__7789\,
            PACKAGEPIN => D_UU_040(5)
        );

    \D_UU_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7791\,
            PADOUT => \N__7790\,
            PADIN => \N__7789\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5156\,
            DIN0 => \D_UU_040_in_5\,
            DOUT0 => \N__7214\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7782\,
            DIN => \N__7781\,
            DOUT => \N__7780\,
            PACKAGEPIN => \CLKRAMA_wire\
        );

    \CLKRAMA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7782\,
            PADOUT => \N__7781\,
            PADIN => \N__7780\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5597\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7773\,
            DIN => \N__7772\,
            DOUT => \N__7771\,
            PACKAGEPIN => D_UM_040(2)
        );

    \D_UM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7773\,
            PADOUT => \N__7772\,
            PADIN => \N__7771\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5060\,
            DIN0 => \D_UM_040_in_2\,
            DOUT0 => \N__4262\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7764\,
            DIN => \N__7763\,
            DOUT => \N__7762\,
            PACKAGEPIN => D_LL_040(2)
        );

    \D_LL_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7764\,
            PADOUT => \N__7763\,
            PADIN => \N__7762\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5224\,
            DIN0 => \D_LL_040_in_2\,
            DOUT0 => \N__3299\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7755\,
            DIN => \N__7754\,
            DOUT => \N__7753\,
            PACKAGEPIN => \TCI_CPUn_wire\
        );

    \TCI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7755\,
            PADOUT => \N__7754\,
            PADIN => \N__7753\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4466\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMB_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7746\,
            DIN => \N__7745\,
            DOUT => \N__7744\,
            PACKAGEPIN => \CLKRAMB_wire\
        );

    \CLKRAMB_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7746\,
            PADOUT => \N__7745\,
            PADIN => \N__7744\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5583\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7737\,
            DIN => \N__7736\,
            DOUT => \N__7735\,
            PACKAGEPIN => D_LL_AMIGA(2)
        );

    \D_LL_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7737\,
            PADOUT => \N__7736\,
            PADIN => \N__7735\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2690\,
            DIN0 => \D_LL_AMIGA_in_2\,
            DOUT0 => \N__3226\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7728\,
            DIN => \N__7727\,
            DOUT => \N__7726\,
            PACKAGEPIN => D_UM_AMIGA(4)
        );

    \D_UM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7728\,
            PADOUT => \N__7727\,
            PADIN => \N__7726\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2594\,
            DIN0 => \D_UM_AMIGA_in_4\,
            DOUT0 => \N__3938\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7719\,
            DIN => \N__7718\,
            DOUT => \N__7717\,
            PACKAGEPIN => D_UU_AMIGA(2)
        );

    \D_UU_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7719\,
            PADOUT => \N__7718\,
            PADIN => \N__7717\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2643\,
            DIN0 => \D_UU_AMIGA_in_2\,
            DOUT0 => \N__4106\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7710\,
            DIN => \N__7709\,
            DOUT => \N__7708\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7710\,
            PADOUT => \N__7709\,
            PADIN => \N__7708\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7701\,
            DIN => \N__7700\,
            DOUT => \N__7699\,
            PACKAGEPIN => D_LM_AMIGA(6)
        );

    \D_LM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7701\,
            PADOUT => \N__7700\,
            PADIN => \N__7699\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2490\,
            DIN0 => \D_LM_AMIGA_in_6\,
            DOUT0 => \N__6041\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7692\,
            DIN => \N__7691\,
            DOUT => \N__7690\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7692\,
            PADOUT => \N__7691\,
            PADIN => \N__7690\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7683\,
            DIN => \N__7682\,
            DOUT => \N__7681\,
            PACKAGEPIN => D_LM_040(5)
        );

    \D_LM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7683\,
            PADOUT => \N__7682\,
            PADIN => \N__7681\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5062\,
            DIN0 => \D_LM_040_in_5\,
            DOUT0 => \N__3539\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7674\,
            DIN => \N__7673\,
            DOUT => \N__7672\,
            PACKAGEPIN => D_UM_040(6)
        );

    \D_UM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7674\,
            PADOUT => \N__7673\,
            PADIN => \N__7672\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5023\,
            DIN0 => \D_UM_040_in_6\,
            DOUT0 => \N__6608\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TAn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7665\,
            DIN => \N__7664\,
            DOUT => \N__7663\,
            PACKAGEPIN => \TAn_wire\
        );

    \TAn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7665\,
            PADOUT => \N__7664\,
            PADIN => \N__7663\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4652\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMAn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7656\,
            DIN => \N__7655\,
            DOUT => \N__7654\,
            PACKAGEPIN => \DMAn_wire\
        );

    \DMAn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7656\,
            PADOUT => \N__7655\,
            PADIN => \N__7654\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4465\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7647\,
            DIN => \N__7646\,
            DOUT => \N__7645\,
            PACKAGEPIN => D_LL_040(6)
        );

    \D_LL_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7647\,
            PADOUT => \N__7646\,
            PADIN => \N__7645\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5223\,
            DIN0 => \D_LL_040_in_6\,
            DOUT0 => \N__3578\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7638\,
            DIN => \N__7637\,
            DOUT => \N__7636\,
            PACKAGEPIN => D_LL_AMIGA(5)
        );

    \D_LL_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7638\,
            PADOUT => \N__7637\,
            PADIN => \N__7636\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2669\,
            DIN0 => \D_LL_AMIGA_in_5\,
            DOUT0 => \N__3662\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7629\,
            DIN => \N__7628\,
            DOUT => \N__7627\,
            PACKAGEPIN => D_UM_AMIGA(0)
        );

    \D_UM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7629\,
            PADOUT => \N__7628\,
            PADIN => \N__7627\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2635\,
            DIN0 => \D_UM_AMIGA_in_0\,
            DOUT0 => \N__2228\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7620\,
            DIN => \N__7619\,
            DOUT => \N__7618\,
            PACKAGEPIN => D_UU_040(2)
        );

    \D_UU_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7620\,
            PADOUT => \N__7619\,
            PADIN => \N__7618\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5188\,
            DIN0 => \D_UU_040_in_2\,
            DOUT0 => \N__4838\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7611\,
            DIN => \N__7610\,
            DOUT => \N__7609\,
            PACKAGEPIN => D_LM_AMIGA(2)
        );

    \D_LM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7611\,
            PADOUT => \N__7610\,
            PADIN => \N__7609\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2634\,
            DIN0 => \D_LM_AMIGA_in_2\,
            DOUT0 => \N__4144\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK80_CPU_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7602\,
            DIN => \N__7601\,
            DOUT => \N__7600\,
            PACKAGEPIN => \CLK80_CPU_wire\
        );

    \CLK80_CPU_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7602\,
            PADOUT => \N__7601\,
            PADIN => \N__7600\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5593\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7593\,
            DIN => \N__7592\,
            DOUT => \N__7591\,
            PACKAGEPIN => D_LL_040(3)
        );

    \D_LL_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7593\,
            PADOUT => \N__7592\,
            PADIN => \N__7591\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5245\,
            DIN0 => \D_LL_040_in_3\,
            DOUT0 => \N__2357\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7584\,
            DIN => \N__7583\,
            DOUT => \N__7582\,
            PACKAGEPIN => D_LM_040(1)
        );

    \D_LM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7584\,
            PADOUT => \N__7583\,
            PADIN => \N__7582\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5193\,
            DIN0 => \D_LM_040_in_1\,
            DOUT0 => \N__4775\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7575\,
            DIN => \N__7574\,
            DOUT => \N__7573\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7575\,
            PADOUT => \N__7574\,
            PADIN => \N__7573\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3485\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7566\,
            DIN => \N__7565\,
            DOUT => \N__7564\,
            PACKAGEPIN => D_UM_AMIGA(7)
        );

    \D_UM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7566\,
            PADOUT => \N__7565\,
            PADIN => \N__7564\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2593\,
            DIN0 => \D_UM_AMIGA_in_7\,
            DOUT0 => \N__2999\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7557\,
            DIN => \N__7556\,
            DOUT => \N__7555\,
            PACKAGEPIN => D_LM_AMIGA(7)
        );

    \D_LM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7557\,
            PADOUT => \N__7556\,
            PADIN => \N__7555\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2489\,
            DIN0 => \D_LM_AMIGA_in_7\,
            DOUT0 => \N__2864\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7548\,
            DIN => \N__7547\,
            DOUT => \N__7546\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7548\,
            PADOUT => \N__7547\,
            PADIN => \N__7546\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \PORTSIZE_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7539\,
            DIN => \N__7538\,
            DOUT => \N__7537\,
            PACKAGEPIN => \A_AMIGA_wire\(0)
        );

    \A_AMIGA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7539\,
            PADOUT => \N__7538\,
            PADIN => \N__7537\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2402\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7530\,
            DIN => \N__7529\,
            DOUT => \N__7528\,
            PACKAGEPIN => D_LM_040(4)
        );

    \D_LM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7530\,
            PADOUT => \N__7529\,
            PADIN => \N__7528\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5105\,
            DIN0 => \D_LM_040_in_4\,
            DOUT0 => \N__4613\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7521\,
            DIN => \N__7520\,
            DOUT => \N__7519\,
            PACKAGEPIN => D_UM_040(7)
        );

    \D_UM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7521\,
            PADOUT => \N__7520\,
            PADIN => \N__7519\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5113\,
            DIN0 => \D_UM_040_in_7\,
            DOUT0 => \N__6713\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7512\,
            DIN => \N__7511\,
            DOUT => \N__7510\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7512\,
            PADOUT => \N__7511\,
            PADIN => \N__7510\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7503\,
            DIN => \N__7502\,
            DOUT => \N__7501\,
            PACKAGEPIN => D_UU_AMIGA(1)
        );

    \D_UU_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7503\,
            PADOUT => \N__7502\,
            PADIN => \N__7501\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2573\,
            DIN0 => \D_UU_AMIGA_in_1\,
            DOUT0 => \N__2909\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7494\,
            DIN => \N__7493\,
            DOUT => \N__7492\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7494\,
            PADOUT => \N__7493\,
            PADIN => \N__7492\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4821\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7485\,
            DIN => \N__7484\,
            DOUT => \N__7483\,
            PACKAGEPIN => D_UM_040(0)
        );

    \D_UM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7485\,
            PADOUT => \N__7484\,
            PADIN => \N__7483\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5061\,
            DIN0 => \D_UM_040_in_0\,
            DOUT0 => \N__6629\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7476\,
            DIN => \N__7475\,
            DOUT => \N__7474\,
            PACKAGEPIN => D_LL_AMIGA(0)
        );

    \D_LL_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7476\,
            PADOUT => \N__7475\,
            PADIN => \N__7474\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2567\,
            DIN0 => \D_LL_AMIGA_in_0\,
            DOUT0 => \N__2275\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7467\,
            DIN => \N__7466\,
            DOUT => \N__7465\,
            PACKAGEPIN => D_UU_AMIGA(4)
        );

    \D_UU_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7467\,
            PADOUT => \N__7466\,
            PADIN => \N__7465\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2525\,
            DIN0 => \D_UU_AMIGA_in_4\,
            DOUT0 => \N__3377\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7458\,
            DIN => \N__7457\,
            DOUT => \N__7456\,
            PACKAGEPIN => D_UU_040(7)
        );

    \D_UU_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7458\,
            PADOUT => \N__7457\,
            PADIN => \N__7456\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5157\,
            DIN0 => \D_UU_040_in_7\,
            DOUT0 => \N__6644\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7449\,
            DIN => \N__7448\,
            DOUT => \N__7447\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7449\,
            PADOUT => \N__7448\,
            PADIN => \N__7447\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7440\,
            DIN => \N__7439\,
            DOUT => \N__7438\,
            PACKAGEPIN => D_LL_040(0)
        );

    \D_LL_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7440\,
            PADOUT => \N__7439\,
            PADIN => \N__7438\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5246\,
            DIN0 => \D_LL_040_in_0\,
            DOUT0 => \N__3458\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7431\,
            DIN => \N__7430\,
            DOUT => \N__7429\,
            PACKAGEPIN => D_UM_AMIGA(2)
        );

    \D_UM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7431\,
            PADOUT => \N__7430\,
            PADIN => \N__7429\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2633\,
            DIN0 => \D_UM_AMIGA_in_2\,
            DOUT0 => \N__3179\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7422\,
            DIN => \N__7421\,
            DOUT => \N__7420\,
            PACKAGEPIN => D_UU_040(0)
        );

    \D_UU_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7422\,
            PADOUT => \N__7421\,
            PADIN => \N__7420\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5099\,
            DIN0 => \D_UU_040_in_0\,
            DOUT0 => \N__6416\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1925\ : InMux
    port map (
            O => \N__7403\,
            I => \N__7400\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__7400\,
            I => \N__7397\
        );

    \I__1923\ : Odrv12
    port map (
            O => \N__7397\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\
        );

    \I__1922\ : InMux
    port map (
            O => \N__7394\,
            I => \N__7390\
        );

    \I__1921\ : CascadeMux
    port map (
            O => \N__7393\,
            I => \N__7386\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__7390\,
            I => \N__7383\
        );

    \I__1919\ : InMux
    port map (
            O => \N__7389\,
            I => \N__7380\
        );

    \I__1918\ : InMux
    port map (
            O => \N__7386\,
            I => \N__7377\
        );

    \I__1917\ : Span4Mux_h
    port map (
            O => \N__7383\,
            I => \N__7374\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__7380\,
            I => \N__7371\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__7377\,
            I => \N__7368\
        );

    \I__1914\ : Span4Mux_v
    port map (
            O => \N__7374\,
            I => \N__7363\
        );

    \I__1913\ : Span4Mux_h
    port map (
            O => \N__7371\,
            I => \N__7363\
        );

    \I__1912\ : Span4Mux_v
    port map (
            O => \N__7368\,
            I => \N__7360\
        );

    \I__1911\ : Span4Mux_h
    port map (
            O => \N__7363\,
            I => \N__7355\
        );

    \I__1910\ : Span4Mux_v
    port map (
            O => \N__7360\,
            I => \N__7355\
        );

    \I__1909\ : Span4Mux_v
    port map (
            O => \N__7355\,
            I => \N__7352\
        );

    \I__1908\ : Sp12to4
    port map (
            O => \N__7352\,
            I => \N__7349\
        );

    \I__1907\ : Odrv12
    port map (
            O => \N__7349\,
            I => \D_UU_AMIGA_in_5\
        );

    \I__1906\ : InMux
    port map (
            O => \N__7346\,
            I => \N__7340\
        );

    \I__1905\ : InMux
    port map (
            O => \N__7345\,
            I => \N__7340\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__7340\,
            I => \N__7335\
        );

    \I__1903\ : InMux
    port map (
            O => \N__7339\,
            I => \N__7326\
        );

    \I__1902\ : InMux
    port map (
            O => \N__7338\,
            I => \N__7326\
        );

    \I__1901\ : Span4Mux_v
    port map (
            O => \N__7335\,
            I => \N__7318\
        );

    \I__1900\ : InMux
    port map (
            O => \N__7334\,
            I => \N__7308\
        );

    \I__1899\ : InMux
    port map (
            O => \N__7333\,
            I => \N__7308\
        );

    \I__1898\ : InMux
    port map (
            O => \N__7332\,
            I => \N__7308\
        );

    \I__1897\ : InMux
    port map (
            O => \N__7331\,
            I => \N__7305\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__7326\,
            I => \N__7301\
        );

    \I__1895\ : InMux
    port map (
            O => \N__7325\,
            I => \N__7296\
        );

    \I__1894\ : InMux
    port map (
            O => \N__7324\,
            I => \N__7296\
        );

    \I__1893\ : InMux
    port map (
            O => \N__7323\,
            I => \N__7293\
        );

    \I__1892\ : InMux
    port map (
            O => \N__7322\,
            I => \N__7288\
        );

    \I__1891\ : InMux
    port map (
            O => \N__7321\,
            I => \N__7288\
        );

    \I__1890\ : Sp12to4
    port map (
            O => \N__7318\,
            I => \N__7283\
        );

    \I__1889\ : InMux
    port map (
            O => \N__7317\,
            I => \N__7280\
        );

    \I__1888\ : InMux
    port map (
            O => \N__7316\,
            I => \N__7275\
        );

    \I__1887\ : InMux
    port map (
            O => \N__7315\,
            I => \N__7275\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__7308\,
            I => \N__7270\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__7305\,
            I => \N__7270\
        );

    \I__1884\ : InMux
    port map (
            O => \N__7304\,
            I => \N__7267\
        );

    \I__1883\ : Span4Mux_v
    port map (
            O => \N__7301\,
            I => \N__7258\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__7296\,
            I => \N__7258\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__7293\,
            I => \N__7258\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__7288\,
            I => \N__7258\
        );

    \I__1879\ : InMux
    port map (
            O => \N__7287\,
            I => \N__7253\
        );

    \I__1878\ : InMux
    port map (
            O => \N__7286\,
            I => \N__7253\
        );

    \I__1877\ : Span12Mux_h
    port map (
            O => \N__7283\,
            I => \N__7248\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__7280\,
            I => \N__7243\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__7275\,
            I => \N__7243\
        );

    \I__1874\ : Span4Mux_v
    port map (
            O => \N__7270\,
            I => \N__7238\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__7267\,
            I => \N__7238\
        );

    \I__1872\ : Span4Mux_v
    port map (
            O => \N__7258\,
            I => \N__7233\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__7253\,
            I => \N__7233\
        );

    \I__1870\ : InMux
    port map (
            O => \N__7252\,
            I => \N__7230\
        );

    \I__1869\ : InMux
    port map (
            O => \N__7251\,
            I => \N__7227\
        );

    \I__1868\ : Odrv12
    port map (
            O => \N__7248\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1867\ : Odrv12
    port map (
            O => \N__7243\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__7238\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1865\ : Odrv4
    port map (
            O => \N__7233\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__7230\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__7227\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1862\ : IoInMux
    port map (
            O => \N__7214\,
            I => \N__7211\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__7211\,
            I => \N__7208\
        );

    \I__1860\ : Span4Mux_s2_v
    port map (
            O => \N__7208\,
            I => \N__7205\
        );

    \I__1859\ : Span4Mux_v
    port map (
            O => \N__7205\,
            I => \N__7202\
        );

    \I__1858\ : Sp12to4
    port map (
            O => \N__7202\,
            I => \N__7199\
        );

    \I__1857\ : Span12Mux_s10_h
    port map (
            O => \N__7199\,
            I => \N__7196\
        );

    \I__1856\ : Odrv12
    port map (
            O => \N__7196\,
            I => \un1_D_UU_AMIGA_5\
        );

    \I__1855\ : CEMux
    port map (
            O => \N__7193\,
            I => \N__7185\
        );

    \I__1854\ : CEMux
    port map (
            O => \N__7192\,
            I => \N__7182\
        );

    \I__1853\ : CEMux
    port map (
            O => \N__7191\,
            I => \N__7179\
        );

    \I__1852\ : CEMux
    port map (
            O => \N__7190\,
            I => \N__7176\
        );

    \I__1851\ : CEMux
    port map (
            O => \N__7189\,
            I => \N__7173\
        );

    \I__1850\ : CEMux
    port map (
            O => \N__7188\,
            I => \N__7170\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__7185\,
            I => \N__7165\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__7182\,
            I => \N__7165\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__7179\,
            I => \N__7160\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__7176\,
            I => \N__7160\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__7173\,
            I => \N__7157\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__7170\,
            I => \N__7154\
        );

    \I__1843\ : Odrv4
    port map (
            O => \N__7165\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\
        );

    \I__1842\ : Odrv4
    port map (
            O => \N__7160\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\
        );

    \I__1841\ : Odrv4
    port map (
            O => \N__7157\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__7154\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\
        );

    \I__1839\ : SRMux
    port map (
            O => \N__7145\,
            I => \N__7140\
        );

    \I__1838\ : SRMux
    port map (
            O => \N__7144\,
            I => \N__7135\
        );

    \I__1837\ : SRMux
    port map (
            O => \N__7143\,
            I => \N__7132\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__7140\,
            I => \N__7129\
        );

    \I__1835\ : SRMux
    port map (
            O => \N__7139\,
            I => \N__7126\
        );

    \I__1834\ : SRMux
    port map (
            O => \N__7138\,
            I => \N__7122\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__7135\,
            I => \N__7119\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__7132\,
            I => \N__7116\
        );

    \I__1831\ : Span4Mux_h
    port map (
            O => \N__7129\,
            I => \N__7111\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__7126\,
            I => \N__7111\
        );

    \I__1829\ : SRMux
    port map (
            O => \N__7125\,
            I => \N__7108\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__7122\,
            I => \N__7105\
        );

    \I__1827\ : Span4Mux_h
    port map (
            O => \N__7119\,
            I => \N__7100\
        );

    \I__1826\ : Span4Mux_h
    port map (
            O => \N__7116\,
            I => \N__7100\
        );

    \I__1825\ : Span4Mux_h
    port map (
            O => \N__7111\,
            I => \N__7093\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__7108\,
            I => \N__7093\
        );

    \I__1823\ : Span4Mux_h
    port map (
            O => \N__7105\,
            I => \N__7093\
        );

    \I__1822\ : Odrv4
    port map (
            O => \N__7100\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0\
        );

    \I__1821\ : Odrv4
    port map (
            O => \N__7093\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0\
        );

    \I__1820\ : InMux
    port map (
            O => \N__7088\,
            I => \N__7085\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__7085\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\
        );

    \I__1818\ : InMux
    port map (
            O => \N__7082\,
            I => \N__7077\
        );

    \I__1817\ : InMux
    port map (
            O => \N__7081\,
            I => \N__7074\
        );

    \I__1816\ : InMux
    port map (
            O => \N__7080\,
            I => \N__7071\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__7077\,
            I => \N__7068\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__7074\,
            I => \N__7065\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__7071\,
            I => \N__7062\
        );

    \I__1812\ : Span4Mux_h
    port map (
            O => \N__7068\,
            I => \N__7059\
        );

    \I__1811\ : Span4Mux_v
    port map (
            O => \N__7065\,
            I => \N__7056\
        );

    \I__1810\ : Span4Mux_h
    port map (
            O => \N__7062\,
            I => \N__7053\
        );

    \I__1809\ : Sp12to4
    port map (
            O => \N__7059\,
            I => \N__7050\
        );

    \I__1808\ : Span4Mux_v
    port map (
            O => \N__7056\,
            I => \N__7047\
        );

    \I__1807\ : Span4Mux_v
    port map (
            O => \N__7053\,
            I => \N__7044\
        );

    \I__1806\ : Span12Mux_v
    port map (
            O => \N__7050\,
            I => \N__7041\
        );

    \I__1805\ : Sp12to4
    port map (
            O => \N__7047\,
            I => \N__7038\
        );

    \I__1804\ : Span4Mux_h
    port map (
            O => \N__7044\,
            I => \N__7035\
        );

    \I__1803\ : Span12Mux_v
    port map (
            O => \N__7041\,
            I => \N__7032\
        );

    \I__1802\ : Span12Mux_h
    port map (
            O => \N__7038\,
            I => \N__7027\
        );

    \I__1801\ : Sp12to4
    port map (
            O => \N__7035\,
            I => \N__7027\
        );

    \I__1800\ : Odrv12
    port map (
            O => \N__7032\,
            I => \D_UM_AMIGA_in_3\
        );

    \I__1799\ : Odrv12
    port map (
            O => \N__7027\,
            I => \D_UM_AMIGA_in_3\
        );

    \I__1798\ : IoInMux
    port map (
            O => \N__7022\,
            I => \N__7019\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__7019\,
            I => \N__7016\
        );

    \I__1796\ : Span4Mux_s3_h
    port map (
            O => \N__7016\,
            I => \N__7013\
        );

    \I__1795\ : Span4Mux_h
    port map (
            O => \N__7013\,
            I => \N__7010\
        );

    \I__1794\ : Span4Mux_h
    port map (
            O => \N__7010\,
            I => \N__7007\
        );

    \I__1793\ : Span4Mux_h
    port map (
            O => \N__7007\,
            I => \N__7004\
        );

    \I__1792\ : Span4Mux_v
    port map (
            O => \N__7004\,
            I => \N__7001\
        );

    \I__1791\ : Odrv4
    port map (
            O => \N__7001\,
            I => \un1_D_UM_AMIGA_3\
        );

    \I__1790\ : InMux
    port map (
            O => \N__6998\,
            I => \N__6993\
        );

    \I__1789\ : InMux
    port map (
            O => \N__6997\,
            I => \N__6990\
        );

    \I__1788\ : InMux
    port map (
            O => \N__6996\,
            I => \N__6987\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__6993\,
            I => \N__6984\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__6990\,
            I => \N__6981\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__6987\,
            I => \N__6978\
        );

    \I__1784\ : Sp12to4
    port map (
            O => \N__6984\,
            I => \N__6975\
        );

    \I__1783\ : Span4Mux_v
    port map (
            O => \N__6981\,
            I => \N__6970\
        );

    \I__1782\ : Span4Mux_v
    port map (
            O => \N__6978\,
            I => \N__6970\
        );

    \I__1781\ : Span12Mux_v
    port map (
            O => \N__6975\,
            I => \N__6967\
        );

    \I__1780\ : Sp12to4
    port map (
            O => \N__6970\,
            I => \N__6964\
        );

    \I__1779\ : Span12Mux_h
    port map (
            O => \N__6967\,
            I => \N__6961\
        );

    \I__1778\ : Span12Mux_h
    port map (
            O => \N__6964\,
            I => \N__6958\
        );

    \I__1777\ : Odrv12
    port map (
            O => \N__6961\,
            I => \D_UM_AMIGA_in_1\
        );

    \I__1776\ : Odrv12
    port map (
            O => \N__6958\,
            I => \D_UM_AMIGA_in_1\
        );

    \I__1775\ : InMux
    port map (
            O => \N__6953\,
            I => \N__6950\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__6950\,
            I => \N__6947\
        );

    \I__1773\ : Odrv4
    port map (
            O => \N__6947\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\
        );

    \I__1772\ : IoInMux
    port map (
            O => \N__6944\,
            I => \N__6941\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__6941\,
            I => \N__6938\
        );

    \I__1770\ : Span4Mux_s3_h
    port map (
            O => \N__6938\,
            I => \N__6935\
        );

    \I__1769\ : Sp12to4
    port map (
            O => \N__6935\,
            I => \N__6932\
        );

    \I__1768\ : Span12Mux_s10_v
    port map (
            O => \N__6932\,
            I => \N__6929\
        );

    \I__1767\ : Span12Mux_h
    port map (
            O => \N__6929\,
            I => \N__6926\
        );

    \I__1766\ : Odrv12
    port map (
            O => \N__6926\,
            I => \un1_D_UM_AMIGA_1\
        );

    \I__1765\ : InMux
    port map (
            O => \N__6923\,
            I => \N__6920\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__6920\,
            I => \N__6917\
        );

    \I__1763\ : Odrv4
    port map (
            O => \N__6917\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\
        );

    \I__1762\ : InMux
    port map (
            O => \N__6914\,
            I => \N__6911\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__6911\,
            I => \N__6906\
        );

    \I__1760\ : InMux
    port map (
            O => \N__6910\,
            I => \N__6903\
        );

    \I__1759\ : InMux
    port map (
            O => \N__6909\,
            I => \N__6900\
        );

    \I__1758\ : Span4Mux_v
    port map (
            O => \N__6906\,
            I => \N__6895\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__6903\,
            I => \N__6895\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__6900\,
            I => \N__6892\
        );

    \I__1755\ : Span4Mux_v
    port map (
            O => \N__6895\,
            I => \N__6889\
        );

    \I__1754\ : Span12Mux_v
    port map (
            O => \N__6892\,
            I => \N__6886\
        );

    \I__1753\ : Sp12to4
    port map (
            O => \N__6889\,
            I => \N__6883\
        );

    \I__1752\ : Span12Mux_h
    port map (
            O => \N__6886\,
            I => \N__6880\
        );

    \I__1751\ : Span12Mux_h
    port map (
            O => \N__6883\,
            I => \N__6877\
        );

    \I__1750\ : Odrv12
    port map (
            O => \N__6880\,
            I => \D_UU_AMIGA_in_1\
        );

    \I__1749\ : Odrv12
    port map (
            O => \N__6877\,
            I => \D_UU_AMIGA_in_1\
        );

    \I__1748\ : IoInMux
    port map (
            O => \N__6872\,
            I => \N__6869\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__6869\,
            I => \N__6866\
        );

    \I__1746\ : IoSpan4Mux
    port map (
            O => \N__6866\,
            I => \N__6863\
        );

    \I__1745\ : IoSpan4Mux
    port map (
            O => \N__6863\,
            I => \N__6860\
        );

    \I__1744\ : Span4Mux_s2_h
    port map (
            O => \N__6860\,
            I => \N__6857\
        );

    \I__1743\ : Sp12to4
    port map (
            O => \N__6857\,
            I => \N__6854\
        );

    \I__1742\ : Odrv12
    port map (
            O => \N__6854\,
            I => \un1_D_UU_AMIGA_1\
        );

    \I__1741\ : InMux
    port map (
            O => \N__6851\,
            I => \N__6848\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__6848\,
            I => \N__6845\
        );

    \I__1739\ : Odrv4
    port map (
            O => \N__6845\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\
        );

    \I__1738\ : InMux
    port map (
            O => \N__6842\,
            I => \N__6839\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__6839\,
            I => \N__6835\
        );

    \I__1736\ : InMux
    port map (
            O => \N__6838\,
            I => \N__6832\
        );

    \I__1735\ : Span4Mux_v
    port map (
            O => \N__6835\,
            I => \N__6828\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__6832\,
            I => \N__6825\
        );

    \I__1733\ : InMux
    port map (
            O => \N__6831\,
            I => \N__6822\
        );

    \I__1732\ : Span4Mux_v
    port map (
            O => \N__6828\,
            I => \N__6819\
        );

    \I__1731\ : Span4Mux_v
    port map (
            O => \N__6825\,
            I => \N__6814\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__6822\,
            I => \N__6814\
        );

    \I__1729\ : Sp12to4
    port map (
            O => \N__6819\,
            I => \N__6811\
        );

    \I__1728\ : Span4Mux_v
    port map (
            O => \N__6814\,
            I => \N__6808\
        );

    \I__1727\ : Span12Mux_s5_h
    port map (
            O => \N__6811\,
            I => \N__6805\
        );

    \I__1726\ : Sp12to4
    port map (
            O => \N__6808\,
            I => \N__6802\
        );

    \I__1725\ : Span12Mux_v
    port map (
            O => \N__6805\,
            I => \N__6797\
        );

    \I__1724\ : Span12Mux_h
    port map (
            O => \N__6802\,
            I => \N__6797\
        );

    \I__1723\ : Odrv12
    port map (
            O => \N__6797\,
            I => \D_UM_AMIGA_in_4\
        );

    \I__1722\ : IoInMux
    port map (
            O => \N__6794\,
            I => \N__6791\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__6791\,
            I => \N__6788\
        );

    \I__1720\ : IoSpan4Mux
    port map (
            O => \N__6788\,
            I => \N__6785\
        );

    \I__1719\ : IoSpan4Mux
    port map (
            O => \N__6785\,
            I => \N__6782\
        );

    \I__1718\ : Span4Mux_s3_v
    port map (
            O => \N__6782\,
            I => \N__6779\
        );

    \I__1717\ : Span4Mux_h
    port map (
            O => \N__6779\,
            I => \N__6776\
        );

    \I__1716\ : Span4Mux_v
    port map (
            O => \N__6776\,
            I => \N__6773\
        );

    \I__1715\ : Odrv4
    port map (
            O => \N__6773\,
            I => \un1_D_UM_AMIGA_4\
        );

    \I__1714\ : InMux
    port map (
            O => \N__6770\,
            I => \N__6766\
        );

    \I__1713\ : InMux
    port map (
            O => \N__6769\,
            I => \N__6763\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__6766\,
            I => \N__6759\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__6763\,
            I => \N__6756\
        );

    \I__1710\ : InMux
    port map (
            O => \N__6762\,
            I => \N__6753\
        );

    \I__1709\ : Span4Mux_h
    port map (
            O => \N__6759\,
            I => \N__6750\
        );

    \I__1708\ : Span4Mux_v
    port map (
            O => \N__6756\,
            I => \N__6745\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__6753\,
            I => \N__6745\
        );

    \I__1706\ : Span4Mux_v
    port map (
            O => \N__6750\,
            I => \N__6742\
        );

    \I__1705\ : Span4Mux_v
    port map (
            O => \N__6745\,
            I => \N__6739\
        );

    \I__1704\ : Sp12to4
    port map (
            O => \N__6742\,
            I => \N__6736\
        );

    \I__1703\ : Sp12to4
    port map (
            O => \N__6739\,
            I => \N__6733\
        );

    \I__1702\ : Span12Mux_v
    port map (
            O => \N__6736\,
            I => \N__6730\
        );

    \I__1701\ : Span12Mux_h
    port map (
            O => \N__6733\,
            I => \N__6727\
        );

    \I__1700\ : Odrv12
    port map (
            O => \N__6730\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__1699\ : Odrv12
    port map (
            O => \N__6727\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__1698\ : InMux
    port map (
            O => \N__6722\,
            I => \N__6719\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__6719\,
            I => \N__6716\
        );

    \I__1696\ : Odrv12
    port map (
            O => \N__6716\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\
        );

    \I__1695\ : IoInMux
    port map (
            O => \N__6713\,
            I => \N__6710\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__6710\,
            I => \N__6707\
        );

    \I__1693\ : IoSpan4Mux
    port map (
            O => \N__6707\,
            I => \N__6704\
        );

    \I__1692\ : Span4Mux_s1_h
    port map (
            O => \N__6704\,
            I => \N__6701\
        );

    \I__1691\ : Sp12to4
    port map (
            O => \N__6701\,
            I => \N__6698\
        );

    \I__1690\ : Span12Mux_h
    port map (
            O => \N__6698\,
            I => \N__6695\
        );

    \I__1689\ : Odrv12
    port map (
            O => \N__6695\,
            I => \un1_D_UM_AMIGA_7\
        );

    \I__1688\ : InMux
    port map (
            O => \N__6692\,
            I => \N__6689\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__6689\,
            I => \N__6686\
        );

    \I__1686\ : Odrv12
    port map (
            O => \N__6686\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\
        );

    \I__1685\ : InMux
    port map (
            O => \N__6683\,
            I => \N__6678\
        );

    \I__1684\ : InMux
    port map (
            O => \N__6682\,
            I => \N__6675\
        );

    \I__1683\ : InMux
    port map (
            O => \N__6681\,
            I => \N__6672\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__6678\,
            I => \N__6669\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__6675\,
            I => \N__6666\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__6672\,
            I => \N__6663\
        );

    \I__1679\ : Span4Mux_v
    port map (
            O => \N__6669\,
            I => \N__6658\
        );

    \I__1678\ : Span4Mux_v
    port map (
            O => \N__6666\,
            I => \N__6658\
        );

    \I__1677\ : Span4Mux_v
    port map (
            O => \N__6663\,
            I => \N__6655\
        );

    \I__1676\ : Sp12to4
    port map (
            O => \N__6658\,
            I => \N__6650\
        );

    \I__1675\ : Sp12to4
    port map (
            O => \N__6655\,
            I => \N__6650\
        );

    \I__1674\ : Span12Mux_h
    port map (
            O => \N__6650\,
            I => \N__6647\
        );

    \I__1673\ : Odrv12
    port map (
            O => \N__6647\,
            I => \D_UU_AMIGA_in_7\
        );

    \I__1672\ : IoInMux
    port map (
            O => \N__6644\,
            I => \N__6641\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__6641\,
            I => \N__6638\
        );

    \I__1670\ : Span12Mux_s10_v
    port map (
            O => \N__6638\,
            I => \N__6635\
        );

    \I__1669\ : Span12Mux_h
    port map (
            O => \N__6635\,
            I => \N__6632\
        );

    \I__1668\ : Odrv12
    port map (
            O => \N__6632\,
            I => \un1_D_UU_AMIGA_7\
        );

    \I__1667\ : IoInMux
    port map (
            O => \N__6629\,
            I => \N__6626\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__6626\,
            I => \N__6623\
        );

    \I__1665\ : Span4Mux_s2_h
    port map (
            O => \N__6623\,
            I => \N__6620\
        );

    \I__1664\ : Span4Mux_h
    port map (
            O => \N__6620\,
            I => \N__6617\
        );

    \I__1663\ : Span4Mux_h
    port map (
            O => \N__6617\,
            I => \N__6614\
        );

    \I__1662\ : Span4Mux_h
    port map (
            O => \N__6614\,
            I => \N__6611\
        );

    \I__1661\ : Odrv4
    port map (
            O => \N__6611\,
            I => \un1_D_UM_AMIGA_0\
        );

    \I__1660\ : IoInMux
    port map (
            O => \N__6608\,
            I => \N__6605\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__6605\,
            I => \N__6602\
        );

    \I__1658\ : Span4Mux_s2_h
    port map (
            O => \N__6602\,
            I => \N__6599\
        );

    \I__1657\ : Span4Mux_h
    port map (
            O => \N__6599\,
            I => \N__6596\
        );

    \I__1656\ : Sp12to4
    port map (
            O => \N__6596\,
            I => \N__6593\
        );

    \I__1655\ : Span12Mux_v
    port map (
            O => \N__6593\,
            I => \N__6590\
        );

    \I__1654\ : Odrv12
    port map (
            O => \N__6590\,
            I => \un1_D_UM_AMIGA_6\
        );

    \I__1653\ : InMux
    port map (
            O => \N__6587\,
            I => \N__6583\
        );

    \I__1652\ : InMux
    port map (
            O => \N__6586\,
            I => \N__6579\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__6583\,
            I => \N__6576\
        );

    \I__1650\ : InMux
    port map (
            O => \N__6582\,
            I => \N__6573\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__6579\,
            I => \N__6570\
        );

    \I__1648\ : Span4Mux_h
    port map (
            O => \N__6576\,
            I => \N__6567\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__6573\,
            I => \N__6564\
        );

    \I__1646\ : Sp12to4
    port map (
            O => \N__6570\,
            I => \N__6561\
        );

    \I__1645\ : Sp12to4
    port map (
            O => \N__6567\,
            I => \N__6558\
        );

    \I__1644\ : Span12Mux_h
    port map (
            O => \N__6564\,
            I => \N__6553\
        );

    \I__1643\ : Span12Mux_v
    port map (
            O => \N__6561\,
            I => \N__6553\
        );

    \I__1642\ : Span12Mux_v
    port map (
            O => \N__6558\,
            I => \N__6550\
        );

    \I__1641\ : Span12Mux_v
    port map (
            O => \N__6553\,
            I => \N__6547\
        );

    \I__1640\ : Span12Mux_h
    port map (
            O => \N__6550\,
            I => \N__6544\
        );

    \I__1639\ : Odrv12
    port map (
            O => \N__6547\,
            I => \D_UM_AMIGA_in_6\
        );

    \I__1638\ : Odrv12
    port map (
            O => \N__6544\,
            I => \D_UM_AMIGA_in_6\
        );

    \I__1637\ : InMux
    port map (
            O => \N__6539\,
            I => \N__6536\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__6536\,
            I => \N__6533\
        );

    \I__1635\ : Odrv4
    port map (
            O => \N__6533\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\
        );

    \I__1634\ : CascadeMux
    port map (
            O => \N__6530\,
            I => \N__6527\
        );

    \I__1633\ : InMux
    port map (
            O => \N__6527\,
            I => \N__6524\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__6524\,
            I => \N__6521\
        );

    \I__1631\ : Span4Mux_v
    port map (
            O => \N__6521\,
            I => \N__6517\
        );

    \I__1630\ : InMux
    port map (
            O => \N__6520\,
            I => \N__6514\
        );

    \I__1629\ : Span4Mux_v
    port map (
            O => \N__6517\,
            I => \N__6511\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__6514\,
            I => \N__6508\
        );

    \I__1627\ : Span4Mux_v
    port map (
            O => \N__6511\,
            I => \N__6502\
        );

    \I__1626\ : Span4Mux_v
    port map (
            O => \N__6508\,
            I => \N__6502\
        );

    \I__1625\ : InMux
    port map (
            O => \N__6507\,
            I => \N__6499\
        );

    \I__1624\ : Sp12to4
    port map (
            O => \N__6502\,
            I => \N__6494\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__6499\,
            I => \N__6494\
        );

    \I__1622\ : Span12Mux_h
    port map (
            O => \N__6494\,
            I => \N__6491\
        );

    \I__1621\ : Odrv12
    port map (
            O => \N__6491\,
            I => \D_UM_AMIGA_in_0\
        );

    \I__1620\ : InMux
    port map (
            O => \N__6488\,
            I => \N__6485\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__6485\,
            I => \N__6482\
        );

    \I__1618\ : Odrv4
    port map (
            O => \N__6482\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\
        );

    \I__1617\ : InMux
    port map (
            O => \N__6479\,
            I => \N__6476\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__6476\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa\
        );

    \I__1615\ : InMux
    port map (
            O => \N__6473\,
            I => \N__6470\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__6470\,
            I => \N__6467\
        );

    \I__1613\ : Odrv4
    port map (
            O => \N__6467\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\
        );

    \I__1612\ : InMux
    port map (
            O => \N__6464\,
            I => \N__6460\
        );

    \I__1611\ : InMux
    port map (
            O => \N__6463\,
            I => \N__6457\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__6460\,
            I => \N__6453\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__6457\,
            I => \N__6450\
        );

    \I__1608\ : InMux
    port map (
            O => \N__6456\,
            I => \N__6447\
        );

    \I__1607\ : Span4Mux_h
    port map (
            O => \N__6453\,
            I => \N__6444\
        );

    \I__1606\ : Span4Mux_v
    port map (
            O => \N__6450\,
            I => \N__6439\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__6447\,
            I => \N__6439\
        );

    \I__1604\ : Span4Mux_h
    port map (
            O => \N__6444\,
            I => \N__6436\
        );

    \I__1603\ : Span4Mux_v
    port map (
            O => \N__6439\,
            I => \N__6433\
        );

    \I__1602\ : Sp12to4
    port map (
            O => \N__6436\,
            I => \N__6430\
        );

    \I__1601\ : Sp12to4
    port map (
            O => \N__6433\,
            I => \N__6427\
        );

    \I__1600\ : Span12Mux_v
    port map (
            O => \N__6430\,
            I => \N__6424\
        );

    \I__1599\ : Span12Mux_h
    port map (
            O => \N__6427\,
            I => \N__6421\
        );

    \I__1598\ : Odrv12
    port map (
            O => \N__6424\,
            I => \D_UU_AMIGA_in_0\
        );

    \I__1597\ : Odrv12
    port map (
            O => \N__6421\,
            I => \D_UU_AMIGA_in_0\
        );

    \I__1596\ : IoInMux
    port map (
            O => \N__6416\,
            I => \N__6413\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__6413\,
            I => \N__6410\
        );

    \I__1594\ : Span12Mux_s7_v
    port map (
            O => \N__6410\,
            I => \N__6407\
        );

    \I__1593\ : Span12Mux_h
    port map (
            O => \N__6407\,
            I => \N__6404\
        );

    \I__1592\ : Odrv12
    port map (
            O => \N__6404\,
            I => \un1_D_UU_AMIGA_0\
        );

    \I__1591\ : InMux
    port map (
            O => \N__6401\,
            I => \N__6398\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__6398\,
            I => \N__6395\
        );

    \I__1589\ : Odrv4
    port map (
            O => \N__6395\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\
        );

    \I__1588\ : CascadeMux
    port map (
            O => \N__6392\,
            I => \N__6389\
        );

    \I__1587\ : InMux
    port map (
            O => \N__6389\,
            I => \N__6386\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__6386\,
            I => \N__6381\
        );

    \I__1585\ : InMux
    port map (
            O => \N__6385\,
            I => \N__6378\
        );

    \I__1584\ : InMux
    port map (
            O => \N__6384\,
            I => \N__6375\
        );

    \I__1583\ : Span4Mux_v
    port map (
            O => \N__6381\,
            I => \N__6372\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__6378\,
            I => \N__6367\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__6375\,
            I => \N__6367\
        );

    \I__1580\ : Sp12to4
    port map (
            O => \N__6372\,
            I => \N__6364\
        );

    \I__1579\ : Span4Mux_v
    port map (
            O => \N__6367\,
            I => \N__6361\
        );

    \I__1578\ : Span12Mux_h
    port map (
            O => \N__6364\,
            I => \N__6358\
        );

    \I__1577\ : Sp12to4
    port map (
            O => \N__6361\,
            I => \N__6355\
        );

    \I__1576\ : Span12Mux_v
    port map (
            O => \N__6358\,
            I => \N__6350\
        );

    \I__1575\ : Span12Mux_h
    port map (
            O => \N__6355\,
            I => \N__6350\
        );

    \I__1574\ : Odrv12
    port map (
            O => \N__6350\,
            I => \D_UM_AMIGA_in_5\
        );

    \I__1573\ : IoInMux
    port map (
            O => \N__6347\,
            I => \N__6344\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__6344\,
            I => \N__6341\
        );

    \I__1571\ : Span4Mux_s1_v
    port map (
            O => \N__6341\,
            I => \N__6338\
        );

    \I__1570\ : Sp12to4
    port map (
            O => \N__6338\,
            I => \N__6335\
        );

    \I__1569\ : Span12Mux_h
    port map (
            O => \N__6335\,
            I => \N__6332\
        );

    \I__1568\ : Odrv12
    port map (
            O => \N__6332\,
            I => \un1_D_UM_AMIGA_5\
        );

    \I__1567\ : InMux
    port map (
            O => \N__6329\,
            I => \N__6323\
        );

    \I__1566\ : InMux
    port map (
            O => \N__6328\,
            I => \N__6318\
        );

    \I__1565\ : InMux
    port map (
            O => \N__6327\,
            I => \N__6311\
        );

    \I__1564\ : InMux
    port map (
            O => \N__6326\,
            I => \N__6311\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__6323\,
            I => \N__6308\
        );

    \I__1562\ : InMux
    port map (
            O => \N__6322\,
            I => \N__6303\
        );

    \I__1561\ : InMux
    port map (
            O => \N__6321\,
            I => \N__6303\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__6318\,
            I => \N__6299\
        );

    \I__1559\ : InMux
    port map (
            O => \N__6317\,
            I => \N__6296\
        );

    \I__1558\ : InMux
    port map (
            O => \N__6316\,
            I => \N__6293\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__6311\,
            I => \N__6285\
        );

    \I__1556\ : Span4Mux_h
    port map (
            O => \N__6308\,
            I => \N__6279\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__6303\,
            I => \N__6279\
        );

    \I__1554\ : InMux
    port map (
            O => \N__6302\,
            I => \N__6276\
        );

    \I__1553\ : Span4Mux_h
    port map (
            O => \N__6299\,
            I => \N__6271\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__6296\,
            I => \N__6271\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__6293\,
            I => \N__6262\
        );

    \I__1550\ : InMux
    port map (
            O => \N__6292\,
            I => \N__6257\
        );

    \I__1549\ : InMux
    port map (
            O => \N__6291\,
            I => \N__6257\
        );

    \I__1548\ : InMux
    port map (
            O => \N__6290\,
            I => \N__6254\
        );

    \I__1547\ : InMux
    port map (
            O => \N__6289\,
            I => \N__6251\
        );

    \I__1546\ : CascadeMux
    port map (
            O => \N__6288\,
            I => \N__6248\
        );

    \I__1545\ : Span4Mux_v
    port map (
            O => \N__6285\,
            I => \N__6241\
        );

    \I__1544\ : InMux
    port map (
            O => \N__6284\,
            I => \N__6238\
        );

    \I__1543\ : Span4Mux_h
    port map (
            O => \N__6279\,
            I => \N__6234\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__6276\,
            I => \N__6231\
        );

    \I__1541\ : Span4Mux_h
    port map (
            O => \N__6271\,
            I => \N__6226\
        );

    \I__1540\ : InMux
    port map (
            O => \N__6270\,
            I => \N__6221\
        );

    \I__1539\ : InMux
    port map (
            O => \N__6269\,
            I => \N__6221\
        );

    \I__1538\ : InMux
    port map (
            O => \N__6268\,
            I => \N__6218\
        );

    \I__1537\ : InMux
    port map (
            O => \N__6267\,
            I => \N__6213\
        );

    \I__1536\ : InMux
    port map (
            O => \N__6266\,
            I => \N__6213\
        );

    \I__1535\ : InMux
    port map (
            O => \N__6265\,
            I => \N__6210\
        );

    \I__1534\ : Span4Mux_v
    port map (
            O => \N__6262\,
            I => \N__6207\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__6257\,
            I => \N__6204\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__6254\,
            I => \N__6201\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__6251\,
            I => \N__6198\
        );

    \I__1530\ : InMux
    port map (
            O => \N__6248\,
            I => \N__6195\
        );

    \I__1529\ : InMux
    port map (
            O => \N__6247\,
            I => \N__6188\
        );

    \I__1528\ : InMux
    port map (
            O => \N__6246\,
            I => \N__6188\
        );

    \I__1527\ : InMux
    port map (
            O => \N__6245\,
            I => \N__6188\
        );

    \I__1526\ : InMux
    port map (
            O => \N__6244\,
            I => \N__6185\
        );

    \I__1525\ : Span4Mux_v
    port map (
            O => \N__6241\,
            I => \N__6179\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__6238\,
            I => \N__6179\
        );

    \I__1523\ : InMux
    port map (
            O => \N__6237\,
            I => \N__6176\
        );

    \I__1522\ : Span4Mux_v
    port map (
            O => \N__6234\,
            I => \N__6171\
        );

    \I__1521\ : Span4Mux_h
    port map (
            O => \N__6231\,
            I => \N__6171\
        );

    \I__1520\ : InMux
    port map (
            O => \N__6230\,
            I => \N__6168\
        );

    \I__1519\ : InMux
    port map (
            O => \N__6229\,
            I => \N__6165\
        );

    \I__1518\ : Sp12to4
    port map (
            O => \N__6226\,
            I => \N__6158\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__6221\,
            I => \N__6158\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__6218\,
            I => \N__6155\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__6213\,
            I => \N__6152\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__6210\,
            I => \N__6149\
        );

    \I__1513\ : Span4Mux_v
    port map (
            O => \N__6207\,
            I => \N__6144\
        );

    \I__1512\ : Span4Mux_v
    port map (
            O => \N__6204\,
            I => \N__6144\
        );

    \I__1511\ : Span4Mux_v
    port map (
            O => \N__6201\,
            I => \N__6139\
        );

    \I__1510\ : Span4Mux_v
    port map (
            O => \N__6198\,
            I => \N__6139\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__6195\,
            I => \N__6134\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__6188\,
            I => \N__6134\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__6185\,
            I => \N__6131\
        );

    \I__1506\ : InMux
    port map (
            O => \N__6184\,
            I => \N__6128\
        );

    \I__1505\ : Span4Mux_h
    port map (
            O => \N__6179\,
            I => \N__6123\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__6176\,
            I => \N__6123\
        );

    \I__1503\ : Span4Mux_v
    port map (
            O => \N__6171\,
            I => \N__6118\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__6168\,
            I => \N__6118\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__6165\,
            I => \N__6115\
        );

    \I__1500\ : InMux
    port map (
            O => \N__6164\,
            I => \N__6110\
        );

    \I__1499\ : InMux
    port map (
            O => \N__6163\,
            I => \N__6110\
        );

    \I__1498\ : Span12Mux_v
    port map (
            O => \N__6158\,
            I => \N__6106\
        );

    \I__1497\ : Span12Mux_h
    port map (
            O => \N__6155\,
            I => \N__6101\
        );

    \I__1496\ : Span12Mux_h
    port map (
            O => \N__6152\,
            I => \N__6101\
        );

    \I__1495\ : Span4Mux_h
    port map (
            O => \N__6149\,
            I => \N__6098\
        );

    \I__1494\ : Span4Mux_h
    port map (
            O => \N__6144\,
            I => \N__6089\
        );

    \I__1493\ : Span4Mux_v
    port map (
            O => \N__6139\,
            I => \N__6089\
        );

    \I__1492\ : Span4Mux_v
    port map (
            O => \N__6134\,
            I => \N__6089\
        );

    \I__1491\ : Span4Mux_v
    port map (
            O => \N__6131\,
            I => \N__6089\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__6128\,
            I => \N__6086\
        );

    \I__1489\ : Span4Mux_h
    port map (
            O => \N__6123\,
            I => \N__6077\
        );

    \I__1488\ : Span4Mux_v
    port map (
            O => \N__6118\,
            I => \N__6077\
        );

    \I__1487\ : Span4Mux_v
    port map (
            O => \N__6115\,
            I => \N__6077\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__6110\,
            I => \N__6077\
        );

    \I__1485\ : InMux
    port map (
            O => \N__6109\,
            I => \N__6074\
        );

    \I__1484\ : Odrv12
    port map (
            O => \N__6106\,
            I => \U111_CYCLE_SM.un1_LW_TRANS_1_0\
        );

    \I__1483\ : Odrv12
    port map (
            O => \N__6101\,
            I => \U111_CYCLE_SM.un1_LW_TRANS_1_0\
        );

    \I__1482\ : Odrv4
    port map (
            O => \N__6098\,
            I => \U111_CYCLE_SM.un1_LW_TRANS_1_0\
        );

    \I__1481\ : Odrv4
    port map (
            O => \N__6089\,
            I => \U111_CYCLE_SM.un1_LW_TRANS_1_0\
        );

    \I__1480\ : Odrv12
    port map (
            O => \N__6086\,
            I => \U111_CYCLE_SM.un1_LW_TRANS_1_0\
        );

    \I__1479\ : Odrv4
    port map (
            O => \N__6077\,
            I => \U111_CYCLE_SM.un1_LW_TRANS_1_0\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__6074\,
            I => \U111_CYCLE_SM.un1_LW_TRANS_1_0\
        );

    \I__1477\ : InMux
    port map (
            O => \N__6059\,
            I => \N__6056\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__6056\,
            I => \N__6053\
        );

    \I__1475\ : Sp12to4
    port map (
            O => \N__6053\,
            I => \N__6050\
        );

    \I__1474\ : Span12Mux_v
    port map (
            O => \N__6050\,
            I => \N__6047\
        );

    \I__1473\ : Span12Mux_h
    port map (
            O => \N__6047\,
            I => \N__6044\
        );

    \I__1472\ : Odrv12
    port map (
            O => \N__6044\,
            I => \D_UU_040_in_6\
        );

    \I__1471\ : IoInMux
    port map (
            O => \N__6041\,
            I => \N__6037\
        );

    \I__1470\ : CascadeMux
    port map (
            O => \N__6040\,
            I => \N__6034\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__6037\,
            I => \N__6031\
        );

    \I__1468\ : InMux
    port map (
            O => \N__6034\,
            I => \N__6028\
        );

    \I__1467\ : Span4Mux_s2_h
    port map (
            O => \N__6031\,
            I => \N__6025\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__6028\,
            I => \N__6022\
        );

    \I__1465\ : Span4Mux_v
    port map (
            O => \N__6025\,
            I => \N__6019\
        );

    \I__1464\ : Span4Mux_v
    port map (
            O => \N__6022\,
            I => \N__6016\
        );

    \I__1463\ : Sp12to4
    port map (
            O => \N__6019\,
            I => \N__6013\
        );

    \I__1462\ : Span4Mux_v
    port map (
            O => \N__6016\,
            I => \N__6010\
        );

    \I__1461\ : Span12Mux_h
    port map (
            O => \N__6013\,
            I => \N__6007\
        );

    \I__1460\ : Sp12to4
    port map (
            O => \N__6010\,
            I => \N__6004\
        );

    \I__1459\ : Span12Mux_h
    port map (
            O => \N__6007\,
            I => \N__6001\
        );

    \I__1458\ : Span12Mux_h
    port map (
            O => \N__6004\,
            I => \N__5998\
        );

    \I__1457\ : Odrv12
    port map (
            O => \N__6001\,
            I => \D_LM_040_in_6\
        );

    \I__1456\ : Odrv12
    port map (
            O => \N__5998\,
            I => \D_LM_040_in_6\
        );

    \I__1455\ : InMux
    port map (
            O => \N__5993\,
            I => \N__5989\
        );

    \I__1454\ : InMux
    port map (
            O => \N__5992\,
            I => \N__5986\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__5989\,
            I => \N__5978\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__5986\,
            I => \N__5978\
        );

    \I__1451\ : InMux
    port map (
            O => \N__5985\,
            I => \N__5971\
        );

    \I__1450\ : InMux
    port map (
            O => \N__5984\,
            I => \N__5971\
        );

    \I__1449\ : InMux
    port map (
            O => \N__5983\,
            I => \N__5971\
        );

    \I__1448\ : Span4Mux_h
    port map (
            O => \N__5978\,
            I => \N__5961\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__5971\,
            I => \N__5961\
        );

    \I__1446\ : InMux
    port map (
            O => \N__5970\,
            I => \N__5958\
        );

    \I__1445\ : InMux
    port map (
            O => \N__5969\,
            I => \N__5950\
        );

    \I__1444\ : InMux
    port map (
            O => \N__5968\,
            I => \N__5950\
        );

    \I__1443\ : CascadeMux
    port map (
            O => \N__5967\,
            I => \N__5946\
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__5966\,
            I => \N__5942\
        );

    \I__1441\ : Span4Mux_v
    port map (
            O => \N__5961\,
            I => \N__5935\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__5958\,
            I => \N__5935\
        );

    \I__1439\ : InMux
    port map (
            O => \N__5957\,
            I => \N__5930\
        );

    \I__1438\ : InMux
    port map (
            O => \N__5956\,
            I => \N__5930\
        );

    \I__1437\ : InMux
    port map (
            O => \N__5955\,
            I => \N__5927\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__5950\,
            I => \N__5923\
        );

    \I__1435\ : InMux
    port map (
            O => \N__5949\,
            I => \N__5920\
        );

    \I__1434\ : InMux
    port map (
            O => \N__5946\,
            I => \N__5914\
        );

    \I__1433\ : InMux
    port map (
            O => \N__5945\,
            I => \N__5914\
        );

    \I__1432\ : InMux
    port map (
            O => \N__5942\,
            I => \N__5909\
        );

    \I__1431\ : CascadeMux
    port map (
            O => \N__5941\,
            I => \N__5906\
        );

    \I__1430\ : CascadeMux
    port map (
            O => \N__5940\,
            I => \N__5903\
        );

    \I__1429\ : Span4Mux_h
    port map (
            O => \N__5935\,
            I => \N__5898\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__5930\,
            I => \N__5898\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__5927\,
            I => \N__5895\
        );

    \I__1426\ : InMux
    port map (
            O => \N__5926\,
            I => \N__5892\
        );

    \I__1425\ : Span4Mux_h
    port map (
            O => \N__5923\,
            I => \N__5887\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__5920\,
            I => \N__5887\
        );

    \I__1423\ : InMux
    port map (
            O => \N__5919\,
            I => \N__5884\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__5914\,
            I => \N__5880\
        );

    \I__1421\ : InMux
    port map (
            O => \N__5913\,
            I => \N__5877\
        );

    \I__1420\ : InMux
    port map (
            O => \N__5912\,
            I => \N__5874\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__5909\,
            I => \N__5871\
        );

    \I__1418\ : InMux
    port map (
            O => \N__5906\,
            I => \N__5868\
        );

    \I__1417\ : InMux
    port map (
            O => \N__5903\,
            I => \N__5865\
        );

    \I__1416\ : Span4Mux_v
    port map (
            O => \N__5898\,
            I => \N__5861\
        );

    \I__1415\ : Span4Mux_v
    port map (
            O => \N__5895\,
            I => \N__5854\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__5892\,
            I => \N__5854\
        );

    \I__1413\ : Span4Mux_v
    port map (
            O => \N__5887\,
            I => \N__5846\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__5884\,
            I => \N__5846\
        );

    \I__1411\ : InMux
    port map (
            O => \N__5883\,
            I => \N__5843\
        );

    \I__1410\ : Span4Mux_v
    port map (
            O => \N__5880\,
            I => \N__5840\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__5877\,
            I => \N__5837\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__5874\,
            I => \N__5834\
        );

    \I__1407\ : Span4Mux_v
    port map (
            O => \N__5871\,
            I => \N__5826\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__5868\,
            I => \N__5826\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__5865\,
            I => \N__5826\
        );

    \I__1404\ : InMux
    port map (
            O => \N__5864\,
            I => \N__5823\
        );

    \I__1403\ : Span4Mux_v
    port map (
            O => \N__5861\,
            I => \N__5820\
        );

    \I__1402\ : InMux
    port map (
            O => \N__5860\,
            I => \N__5817\
        );

    \I__1401\ : InMux
    port map (
            O => \N__5859\,
            I => \N__5814\
        );

    \I__1400\ : Span4Mux_v
    port map (
            O => \N__5854\,
            I => \N__5811\
        );

    \I__1399\ : InMux
    port map (
            O => \N__5853\,
            I => \N__5806\
        );

    \I__1398\ : InMux
    port map (
            O => \N__5852\,
            I => \N__5806\
        );

    \I__1397\ : InMux
    port map (
            O => \N__5851\,
            I => \N__5803\
        );

    \I__1396\ : Span4Mux_v
    port map (
            O => \N__5846\,
            I => \N__5798\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__5843\,
            I => \N__5798\
        );

    \I__1394\ : Span4Mux_h
    port map (
            O => \N__5840\,
            I => \N__5790\
        );

    \I__1393\ : Span4Mux_v
    port map (
            O => \N__5837\,
            I => \N__5790\
        );

    \I__1392\ : Span12Mux_h
    port map (
            O => \N__5834\,
            I => \N__5787\
        );

    \I__1391\ : IoInMux
    port map (
            O => \N__5833\,
            I => \N__5784\
        );

    \I__1390\ : Span4Mux_v
    port map (
            O => \N__5826\,
            I => \N__5779\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__5823\,
            I => \N__5779\
        );

    \I__1388\ : Sp12to4
    port map (
            O => \N__5820\,
            I => \N__5770\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__5817\,
            I => \N__5770\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__5814\,
            I => \N__5770\
        );

    \I__1385\ : Sp12to4
    port map (
            O => \N__5811\,
            I => \N__5770\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__5806\,
            I => \N__5765\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__5803\,
            I => \N__5765\
        );

    \I__1382\ : Span4Mux_h
    port map (
            O => \N__5798\,
            I => \N__5762\
        );

    \I__1381\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5757\
        );

    \I__1380\ : InMux
    port map (
            O => \N__5796\,
            I => \N__5757\
        );

    \I__1379\ : InMux
    port map (
            O => \N__5795\,
            I => \N__5754\
        );

    \I__1378\ : Span4Mux_h
    port map (
            O => \N__5790\,
            I => \N__5751\
        );

    \I__1377\ : Span12Mux_v
    port map (
            O => \N__5787\,
            I => \N__5746\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__5784\,
            I => \N__5746\
        );

    \I__1375\ : Span4Mux_h
    port map (
            O => \N__5779\,
            I => \N__5743\
        );

    \I__1374\ : Span12Mux_h
    port map (
            O => \N__5770\,
            I => \N__5732\
        );

    \I__1373\ : Span12Mux_v
    port map (
            O => \N__5765\,
            I => \N__5732\
        );

    \I__1372\ : Sp12to4
    port map (
            O => \N__5762\,
            I => \N__5732\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__5757\,
            I => \N__5732\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__5754\,
            I => \N__5732\
        );

    \I__1369\ : Odrv4
    port map (
            O => \N__5751\,
            I => \A_AMIGA_c_1\
        );

    \I__1368\ : Odrv12
    port map (
            O => \N__5746\,
            I => \A_AMIGA_c_1\
        );

    \I__1367\ : Odrv4
    port map (
            O => \N__5743\,
            I => \A_AMIGA_c_1\
        );

    \I__1366\ : Odrv12
    port map (
            O => \N__5732\,
            I => \A_AMIGA_c_1\
        );

    \I__1365\ : IoInMux
    port map (
            O => \N__5723\,
            I => \N__5720\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__5720\,
            I => \N__5717\
        );

    \I__1363\ : Span12Mux_s10_v
    port map (
            O => \N__5717\,
            I => \N__5714\
        );

    \I__1362\ : Span12Mux_h
    port map (
            O => \N__5714\,
            I => \N__5711\
        );

    \I__1361\ : Odrv12
    port map (
            O => \N__5711\,
            I => \un1_D_UU_040_6\
        );

    \I__1360\ : CascadeMux
    port map (
            O => \N__5708\,
            I => \N__5705\
        );

    \I__1359\ : InMux
    port map (
            O => \N__5705\,
            I => \N__5702\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__5702\,
            I => \N__5697\
        );

    \I__1357\ : InMux
    port map (
            O => \N__5701\,
            I => \N__5694\
        );

    \I__1356\ : InMux
    port map (
            O => \N__5700\,
            I => \N__5691\
        );

    \I__1355\ : Span4Mux_v
    port map (
            O => \N__5697\,
            I => \N__5686\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__5694\,
            I => \N__5686\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__5691\,
            I => \N__5683\
        );

    \I__1352\ : Span4Mux_v
    port map (
            O => \N__5686\,
            I => \N__5678\
        );

    \I__1351\ : Span4Mux_v
    port map (
            O => \N__5683\,
            I => \N__5678\
        );

    \I__1350\ : Sp12to4
    port map (
            O => \N__5678\,
            I => \N__5675\
        );

    \I__1349\ : Span12Mux_h
    port map (
            O => \N__5675\,
            I => \N__5672\
        );

    \I__1348\ : Odrv12
    port map (
            O => \N__5672\,
            I => \D_UU_AMIGA_in_4\
        );

    \I__1347\ : InMux
    port map (
            O => \N__5669\,
            I => \N__5666\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__5666\,
            I => \N__5663\
        );

    \I__1345\ : Odrv12
    port map (
            O => \N__5663\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\
        );

    \I__1344\ : IoInMux
    port map (
            O => \N__5660\,
            I => \N__5657\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__5657\,
            I => \N__5654\
        );

    \I__1342\ : Span4Mux_s2_v
    port map (
            O => \N__5654\,
            I => \N__5651\
        );

    \I__1341\ : Span4Mux_h
    port map (
            O => \N__5651\,
            I => \N__5648\
        );

    \I__1340\ : Span4Mux_h
    port map (
            O => \N__5648\,
            I => \N__5645\
        );

    \I__1339\ : Span4Mux_v
    port map (
            O => \N__5645\,
            I => \N__5642\
        );

    \I__1338\ : Odrv4
    port map (
            O => \N__5642\,
            I => \un1_D_UU_AMIGA_4\
        );

    \I__1337\ : InMux
    port map (
            O => \N__5639\,
            I => \N__5636\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__5636\,
            I => \N__5633\
        );

    \I__1335\ : Glb2LocalMux
    port map (
            O => \N__5633\,
            I => \N__5600\
        );

    \I__1334\ : ClkMux
    port map (
            O => \N__5632\,
            I => \N__5600\
        );

    \I__1333\ : ClkMux
    port map (
            O => \N__5631\,
            I => \N__5600\
        );

    \I__1332\ : ClkMux
    port map (
            O => \N__5630\,
            I => \N__5600\
        );

    \I__1331\ : ClkMux
    port map (
            O => \N__5629\,
            I => \N__5600\
        );

    \I__1330\ : ClkMux
    port map (
            O => \N__5628\,
            I => \N__5600\
        );

    \I__1329\ : ClkMux
    port map (
            O => \N__5627\,
            I => \N__5600\
        );

    \I__1328\ : ClkMux
    port map (
            O => \N__5626\,
            I => \N__5600\
        );

    \I__1327\ : ClkMux
    port map (
            O => \N__5625\,
            I => \N__5600\
        );

    \I__1326\ : ClkMux
    port map (
            O => \N__5624\,
            I => \N__5600\
        );

    \I__1325\ : ClkMux
    port map (
            O => \N__5623\,
            I => \N__5600\
        );

    \I__1324\ : GlobalMux
    port map (
            O => \N__5600\,
            I => \CLK80\
        );

    \I__1323\ : IoInMux
    port map (
            O => \N__5597\,
            I => \N__5594\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__5594\,
            I => \N__5590\
        );

    \I__1321\ : IoInMux
    port map (
            O => \N__5593\,
            I => \N__5587\
        );

    \I__1320\ : IoSpan4Mux
    port map (
            O => \N__5590\,
            I => \N__5584\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__5587\,
            I => \N__5580\
        );

    \I__1318\ : IoSpan4Mux
    port map (
            O => \N__5584\,
            I => \N__5577\
        );

    \I__1317\ : IoInMux
    port map (
            O => \N__5583\,
            I => \N__5574\
        );

    \I__1316\ : IoSpan4Mux
    port map (
            O => \N__5580\,
            I => \N__5571\
        );

    \I__1315\ : Sp12to4
    port map (
            O => \N__5577\,
            I => \N__5566\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__5574\,
            I => \N__5566\
        );

    \I__1313\ : Span4Mux_s2_h
    port map (
            O => \N__5571\,
            I => \N__5563\
        );

    \I__1312\ : Span12Mux_s9_v
    port map (
            O => \N__5566\,
            I => \N__5560\
        );

    \I__1311\ : Sp12to4
    port map (
            O => \N__5563\,
            I => \N__5557\
        );

    \I__1310\ : Odrv12
    port map (
            O => \N__5560\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__1309\ : Odrv12
    port map (
            O => \N__5557\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__1308\ : InMux
    port map (
            O => \N__5552\,
            I => \N__5549\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__5549\,
            I => \U111_CYCLE_SM.A_OUT_0_sqmuxa_0_a3_0\
        );

    \I__1306\ : InMux
    port map (
            O => \N__5546\,
            I => \N__5540\
        );

    \I__1305\ : InMux
    port map (
            O => \N__5545\,
            I => \N__5537\
        );

    \I__1304\ : InMux
    port map (
            O => \N__5544\,
            I => \N__5532\
        );

    \I__1303\ : InMux
    port map (
            O => \N__5543\,
            I => \N__5532\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__5540\,
            I => \N__5528\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__5537\,
            I => \N__5525\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__5532\,
            I => \N__5522\
        );

    \I__1299\ : ClkMux
    port map (
            O => \N__5531\,
            I => \N__5513\
        );

    \I__1298\ : Glb2LocalMux
    port map (
            O => \N__5528\,
            I => \N__5513\
        );

    \I__1297\ : Glb2LocalMux
    port map (
            O => \N__5525\,
            I => \N__5513\
        );

    \I__1296\ : Glb2LocalMux
    port map (
            O => \N__5522\,
            I => \N__5513\
        );

    \I__1295\ : GlobalMux
    port map (
            O => \N__5513\,
            I => \CLK40\
        );

    \I__1294\ : CascadeMux
    port map (
            O => \N__5510\,
            I => \U111_CYCLE_SM.N_91_cascade_\
        );

    \I__1293\ : InMux
    port map (
            O => \N__5507\,
            I => \N__5504\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__5504\,
            I => \N__5497\
        );

    \I__1291\ : InMux
    port map (
            O => \N__5503\,
            I => \N__5494\
        );

    \I__1290\ : InMux
    port map (
            O => \N__5502\,
            I => \N__5489\
        );

    \I__1289\ : InMux
    port map (
            O => \N__5501\,
            I => \N__5489\
        );

    \I__1288\ : InMux
    port map (
            O => \N__5500\,
            I => \N__5486\
        );

    \I__1287\ : Odrv4
    port map (
            O => \N__5497\,
            I => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__5494\,
            I => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__5489\,
            I => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__5486\,
            I => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\
        );

    \I__1283\ : CascadeMux
    port map (
            O => \N__5477\,
            I => \U111_CYCLE_SM.A_OUT_0_cascade_\
        );

    \I__1282\ : InMux
    port map (
            O => \N__5474\,
            I => \N__5471\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__5471\,
            I => \N__5468\
        );

    \I__1280\ : Span4Mux_v
    port map (
            O => \N__5468\,
            I => \N__5465\
        );

    \I__1279\ : Sp12to4
    port map (
            O => \N__5465\,
            I => \N__5462\
        );

    \I__1278\ : Span12Mux_h
    port map (
            O => \N__5462\,
            I => \N__5459\
        );

    \I__1277\ : Span12Mux_v
    port map (
            O => \N__5459\,
            I => \N__5455\
        );

    \I__1276\ : InMux
    port map (
            O => \N__5458\,
            I => \N__5452\
        );

    \I__1275\ : Odrv12
    port map (
            O => \N__5455\,
            I => \U111_CYCLE_SM.A_OUTZ0\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__5452\,
            I => \U111_CYCLE_SM.A_OUTZ0\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__5447\,
            I => \N__5441\
        );

    \I__1272\ : InMux
    port map (
            O => \N__5446\,
            I => \N__5434\
        );

    \I__1271\ : InMux
    port map (
            O => \N__5445\,
            I => \N__5434\
        );

    \I__1270\ : InMux
    port map (
            O => \N__5444\,
            I => \N__5434\
        );

    \I__1269\ : InMux
    port map (
            O => \N__5441\,
            I => \N__5431\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__5434\,
            I => \N__5426\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__5431\,
            I => \N__5426\
        );

    \I__1266\ : Span4Mux_v
    port map (
            O => \N__5426\,
            I => \N__5422\
        );

    \I__1265\ : InMux
    port map (
            O => \N__5425\,
            I => \N__5419\
        );

    \I__1264\ : Sp12to4
    port map (
            O => \N__5422\,
            I => \N__5414\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__5419\,
            I => \N__5414\
        );

    \I__1262\ : Span12Mux_h
    port map (
            O => \N__5414\,
            I => \N__5411\
        );

    \I__1261\ : Span12Mux_v
    port map (
            O => \N__5411\,
            I => \N__5408\
        );

    \I__1260\ : Odrv12
    port map (
            O => \N__5408\,
            I => \TACKn_c\
        );

    \I__1259\ : InMux
    port map (
            O => \N__5405\,
            I => \N__5402\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__5402\,
            I => \N__5391\
        );

    \I__1257\ : InMux
    port map (
            O => \N__5401\,
            I => \N__5386\
        );

    \I__1256\ : InMux
    port map (
            O => \N__5400\,
            I => \N__5386\
        );

    \I__1255\ : InMux
    port map (
            O => \N__5399\,
            I => \N__5381\
        );

    \I__1254\ : InMux
    port map (
            O => \N__5398\,
            I => \N__5381\
        );

    \I__1253\ : InMux
    port map (
            O => \N__5397\,
            I => \N__5372\
        );

    \I__1252\ : InMux
    port map (
            O => \N__5396\,
            I => \N__5372\
        );

    \I__1251\ : InMux
    port map (
            O => \N__5395\,
            I => \N__5372\
        );

    \I__1250\ : InMux
    port map (
            O => \N__5394\,
            I => \N__5372\
        );

    \I__1249\ : Odrv4
    port map (
            O => \N__5391\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__5386\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__5381\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__5372\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1245\ : InMux
    port map (
            O => \N__5363\,
            I => \N__5358\
        );

    \I__1244\ : CascadeMux
    port map (
            O => \N__5362\,
            I => \N__5351\
        );

    \I__1243\ : CascadeMux
    port map (
            O => \N__5361\,
            I => \N__5347\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__5358\,
            I => \N__5343\
        );

    \I__1241\ : InMux
    port map (
            O => \N__5357\,
            I => \N__5338\
        );

    \I__1240\ : InMux
    port map (
            O => \N__5356\,
            I => \N__5338\
        );

    \I__1239\ : InMux
    port map (
            O => \N__5355\,
            I => \N__5333\
        );

    \I__1238\ : InMux
    port map (
            O => \N__5354\,
            I => \N__5333\
        );

    \I__1237\ : InMux
    port map (
            O => \N__5351\,
            I => \N__5324\
        );

    \I__1236\ : InMux
    port map (
            O => \N__5350\,
            I => \N__5324\
        );

    \I__1235\ : InMux
    port map (
            O => \N__5347\,
            I => \N__5324\
        );

    \I__1234\ : InMux
    port map (
            O => \N__5346\,
            I => \N__5324\
        );

    \I__1233\ : Odrv4
    port map (
            O => \N__5343\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__5338\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__5333\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__5324\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1229\ : CascadeMux
    port map (
            O => \N__5315\,
            I => \N__5306\
        );

    \I__1228\ : InMux
    port map (
            O => \N__5314\,
            I => \N__5303\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5313\,
            I => \N__5296\
        );

    \I__1226\ : InMux
    port map (
            O => \N__5312\,
            I => \N__5296\
        );

    \I__1225\ : InMux
    port map (
            O => \N__5311\,
            I => \N__5296\
        );

    \I__1224\ : InMux
    port map (
            O => \N__5310\,
            I => \N__5291\
        );

    \I__1223\ : InMux
    port map (
            O => \N__5309\,
            I => \N__5291\
        );

    \I__1222\ : InMux
    port map (
            O => \N__5306\,
            I => \N__5288\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__5303\,
            I => \N__5278\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__5296\,
            I => \N__5278\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__5291\,
            I => \N__5278\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__5288\,
            I => \N__5278\
        );

    \I__1217\ : InMux
    port map (
            O => \N__5287\,
            I => \N__5275\
        );

    \I__1216\ : Span4Mux_v
    port map (
            O => \N__5278\,
            I => \N__5270\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__5275\,
            I => \N__5270\
        );

    \I__1214\ : Span4Mux_h
    port map (
            O => \N__5270\,
            I => \N__5267\
        );

    \I__1213\ : Span4Mux_v
    port map (
            O => \N__5267\,
            I => \N__5263\
        );

    \I__1212\ : InMux
    port map (
            O => \N__5266\,
            I => \N__5260\
        );

    \I__1211\ : Sp12to4
    port map (
            O => \N__5263\,
            I => \N__5255\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__5260\,
            I => \N__5255\
        );

    \I__1209\ : Span12Mux_v
    port map (
            O => \N__5255\,
            I => \N__5252\
        );

    \I__1208\ : Odrv12
    port map (
            O => \N__5252\,
            I => \RESETn_c\
        );

    \I__1207\ : CascadeMux
    port map (
            O => \N__5249\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_\
        );

    \I__1206\ : IoInMux
    port map (
            O => \N__5246\,
            I => \N__5242\
        );

    \I__1205\ : IoInMux
    port map (
            O => \N__5245\,
            I => \N__5239\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__5242\,
            I => \N__5231\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__5239\,
            I => \N__5231\
        );

    \I__1202\ : IoInMux
    port map (
            O => \N__5238\,
            I => \N__5228\
        );

    \I__1201\ : IoInMux
    port map (
            O => \N__5237\,
            I => \N__5225\
        );

    \I__1200\ : IoInMux
    port map (
            O => \N__5236\,
            I => \N__5217\
        );

    \I__1199\ : IoSpan4Mux
    port map (
            O => \N__5231\,
            I => \N__5210\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__5228\,
            I => \N__5210\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__5225\,
            I => \N__5210\
        );

    \I__1196\ : IoInMux
    port map (
            O => \N__5224\,
            I => \N__5207\
        );

    \I__1195\ : IoInMux
    port map (
            O => \N__5223\,
            I => \N__5204\
        );

    \I__1194\ : IoInMux
    port map (
            O => \N__5222\,
            I => \N__5201\
        );

    \I__1193\ : IoInMux
    port map (
            O => \N__5221\,
            I => \N__5198\
        );

    \I__1192\ : IoInMux
    port map (
            O => \N__5220\,
            I => \N__5195\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__5217\,
            I => \N__5190\
        );

    \I__1190\ : IoSpan4Mux
    port map (
            O => \N__5210\,
            I => \N__5175\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5207\,
            I => \N__5175\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__5204\,
            I => \N__5175\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__5201\,
            I => \N__5175\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__5198\,
            I => \N__5175\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__5195\,
            I => \N__5175\
        );

    \I__1184\ : IoInMux
    port map (
            O => \N__5194\,
            I => \N__5172\
        );

    \I__1183\ : IoInMux
    port map (
            O => \N__5193\,
            I => \N__5169\
        );

    \I__1182\ : Span4Mux_s3_v
    port map (
            O => \N__5190\,
            I => \N__5166\
        );

    \I__1181\ : IoInMux
    port map (
            O => \N__5189\,
            I => \N__5162\
        );

    \I__1180\ : IoInMux
    port map (
            O => \N__5188\,
            I => \N__5159\
        );

    \I__1179\ : IoSpan4Mux
    port map (
            O => \N__5175\,
            I => \N__5146\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__5172\,
            I => \N__5146\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__5169\,
            I => \N__5146\
        );

    \I__1176\ : Span4Mux_h
    port map (
            O => \N__5166\,
            I => \N__5142\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5165\,
            I => \N__5139\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__5162\,
            I => \N__5134\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__5159\,
            I => \N__5134\
        );

    \I__1172\ : IoInMux
    port map (
            O => \N__5158\,
            I => \N__5131\
        );

    \I__1171\ : IoInMux
    port map (
            O => \N__5157\,
            I => \N__5128\
        );

    \I__1170\ : IoInMux
    port map (
            O => \N__5156\,
            I => \N__5125\
        );

    \I__1169\ : IoInMux
    port map (
            O => \N__5155\,
            I => \N__5122\
        );

    \I__1168\ : IoInMux
    port map (
            O => \N__5154\,
            I => \N__5119\
        );

    \I__1167\ : IoInMux
    port map (
            O => \N__5153\,
            I => \N__5116\
        );

    \I__1166\ : IoSpan4Mux
    port map (
            O => \N__5146\,
            I => \N__5109\
        );

    \I__1165\ : IoInMux
    port map (
            O => \N__5145\,
            I => \N__5106\
        );

    \I__1164\ : Span4Mux_v
    port map (
            O => \N__5142\,
            I => \N__5100\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__5139\,
            I => \N__5100\
        );

    \I__1162\ : IoSpan4Mux
    port map (
            O => \N__5134\,
            I => \N__5083\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__5131\,
            I => \N__5083\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__5128\,
            I => \N__5083\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__5125\,
            I => \N__5083\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__5122\,
            I => \N__5083\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__5119\,
            I => \N__5083\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__5116\,
            I => \N__5083\
        );

    \I__1155\ : IoInMux
    port map (
            O => \N__5115\,
            I => \N__5080\
        );

    \I__1154\ : IoInMux
    port map (
            O => \N__5114\,
            I => \N__5077\
        );

    \I__1153\ : IoInMux
    port map (
            O => \N__5113\,
            I => \N__5074\
        );

    \I__1152\ : IoInMux
    port map (
            O => \N__5112\,
            I => \N__5071\
        );

    \I__1151\ : IoSpan4Mux
    port map (
            O => \N__5109\,
            I => \N__5066\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__5106\,
            I => \N__5066\
        );

    \I__1149\ : IoInMux
    port map (
            O => \N__5105\,
            I => \N__5063\
        );

    \I__1148\ : Span4Mux_v
    port map (
            O => \N__5100\,
            I => \N__5057\
        );

    \I__1147\ : IoInMux
    port map (
            O => \N__5099\,
            I => \N__5054\
        );

    \I__1146\ : InMux
    port map (
            O => \N__5098\,
            I => \N__5051\
        );

    \I__1145\ : IoSpan4Mux
    port map (
            O => \N__5083\,
            I => \N__5040\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__5080\,
            I => \N__5040\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__5077\,
            I => \N__5040\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__5074\,
            I => \N__5040\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__5071\,
            I => \N__5040\
        );

    \I__1140\ : IoSpan4Mux
    port map (
            O => \N__5066\,
            I => \N__5036\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__5063\,
            I => \N__5033\
        );

    \I__1138\ : IoInMux
    port map (
            O => \N__5062\,
            I => \N__5030\
        );

    \I__1137\ : IoInMux
    port map (
            O => \N__5061\,
            I => \N__5027\
        );

    \I__1136\ : IoInMux
    port map (
            O => \N__5060\,
            I => \N__5024\
        );

    \I__1135\ : Sp12to4
    port map (
            O => \N__5057\,
            I => \N__5019\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__5054\,
            I => \N__5016\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__5051\,
            I => \N__5013\
        );

    \I__1132\ : IoSpan4Mux
    port map (
            O => \N__5040\,
            I => \N__5010\
        );

    \I__1131\ : IoInMux
    port map (
            O => \N__5039\,
            I => \N__5007\
        );

    \I__1130\ : IoSpan4Mux
    port map (
            O => \N__5036\,
            I => \N__4996\
        );

    \I__1129\ : IoSpan4Mux
    port map (
            O => \N__5033\,
            I => \N__4996\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__5030\,
            I => \N__4996\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__5027\,
            I => \N__4996\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__5024\,
            I => \N__4996\
        );

    \I__1125\ : IoInMux
    port map (
            O => \N__5023\,
            I => \N__4993\
        );

    \I__1124\ : IoInMux
    port map (
            O => \N__5022\,
            I => \N__4990\
        );

    \I__1123\ : Span12Mux_h
    port map (
            O => \N__5019\,
            I => \N__4987\
        );

    \I__1122\ : Span12Mux_s11_v
    port map (
            O => \N__5016\,
            I => \N__4982\
        );

    \I__1121\ : Span12Mux_h
    port map (
            O => \N__5013\,
            I => \N__4982\
        );

    \I__1120\ : IoSpan4Mux
    port map (
            O => \N__5010\,
            I => \N__4977\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__5007\,
            I => \N__4977\
        );

    \I__1118\ : IoSpan4Mux
    port map (
            O => \N__4996\,
            I => \N__4972\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__4993\,
            I => \N__4972\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__4990\,
            I => \N__4969\
        );

    \I__1115\ : Odrv12
    port map (
            O => \N__4987\,
            I => \RnW_c\
        );

    \I__1114\ : Odrv12
    port map (
            O => \N__4982\,
            I => \RnW_c\
        );

    \I__1113\ : Odrv4
    port map (
            O => \N__4977\,
            I => \RnW_c\
        );

    \I__1112\ : Odrv4
    port map (
            O => \N__4972\,
            I => \RnW_c\
        );

    \I__1111\ : Odrv12
    port map (
            O => \N__4969\,
            I => \RnW_c\
        );

    \I__1110\ : CascadeMux
    port map (
            O => \N__4958\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0_cascade_\
        );

    \I__1109\ : InMux
    port map (
            O => \N__4955\,
            I => \N__4952\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__4952\,
            I => \N__4949\
        );

    \I__1107\ : Odrv4
    port map (
            O => \N__4949\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\
        );

    \I__1106\ : InMux
    port map (
            O => \N__4946\,
            I => \N__4941\
        );

    \I__1105\ : InMux
    port map (
            O => \N__4945\,
            I => \N__4938\
        );

    \I__1104\ : InMux
    port map (
            O => \N__4944\,
            I => \N__4935\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__4941\,
            I => \N__4930\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__4938\,
            I => \N__4930\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__4935\,
            I => \N__4927\
        );

    \I__1100\ : Span4Mux_v
    port map (
            O => \N__4930\,
            I => \N__4924\
        );

    \I__1099\ : Sp12to4
    port map (
            O => \N__4927\,
            I => \N__4921\
        );

    \I__1098\ : Sp12to4
    port map (
            O => \N__4924\,
            I => \N__4918\
        );

    \I__1097\ : Span12Mux_v
    port map (
            O => \N__4921\,
            I => \N__4915\
        );

    \I__1096\ : Span12Mux_h
    port map (
            O => \N__4918\,
            I => \N__4912\
        );

    \I__1095\ : Span12Mux_h
    port map (
            O => \N__4915\,
            I => \N__4909\
        );

    \I__1094\ : Odrv12
    port map (
            O => \N__4912\,
            I => \D_UU_AMIGA_in_6\
        );

    \I__1093\ : Odrv12
    port map (
            O => \N__4909\,
            I => \D_UU_AMIGA_in_6\
        );

    \I__1092\ : IoInMux
    port map (
            O => \N__4904\,
            I => \N__4901\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__4901\,
            I => \N__4898\
        );

    \I__1090\ : Span4Mux_s1_v
    port map (
            O => \N__4898\,
            I => \N__4895\
        );

    \I__1089\ : Span4Mux_v
    port map (
            O => \N__4895\,
            I => \N__4892\
        );

    \I__1088\ : Sp12to4
    port map (
            O => \N__4892\,
            I => \N__4889\
        );

    \I__1087\ : Span12Mux_h
    port map (
            O => \N__4889\,
            I => \N__4886\
        );

    \I__1086\ : Odrv12
    port map (
            O => \N__4886\,
            I => \un1_D_UU_AMIGA_6\
        );

    \I__1085\ : InMux
    port map (
            O => \N__4883\,
            I => \N__4880\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__4880\,
            I => \N__4877\
        );

    \I__1083\ : Odrv12
    port map (
            O => \N__4877\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\
        );

    \I__1082\ : CascadeMux
    port map (
            O => \N__4874\,
            I => \N__4871\
        );

    \I__1081\ : InMux
    port map (
            O => \N__4871\,
            I => \N__4868\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__4868\,
            I => \N__4863\
        );

    \I__1079\ : InMux
    port map (
            O => \N__4867\,
            I => \N__4860\
        );

    \I__1078\ : InMux
    port map (
            O => \N__4866\,
            I => \N__4857\
        );

    \I__1077\ : Span4Mux_v
    port map (
            O => \N__4863\,
            I => \N__4850\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__4860\,
            I => \N__4850\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__4857\,
            I => \N__4850\
        );

    \I__1074\ : Span4Mux_v
    port map (
            O => \N__4850\,
            I => \N__4847\
        );

    \I__1073\ : Sp12to4
    port map (
            O => \N__4847\,
            I => \N__4844\
        );

    \I__1072\ : Span12Mux_h
    port map (
            O => \N__4844\,
            I => \N__4841\
        );

    \I__1071\ : Odrv12
    port map (
            O => \N__4841\,
            I => \D_UU_AMIGA_in_2\
        );

    \I__1070\ : IoInMux
    port map (
            O => \N__4838\,
            I => \N__4835\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__4835\,
            I => \N__4832\
        );

    \I__1068\ : Span12Mux_s1_v
    port map (
            O => \N__4832\,
            I => \N__4829\
        );

    \I__1067\ : Span12Mux_h
    port map (
            O => \N__4829\,
            I => \N__4826\
        );

    \I__1066\ : Odrv12
    port map (
            O => \N__4826\,
            I => \un1_D_UU_AMIGA_2\
        );

    \I__1065\ : IoInMux
    port map (
            O => \N__4823\,
            I => \N__4818\
        );

    \I__1064\ : IoInMux
    port map (
            O => \N__4822\,
            I => \N__4815\
        );

    \I__1063\ : IoInMux
    port map (
            O => \N__4821\,
            I => \N__4812\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__4818\,
            I => \N__4809\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__4815\,
            I => \N__4806\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__4812\,
            I => \N__4803\
        );

    \I__1059\ : Span12Mux_s5_v
    port map (
            O => \N__4809\,
            I => \N__4800\
        );

    \I__1058\ : Span12Mux_s10_h
    port map (
            O => \N__4806\,
            I => \N__4795\
        );

    \I__1057\ : Span12Mux_s9_h
    port map (
            O => \N__4803\,
            I => \N__4795\
        );

    \I__1056\ : Odrv12
    port map (
            O => \N__4800\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__1055\ : Odrv12
    port map (
            O => \N__4795\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__1054\ : CascadeMux
    port map (
            O => \N__4790\,
            I => \N__4787\
        );

    \I__1053\ : InMux
    port map (
            O => \N__4787\,
            I => \N__4784\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__4784\,
            I => \N__4781\
        );

    \I__1051\ : Span12Mux_h
    port map (
            O => \N__4781\,
            I => \N__4778\
        );

    \I__1050\ : Odrv12
    port map (
            O => \N__4778\,
            I => \D_LM_AMIGA_in_1\
        );

    \I__1049\ : IoInMux
    port map (
            O => \N__4775\,
            I => \N__4772\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__4772\,
            I => \N__4769\
        );

    \I__1047\ : IoSpan4Mux
    port map (
            O => \N__4769\,
            I => \N__4766\
        );

    \I__1046\ : Span4Mux_s2_h
    port map (
            O => \N__4766\,
            I => \N__4763\
        );

    \I__1045\ : Sp12to4
    port map (
            O => \N__4763\,
            I => \N__4760\
        );

    \I__1044\ : Span12Mux_h
    port map (
            O => \N__4760\,
            I => \N__4757\
        );

    \I__1043\ : Odrv12
    port map (
            O => \N__4757\,
            I => \un1_D_LM_AMIGA_1\
        );

    \I__1042\ : InMux
    port map (
            O => \N__4754\,
            I => \N__4751\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__4751\,
            I => \N__4748\
        );

    \I__1040\ : Span4Mux_v
    port map (
            O => \N__4748\,
            I => \N__4745\
        );

    \I__1039\ : Sp12to4
    port map (
            O => \N__4745\,
            I => \N__4742\
        );

    \I__1038\ : Span12Mux_h
    port map (
            O => \N__4742\,
            I => \N__4739\
        );

    \I__1037\ : Odrv12
    port map (
            O => \N__4739\,
            I => \D_UM_040_in_6\
        );

    \I__1036\ : IoInMux
    port map (
            O => \N__4736\,
            I => \N__4733\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__4733\,
            I => \N__4729\
        );

    \I__1034\ : CascadeMux
    port map (
            O => \N__4732\,
            I => \N__4726\
        );

    \I__1033\ : IoSpan4Mux
    port map (
            O => \N__4729\,
            I => \N__4723\
        );

    \I__1032\ : InMux
    port map (
            O => \N__4726\,
            I => \N__4720\
        );

    \I__1031\ : IoSpan4Mux
    port map (
            O => \N__4723\,
            I => \N__4717\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__4720\,
            I => \N__4714\
        );

    \I__1029\ : Span4Mux_s2_h
    port map (
            O => \N__4717\,
            I => \N__4711\
        );

    \I__1028\ : Span4Mux_v
    port map (
            O => \N__4714\,
            I => \N__4708\
        );

    \I__1027\ : Sp12to4
    port map (
            O => \N__4711\,
            I => \N__4705\
        );

    \I__1026\ : Sp12to4
    port map (
            O => \N__4708\,
            I => \N__4702\
        );

    \I__1025\ : Span12Mux_h
    port map (
            O => \N__4705\,
            I => \N__4699\
        );

    \I__1024\ : Span12Mux_h
    port map (
            O => \N__4702\,
            I => \N__4696\
        );

    \I__1023\ : Span12Mux_h
    port map (
            O => \N__4699\,
            I => \N__4693\
        );

    \I__1022\ : Span12Mux_v
    port map (
            O => \N__4696\,
            I => \N__4690\
        );

    \I__1021\ : Odrv12
    port map (
            O => \N__4693\,
            I => \D_LL_040_in_6\
        );

    \I__1020\ : Odrv12
    port map (
            O => \N__4690\,
            I => \D_LL_040_in_6\
        );

    \I__1019\ : IoInMux
    port map (
            O => \N__4685\,
            I => \N__4682\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__4682\,
            I => \N__4679\
        );

    \I__1017\ : Span12Mux_s2_h
    port map (
            O => \N__4679\,
            I => \N__4676\
        );

    \I__1016\ : Span12Mux_v
    port map (
            O => \N__4676\,
            I => \N__4673\
        );

    \I__1015\ : Span12Mux_h
    port map (
            O => \N__4673\,
            I => \N__4670\
        );

    \I__1014\ : Odrv12
    port map (
            O => \N__4670\,
            I => \un1_D_UM_040_6\
        );

    \I__1013\ : CascadeMux
    port map (
            O => \N__4667\,
            I => \N__4663\
        );

    \I__1012\ : InMux
    port map (
            O => \N__4666\,
            I => \N__4660\
        );

    \I__1011\ : InMux
    port map (
            O => \N__4663\,
            I => \N__4657\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__4660\,
            I => \U111_CYCLE_SM.TA_ENZ0\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__4657\,
            I => \U111_CYCLE_SM.TA_ENZ0\
        );

    \I__1008\ : IoInMux
    port map (
            O => \N__4652\,
            I => \N__4649\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__4649\,
            I => \N__4646\
        );

    \I__1006\ : Span4Mux_s1_v
    port map (
            O => \N__4646\,
            I => \N__4643\
        );

    \I__1005\ : Span4Mux_v
    port map (
            O => \N__4643\,
            I => \N__4640\
        );

    \I__1004\ : Span4Mux_v
    port map (
            O => \N__4640\,
            I => \N__4637\
        );

    \I__1003\ : Span4Mux_v
    port map (
            O => \N__4637\,
            I => \N__4634\
        );

    \I__1002\ : Odrv4
    port map (
            O => \N__4634\,
            I => \U111_CYCLE_SM_TAn_0_i\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4631\,
            I => \N__4628\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__4628\,
            I => \N__4625\
        );

    \I__999\ : Span4Mux_v
    port map (
            O => \N__4625\,
            I => \N__4622\
        );

    \I__998\ : Sp12to4
    port map (
            O => \N__4622\,
            I => \N__4619\
        );

    \I__997\ : Span12Mux_h
    port map (
            O => \N__4619\,
            I => \N__4616\
        );

    \I__996\ : Odrv12
    port map (
            O => \N__4616\,
            I => \D_LM_AMIGA_in_4\
        );

    \I__995\ : IoInMux
    port map (
            O => \N__4613\,
            I => \N__4610\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__4610\,
            I => \N__4607\
        );

    \I__993\ : IoSpan4Mux
    port map (
            O => \N__4607\,
            I => \N__4604\
        );

    \I__992\ : Span4Mux_s2_h
    port map (
            O => \N__4604\,
            I => \N__4601\
        );

    \I__991\ : Sp12to4
    port map (
            O => \N__4601\,
            I => \N__4598\
        );

    \I__990\ : Span12Mux_h
    port map (
            O => \N__4598\,
            I => \N__4595\
        );

    \I__989\ : Odrv12
    port map (
            O => \N__4595\,
            I => \un1_D_LM_AMIGA_4\
        );

    \I__988\ : InMux
    port map (
            O => \N__4592\,
            I => \N__4589\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__4589\,
            I => \U111_CYCLE_SM.LW_CYCLE_0\
        );

    \I__986\ : CascadeMux
    port map (
            O => \N__4586\,
            I => \U111_CYCLE_SM.N_69_0_cascade_\
        );

    \I__985\ : InMux
    port map (
            O => \N__4583\,
            I => \N__4580\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__4580\,
            I => \U111_CYCLE_SM.TS_EN_5\
        );

    \I__983\ : InMux
    port map (
            O => \N__4577\,
            I => \N__4574\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__4574\,
            I => \N__4570\
        );

    \I__981\ : CascadeMux
    port map (
            O => \N__4573\,
            I => \N__4566\
        );

    \I__980\ : Span12Mux_s8_v
    port map (
            O => \N__4570\,
            I => \N__4563\
        );

    \I__979\ : InMux
    port map (
            O => \N__4569\,
            I => \N__4558\
        );

    \I__978\ : InMux
    port map (
            O => \N__4566\,
            I => \N__4558\
        );

    \I__977\ : Span12Mux_v
    port map (
            O => \N__4563\,
            I => \N__4555\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__4558\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__975\ : Odrv12
    port map (
            O => \N__4555\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__974\ : InMux
    port map (
            O => \N__4550\,
            I => \N__4547\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__4547\,
            I => \N__4544\
        );

    \I__972\ : Span4Mux_v
    port map (
            O => \N__4544\,
            I => \N__4540\
        );

    \I__971\ : InMux
    port map (
            O => \N__4543\,
            I => \N__4537\
        );

    \I__970\ : Sp12to4
    port map (
            O => \N__4540\,
            I => \N__4532\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__4537\,
            I => \N__4532\
        );

    \I__968\ : Span12Mux_h
    port map (
            O => \N__4532\,
            I => \N__4529\
        );

    \I__967\ : Span12Mux_v
    port map (
            O => \N__4529\,
            I => \N__4526\
        );

    \I__966\ : Odrv12
    port map (
            O => \N__4526\,
            I => \PORTSIZE_c\
        );

    \I__965\ : InMux
    port map (
            O => \N__4523\,
            I => \N__4520\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__4520\,
            I => \N__4516\
        );

    \I__963\ : InMux
    port map (
            O => \N__4519\,
            I => \N__4513\
        );

    \I__962\ : Span4Mux_h
    port map (
            O => \N__4516\,
            I => \N__4508\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__4513\,
            I => \N__4508\
        );

    \I__960\ : Span4Mux_v
    port map (
            O => \N__4508\,
            I => \N__4505\
        );

    \I__959\ : Sp12to4
    port map (
            O => \N__4505\,
            I => \N__4502\
        );

    \I__958\ : Span12Mux_h
    port map (
            O => \N__4502\,
            I => \N__4499\
        );

    \I__957\ : Odrv12
    port map (
            O => \N__4499\,
            I => \SIZ_c_1\
        );

    \I__956\ : InMux
    port map (
            O => \N__4496\,
            I => \N__4492\
        );

    \I__955\ : CascadeMux
    port map (
            O => \N__4495\,
            I => \N__4489\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__4492\,
            I => \N__4486\
        );

    \I__953\ : InMux
    port map (
            O => \N__4489\,
            I => \N__4483\
        );

    \I__952\ : Span4Mux_h
    port map (
            O => \N__4486\,
            I => \N__4478\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__4483\,
            I => \N__4478\
        );

    \I__950\ : Span4Mux_v
    port map (
            O => \N__4478\,
            I => \N__4475\
        );

    \I__949\ : Sp12to4
    port map (
            O => \N__4475\,
            I => \N__4472\
        );

    \I__948\ : Span12Mux_h
    port map (
            O => \N__4472\,
            I => \N__4469\
        );

    \I__947\ : Odrv12
    port map (
            O => \N__4469\,
            I => \SIZ_c_0\
        );

    \I__946\ : IoInMux
    port map (
            O => \N__4466\,
            I => \N__4462\
        );

    \I__945\ : IoInMux
    port map (
            O => \N__4465\,
            I => \N__4459\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4462\,
            I => \N__4455\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__4459\,
            I => \N__4452\
        );

    \I__942\ : IoInMux
    port map (
            O => \N__4458\,
            I => \N__4449\
        );

    \I__941\ : Span4Mux_s2_h
    port map (
            O => \N__4455\,
            I => \N__4446\
        );

    \I__940\ : IoSpan4Mux
    port map (
            O => \N__4452\,
            I => \N__4443\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__4449\,
            I => \N__4440\
        );

    \I__938\ : Span4Mux_h
    port map (
            O => \N__4446\,
            I => \N__4437\
        );

    \I__937\ : IoSpan4Mux
    port map (
            O => \N__4443\,
            I => \N__4434\
        );

    \I__936\ : Span4Mux_s2_v
    port map (
            O => \N__4440\,
            I => \N__4431\
        );

    \I__935\ : Span4Mux_v
    port map (
            O => \N__4437\,
            I => \N__4428\
        );

    \I__934\ : Span4Mux_s2_v
    port map (
            O => \N__4434\,
            I => \N__4423\
        );

    \I__933\ : Span4Mux_h
    port map (
            O => \N__4431\,
            I => \N__4423\
        );

    \I__932\ : Sp12to4
    port map (
            O => \N__4428\,
            I => \N__4420\
        );

    \I__931\ : Span4Mux_v
    port map (
            O => \N__4423\,
            I => \N__4417\
        );

    \I__930\ : Odrv12
    port map (
            O => \N__4420\,
            I => \CONSTANT_ONE_NET\
        );

    \I__929\ : Odrv4
    port map (
            O => \N__4417\,
            I => \CONSTANT_ONE_NET\
        );

    \I__928\ : InMux
    port map (
            O => \N__4412\,
            I => \N__4409\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__4409\,
            I => \N__4406\
        );

    \I__926\ : Odrv4
    port map (
            O => \N__4406\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\
        );

    \I__925\ : CascadeMux
    port map (
            O => \N__4403\,
            I => \N__4400\
        );

    \I__924\ : InMux
    port map (
            O => \N__4400\,
            I => \N__4397\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__4397\,
            I => \N__4394\
        );

    \I__922\ : Span4Mux_v
    port map (
            O => \N__4394\,
            I => \N__4389\
        );

    \I__921\ : InMux
    port map (
            O => \N__4393\,
            I => \N__4386\
        );

    \I__920\ : InMux
    port map (
            O => \N__4392\,
            I => \N__4383\
        );

    \I__919\ : Sp12to4
    port map (
            O => \N__4389\,
            I => \N__4380\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__4386\,
            I => \N__4375\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__4383\,
            I => \N__4375\
        );

    \I__916\ : Span12Mux_h
    port map (
            O => \N__4380\,
            I => \N__4372\
        );

    \I__915\ : Span12Mux_v
    port map (
            O => \N__4375\,
            I => \N__4369\
        );

    \I__914\ : Span12Mux_v
    port map (
            O => \N__4372\,
            I => \N__4364\
        );

    \I__913\ : Span12Mux_h
    port map (
            O => \N__4369\,
            I => \N__4364\
        );

    \I__912\ : Odrv12
    port map (
            O => \N__4364\,
            I => \D_UU_AMIGA_in_3\
        );

    \I__911\ : IoInMux
    port map (
            O => \N__4361\,
            I => \N__4358\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__4358\,
            I => \N__4355\
        );

    \I__909\ : Span4Mux_s3_v
    port map (
            O => \N__4355\,
            I => \N__4352\
        );

    \I__908\ : Span4Mux_h
    port map (
            O => \N__4352\,
            I => \N__4349\
        );

    \I__907\ : Span4Mux_v
    port map (
            O => \N__4349\,
            I => \N__4346\
        );

    \I__906\ : Sp12to4
    port map (
            O => \N__4346\,
            I => \N__4343\
        );

    \I__905\ : Span12Mux_h
    port map (
            O => \N__4343\,
            I => \N__4340\
        );

    \I__904\ : Odrv12
    port map (
            O => \N__4340\,
            I => \un1_D_UU_AMIGA_3\
        );

    \I__903\ : InMux
    port map (
            O => \N__4337\,
            I => \N__4334\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__4334\,
            I => \N__4331\
        );

    \I__901\ : Span4Mux_v
    port map (
            O => \N__4331\,
            I => \N__4328\
        );

    \I__900\ : Sp12to4
    port map (
            O => \N__4328\,
            I => \N__4325\
        );

    \I__899\ : Span12Mux_h
    port map (
            O => \N__4325\,
            I => \N__4322\
        );

    \I__898\ : Odrv12
    port map (
            O => \N__4322\,
            I => \D_LL_AMIGA_in_5\
        );

    \I__897\ : IoInMux
    port map (
            O => \N__4319\,
            I => \N__4316\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__4316\,
            I => \N__4313\
        );

    \I__895\ : Span4Mux_s2_h
    port map (
            O => \N__4313\,
            I => \N__4310\
        );

    \I__894\ : Span4Mux_v
    port map (
            O => \N__4310\,
            I => \N__4307\
        );

    \I__893\ : Span4Mux_v
    port map (
            O => \N__4307\,
            I => \N__4304\
        );

    \I__892\ : Sp12to4
    port map (
            O => \N__4304\,
            I => \N__4301\
        );

    \I__891\ : Span12Mux_s9_h
    port map (
            O => \N__4301\,
            I => \N__4298\
        );

    \I__890\ : Odrv12
    port map (
            O => \N__4298\,
            I => \un1_D_LL_AMIGA_5\
        );

    \I__889\ : InMux
    port map (
            O => \N__4295\,
            I => \N__4292\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__4292\,
            I => \N__4289\
        );

    \I__887\ : Span12Mux_h
    port map (
            O => \N__4289\,
            I => \N__4286\
        );

    \I__886\ : Odrv12
    port map (
            O => \N__4286\,
            I => \D_LL_AMIGA_in_7\
        );

    \I__885\ : IoInMux
    port map (
            O => \N__4283\,
            I => \N__4280\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__4280\,
            I => \N__4277\
        );

    \I__883\ : Span4Mux_s3_h
    port map (
            O => \N__4277\,
            I => \N__4274\
        );

    \I__882\ : Span4Mux_v
    port map (
            O => \N__4274\,
            I => \N__4271\
        );

    \I__881\ : Sp12to4
    port map (
            O => \N__4271\,
            I => \N__4268\
        );

    \I__880\ : Span12Mux_h
    port map (
            O => \N__4268\,
            I => \N__4265\
        );

    \I__879\ : Odrv12
    port map (
            O => \N__4265\,
            I => \un1_D_LL_AMIGA_7\
        );

    \I__878\ : IoInMux
    port map (
            O => \N__4262\,
            I => \N__4259\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__4259\,
            I => \N__4256\
        );

    \I__876\ : Span12Mux_s5_h
    port map (
            O => \N__4256\,
            I => \N__4253\
        );

    \I__875\ : Span12Mux_h
    port map (
            O => \N__4253\,
            I => \N__4250\
        );

    \I__874\ : Odrv12
    port map (
            O => \N__4250\,
            I => \un1_D_UM_AMIGA_2\
        );

    \I__873\ : SRMux
    port map (
            O => \N__4247\,
            I => \N__4244\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__4244\,
            I => \N__4241\
        );

    \I__871\ : Odrv4
    port map (
            O => \N__4241\,
            I => \U111_CYCLE_SM.RESETn_c_i\
        );

    \I__870\ : InMux
    port map (
            O => \N__4238\,
            I => \N__4234\
        );

    \I__869\ : InMux
    port map (
            O => \N__4237\,
            I => \N__4231\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4234\,
            I => \N__4228\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4231\,
            I => \N__4225\
        );

    \I__866\ : Sp12to4
    port map (
            O => \N__4228\,
            I => \N__4221\
        );

    \I__865\ : Span4Mux_v
    port map (
            O => \N__4225\,
            I => \N__4218\
        );

    \I__864\ : InMux
    port map (
            O => \N__4224\,
            I => \N__4215\
        );

    \I__863\ : Span12Mux_v
    port map (
            O => \N__4221\,
            I => \N__4212\
        );

    \I__862\ : Sp12to4
    port map (
            O => \N__4218\,
            I => \N__4207\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__4215\,
            I => \N__4207\
        );

    \I__860\ : Span12Mux_h
    port map (
            O => \N__4212\,
            I => \N__4204\
        );

    \I__859\ : Span12Mux_h
    port map (
            O => \N__4207\,
            I => \N__4201\
        );

    \I__858\ : Odrv12
    port map (
            O => \N__4204\,
            I => \D_UM_AMIGA_in_2\
        );

    \I__857\ : Odrv12
    port map (
            O => \N__4201\,
            I => \D_UM_AMIGA_in_2\
        );

    \I__856\ : InMux
    port map (
            O => \N__4196\,
            I => \N__4193\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__4193\,
            I => \N__4190\
        );

    \I__854\ : Odrv4
    port map (
            O => \N__4190\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\
        );

    \I__853\ : CascadeMux
    port map (
            O => \N__4187\,
            I => \U111_CYCLE_SM.un3_LW_CYCLE_START_cascade_\
        );

    \I__852\ : CascadeMux
    port map (
            O => \N__4184\,
            I => \N__4181\
        );

    \I__851\ : InMux
    port map (
            O => \N__4181\,
            I => \N__4178\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__4178\,
            I => \N__4175\
        );

    \I__849\ : Span4Mux_h
    port map (
            O => \N__4175\,
            I => \N__4172\
        );

    \I__848\ : Sp12to4
    port map (
            O => \N__4172\,
            I => \N__4169\
        );

    \I__847\ : Odrv12
    port map (
            O => \N__4169\,
            I => \TS_CPUn_c\
        );

    \I__846\ : InMux
    port map (
            O => \N__4166\,
            I => \N__4163\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__4163\,
            I => \N__4160\
        );

    \I__844\ : Span4Mux_v
    port map (
            O => \N__4160\,
            I => \N__4157\
        );

    \I__843\ : Sp12to4
    port map (
            O => \N__4157\,
            I => \N__4154\
        );

    \I__842\ : Span12Mux_h
    port map (
            O => \N__4154\,
            I => \N__4151\
        );

    \I__841\ : Odrv12
    port map (
            O => \N__4151\,
            I => \D_UU_040_in_2\
        );

    \I__840\ : CascadeMux
    port map (
            O => \N__4148\,
            I => \N__4145\
        );

    \I__839\ : InMux
    port map (
            O => \N__4145\,
            I => \N__4141\
        );

    \I__838\ : IoInMux
    port map (
            O => \N__4144\,
            I => \N__4138\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__4141\,
            I => \N__4135\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__4138\,
            I => \N__4132\
        );

    \I__835\ : Sp12to4
    port map (
            O => \N__4135\,
            I => \N__4129\
        );

    \I__834\ : Span12Mux_s9_h
    port map (
            O => \N__4132\,
            I => \N__4126\
        );

    \I__833\ : Span12Mux_v
    port map (
            O => \N__4129\,
            I => \N__4123\
        );

    \I__832\ : Span12Mux_v
    port map (
            O => \N__4126\,
            I => \N__4120\
        );

    \I__831\ : Span12Mux_v
    port map (
            O => \N__4123\,
            I => \N__4117\
        );

    \I__830\ : Span12Mux_h
    port map (
            O => \N__4120\,
            I => \N__4114\
        );

    \I__829\ : Span12Mux_h
    port map (
            O => \N__4117\,
            I => \N__4111\
        );

    \I__828\ : Odrv12
    port map (
            O => \N__4114\,
            I => \D_LM_040_in_2\
        );

    \I__827\ : Odrv12
    port map (
            O => \N__4111\,
            I => \D_LM_040_in_2\
        );

    \I__826\ : IoInMux
    port map (
            O => \N__4106\,
            I => \N__4103\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__4103\,
            I => \N__4100\
        );

    \I__824\ : Span12Mux_s6_v
    port map (
            O => \N__4100\,
            I => \N__4097\
        );

    \I__823\ : Odrv12
    port map (
            O => \N__4097\,
            I => \un1_D_UU_040_2\
        );

    \I__822\ : CascadeMux
    port map (
            O => \N__4094\,
            I => \N__4091\
        );

    \I__821\ : InMux
    port map (
            O => \N__4091\,
            I => \N__4088\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__4088\,
            I => \N__4085\
        );

    \I__819\ : Span4Mux_v
    port map (
            O => \N__4085\,
            I => \N__4082\
        );

    \I__818\ : Span4Mux_h
    port map (
            O => \N__4082\,
            I => \N__4079\
        );

    \I__817\ : Sp12to4
    port map (
            O => \N__4079\,
            I => \N__4076\
        );

    \I__816\ : Span12Mux_h
    port map (
            O => \N__4076\,
            I => \N__4073\
        );

    \I__815\ : Odrv12
    port map (
            O => \N__4073\,
            I => \D_UU_040_in_0\
        );

    \I__814\ : IoInMux
    port map (
            O => \N__4070\,
            I => \N__4067\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__4067\,
            I => \N__4063\
        );

    \I__812\ : InMux
    port map (
            O => \N__4066\,
            I => \N__4060\
        );

    \I__811\ : IoSpan4Mux
    port map (
            O => \N__4063\,
            I => \N__4057\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__4060\,
            I => \N__4054\
        );

    \I__809\ : Span4Mux_s2_h
    port map (
            O => \N__4057\,
            I => \N__4051\
        );

    \I__808\ : Sp12to4
    port map (
            O => \N__4054\,
            I => \N__4048\
        );

    \I__807\ : Span4Mux_v
    port map (
            O => \N__4051\,
            I => \N__4045\
        );

    \I__806\ : Span12Mux_v
    port map (
            O => \N__4048\,
            I => \N__4042\
        );

    \I__805\ : Sp12to4
    port map (
            O => \N__4045\,
            I => \N__4039\
        );

    \I__804\ : Span12Mux_v
    port map (
            O => \N__4042\,
            I => \N__4036\
        );

    \I__803\ : Span12Mux_s9_h
    port map (
            O => \N__4039\,
            I => \N__4033\
        );

    \I__802\ : Span12Mux_h
    port map (
            O => \N__4036\,
            I => \N__4030\
        );

    \I__801\ : Span12Mux_h
    port map (
            O => \N__4033\,
            I => \N__4027\
        );

    \I__800\ : Odrv12
    port map (
            O => \N__4030\,
            I => \D_LM_040_in_0\
        );

    \I__799\ : Odrv12
    port map (
            O => \N__4027\,
            I => \D_LM_040_in_0\
        );

    \I__798\ : IoInMux
    port map (
            O => \N__4022\,
            I => \N__4019\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__4019\,
            I => \N__4016\
        );

    \I__796\ : IoSpan4Mux
    port map (
            O => \N__4016\,
            I => \N__4013\
        );

    \I__795\ : IoSpan4Mux
    port map (
            O => \N__4013\,
            I => \N__4010\
        );

    \I__794\ : Span4Mux_s3_v
    port map (
            O => \N__4010\,
            I => \N__4007\
        );

    \I__793\ : Odrv4
    port map (
            O => \N__4007\,
            I => \un1_D_UU_040_0\
        );

    \I__792\ : IoInMux
    port map (
            O => \N__4004\,
            I => \N__4001\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__4001\,
            I => \N__3997\
        );

    \I__790\ : InMux
    port map (
            O => \N__4000\,
            I => \N__3994\
        );

    \I__789\ : Span4Mux_s2_h
    port map (
            O => \N__3997\,
            I => \N__3991\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__3994\,
            I => \N__3988\
        );

    \I__787\ : Span4Mux_v
    port map (
            O => \N__3991\,
            I => \N__3985\
        );

    \I__786\ : Span12Mux_h
    port map (
            O => \N__3988\,
            I => \N__3982\
        );

    \I__785\ : Sp12to4
    port map (
            O => \N__3985\,
            I => \N__3979\
        );

    \I__784\ : Span12Mux_v
    port map (
            O => \N__3982\,
            I => \N__3976\
        );

    \I__783\ : Span12Mux_h
    port map (
            O => \N__3979\,
            I => \N__3973\
        );

    \I__782\ : Span12Mux_v
    port map (
            O => \N__3976\,
            I => \N__3970\
        );

    \I__781\ : Span12Mux_h
    port map (
            O => \N__3973\,
            I => \N__3967\
        );

    \I__780\ : Odrv12
    port map (
            O => \N__3970\,
            I => \D_LL_040_in_4\
        );

    \I__779\ : Odrv12
    port map (
            O => \N__3967\,
            I => \D_LL_040_in_4\
        );

    \I__778\ : CascadeMux
    port map (
            O => \N__3962\,
            I => \N__3959\
        );

    \I__777\ : InMux
    port map (
            O => \N__3959\,
            I => \N__3956\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__3956\,
            I => \N__3953\
        );

    \I__775\ : Span4Mux_v
    port map (
            O => \N__3953\,
            I => \N__3950\
        );

    \I__774\ : Span4Mux_h
    port map (
            O => \N__3950\,
            I => \N__3947\
        );

    \I__773\ : Sp12to4
    port map (
            O => \N__3947\,
            I => \N__3944\
        );

    \I__772\ : Span12Mux_h
    port map (
            O => \N__3944\,
            I => \N__3941\
        );

    \I__771\ : Odrv12
    port map (
            O => \N__3941\,
            I => \D_UM_040_in_4\
        );

    \I__770\ : IoInMux
    port map (
            O => \N__3938\,
            I => \N__3935\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__3935\,
            I => \N__3932\
        );

    \I__768\ : IoSpan4Mux
    port map (
            O => \N__3932\,
            I => \N__3929\
        );

    \I__767\ : Span4Mux_s2_h
    port map (
            O => \N__3929\,
            I => \N__3926\
        );

    \I__766\ : Span4Mux_h
    port map (
            O => \N__3926\,
            I => \N__3923\
        );

    \I__765\ : Span4Mux_h
    port map (
            O => \N__3923\,
            I => \N__3920\
        );

    \I__764\ : Odrv4
    port map (
            O => \N__3920\,
            I => \un1_D_UM_040_4\
        );

    \I__763\ : InMux
    port map (
            O => \N__3917\,
            I => \N__3914\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__3914\,
            I => \N__3911\
        );

    \I__761\ : Span12Mux_h
    port map (
            O => \N__3911\,
            I => \N__3908\
        );

    \I__760\ : Odrv12
    port map (
            O => \N__3908\,
            I => \D_LM_AMIGA_in_2\
        );

    \I__759\ : IoInMux
    port map (
            O => \N__3905\,
            I => \N__3902\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__3902\,
            I => \N__3899\
        );

    \I__757\ : Span12Mux_s7_h
    port map (
            O => \N__3899\,
            I => \N__3896\
        );

    \I__756\ : Span12Mux_v
    port map (
            O => \N__3896\,
            I => \N__3893\
        );

    \I__755\ : Odrv12
    port map (
            O => \N__3893\,
            I => \un1_D_LM_AMIGA_2\
        );

    \I__754\ : CascadeMux
    port map (
            O => \N__3890\,
            I => \N__3887\
        );

    \I__753\ : InMux
    port map (
            O => \N__3887\,
            I => \N__3884\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__3884\,
            I => \N__3881\
        );

    \I__751\ : Span12Mux_v
    port map (
            O => \N__3881\,
            I => \N__3878\
        );

    \I__750\ : Span12Mux_h
    port map (
            O => \N__3878\,
            I => \N__3875\
        );

    \I__749\ : Odrv12
    port map (
            O => \N__3875\,
            I => \D_LM_AMIGA_in_6\
        );

    \I__748\ : IoInMux
    port map (
            O => \N__3872\,
            I => \N__3869\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__3869\,
            I => \N__3866\
        );

    \I__746\ : IoSpan4Mux
    port map (
            O => \N__3866\,
            I => \N__3863\
        );

    \I__745\ : Sp12to4
    port map (
            O => \N__3863\,
            I => \N__3860\
        );

    \I__744\ : Span12Mux_s9_h
    port map (
            O => \N__3860\,
            I => \N__3857\
        );

    \I__743\ : Odrv12
    port map (
            O => \N__3857\,
            I => \un1_D_LM_AMIGA_6\
        );

    \I__742\ : CascadeMux
    port map (
            O => \N__3854\,
            I => \N__3851\
        );

    \I__741\ : InMux
    port map (
            O => \N__3851\,
            I => \N__3848\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__3848\,
            I => \N__3845\
        );

    \I__739\ : Span4Mux_v
    port map (
            O => \N__3845\,
            I => \N__3842\
        );

    \I__738\ : Sp12to4
    port map (
            O => \N__3842\,
            I => \N__3839\
        );

    \I__737\ : Span12Mux_s2_v
    port map (
            O => \N__3839\,
            I => \N__3836\
        );

    \I__736\ : Span12Mux_h
    port map (
            O => \N__3836\,
            I => \N__3833\
        );

    \I__735\ : Odrv12
    port map (
            O => \N__3833\,
            I => \D_UM_040_in_3\
        );

    \I__734\ : IoInMux
    port map (
            O => \N__3830\,
            I => \N__3827\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__3827\,
            I => \N__3823\
        );

    \I__732\ : InMux
    port map (
            O => \N__3826\,
            I => \N__3820\
        );

    \I__731\ : Span4Mux_s3_h
    port map (
            O => \N__3823\,
            I => \N__3817\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__3820\,
            I => \N__3814\
        );

    \I__729\ : Sp12to4
    port map (
            O => \N__3817\,
            I => \N__3811\
        );

    \I__728\ : Span12Mux_h
    port map (
            O => \N__3814\,
            I => \N__3808\
        );

    \I__727\ : Span12Mux_v
    port map (
            O => \N__3811\,
            I => \N__3805\
        );

    \I__726\ : Span12Mux_v
    port map (
            O => \N__3808\,
            I => \N__3802\
        );

    \I__725\ : Span12Mux_h
    port map (
            O => \N__3805\,
            I => \N__3799\
        );

    \I__724\ : Span12Mux_v
    port map (
            O => \N__3802\,
            I => \N__3796\
        );

    \I__723\ : Span12Mux_h
    port map (
            O => \N__3799\,
            I => \N__3793\
        );

    \I__722\ : Odrv12
    port map (
            O => \N__3796\,
            I => \D_LL_040_in_3\
        );

    \I__721\ : Odrv12
    port map (
            O => \N__3793\,
            I => \D_LL_040_in_3\
        );

    \I__720\ : IoInMux
    port map (
            O => \N__3788\,
            I => \N__3785\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__3785\,
            I => \N__3782\
        );

    \I__718\ : IoSpan4Mux
    port map (
            O => \N__3782\,
            I => \N__3779\
        );

    \I__717\ : Span4Mux_s3_h
    port map (
            O => \N__3779\,
            I => \N__3776\
        );

    \I__716\ : Span4Mux_h
    port map (
            O => \N__3776\,
            I => \N__3773\
        );

    \I__715\ : Span4Mux_h
    port map (
            O => \N__3773\,
            I => \N__3770\
        );

    \I__714\ : Odrv4
    port map (
            O => \N__3770\,
            I => \un1_D_UM_040_3\
        );

    \I__713\ : CascadeMux
    port map (
            O => \N__3767\,
            I => \N__3764\
        );

    \I__712\ : InMux
    port map (
            O => \N__3764\,
            I => \N__3761\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__3761\,
            I => \N__3758\
        );

    \I__710\ : Span4Mux_h
    port map (
            O => \N__3758\,
            I => \N__3755\
        );

    \I__709\ : Sp12to4
    port map (
            O => \N__3755\,
            I => \N__3752\
        );

    \I__708\ : Span12Mux_v
    port map (
            O => \N__3752\,
            I => \N__3749\
        );

    \I__707\ : Span12Mux_h
    port map (
            O => \N__3749\,
            I => \N__3746\
        );

    \I__706\ : Odrv12
    port map (
            O => \N__3746\,
            I => \D_UU_040_in_5\
        );

    \I__705\ : IoInMux
    port map (
            O => \N__3743\,
            I => \N__3740\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__3740\,
            I => \N__3737\
        );

    \I__703\ : IoSpan4Mux
    port map (
            O => \N__3737\,
            I => \N__3734\
        );

    \I__702\ : Span4Mux_s0_h
    port map (
            O => \N__3734\,
            I => \N__3731\
        );

    \I__701\ : Span4Mux_v
    port map (
            O => \N__3731\,
            I => \N__3727\
        );

    \I__700\ : InMux
    port map (
            O => \N__3730\,
            I => \N__3724\
        );

    \I__699\ : Sp12to4
    port map (
            O => \N__3727\,
            I => \N__3721\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__3724\,
            I => \N__3718\
        );

    \I__697\ : Span12Mux_h
    port map (
            O => \N__3721\,
            I => \N__3713\
        );

    \I__696\ : Span12Mux_v
    port map (
            O => \N__3718\,
            I => \N__3713\
        );

    \I__695\ : Span12Mux_h
    port map (
            O => \N__3713\,
            I => \N__3710\
        );

    \I__694\ : Odrv12
    port map (
            O => \N__3710\,
            I => \D_LM_040_in_5\
        );

    \I__693\ : IoInMux
    port map (
            O => \N__3707\,
            I => \N__3704\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__3704\,
            I => \N__3701\
        );

    \I__691\ : Span4Mux_s2_h
    port map (
            O => \N__3701\,
            I => \N__3698\
        );

    \I__690\ : Span4Mux_h
    port map (
            O => \N__3698\,
            I => \N__3695\
        );

    \I__689\ : Sp12to4
    port map (
            O => \N__3695\,
            I => \N__3692\
        );

    \I__688\ : Span12Mux_s7_v
    port map (
            O => \N__3692\,
            I => \N__3689\
        );

    \I__687\ : Odrv12
    port map (
            O => \N__3689\,
            I => \un1_D_UU_040_5\
        );

    \I__686\ : CascadeMux
    port map (
            O => \N__3686\,
            I => \N__3683\
        );

    \I__685\ : InMux
    port map (
            O => \N__3683\,
            I => \N__3680\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__3680\,
            I => \N__3677\
        );

    \I__683\ : Span4Mux_v
    port map (
            O => \N__3677\,
            I => \N__3674\
        );

    \I__682\ : Span4Mux_h
    port map (
            O => \N__3674\,
            I => \N__3671\
        );

    \I__681\ : Sp12to4
    port map (
            O => \N__3671\,
            I => \N__3668\
        );

    \I__680\ : Span12Mux_h
    port map (
            O => \N__3668\,
            I => \N__3665\
        );

    \I__679\ : Odrv12
    port map (
            O => \N__3665\,
            I => \D_UM_040_in_5\
        );

    \I__678\ : IoInMux
    port map (
            O => \N__3662\,
            I => \N__3658\
        );

    \I__677\ : InMux
    port map (
            O => \N__3661\,
            I => \N__3655\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__3658\,
            I => \N__3652\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__3655\,
            I => \N__3649\
        );

    \I__674\ : IoSpan4Mux
    port map (
            O => \N__3652\,
            I => \N__3646\
        );

    \I__673\ : Span4Mux_v
    port map (
            O => \N__3649\,
            I => \N__3643\
        );

    \I__672\ : Span4Mux_s3_h
    port map (
            O => \N__3646\,
            I => \N__3640\
        );

    \I__671\ : Sp12to4
    port map (
            O => \N__3643\,
            I => \N__3637\
        );

    \I__670\ : Sp12to4
    port map (
            O => \N__3640\,
            I => \N__3634\
        );

    \I__669\ : Span12Mux_h
    port map (
            O => \N__3637\,
            I => \N__3631\
        );

    \I__668\ : Span12Mux_v
    port map (
            O => \N__3634\,
            I => \N__3628\
        );

    \I__667\ : Span12Mux_v
    port map (
            O => \N__3631\,
            I => \N__3625\
        );

    \I__666\ : Span12Mux_h
    port map (
            O => \N__3628\,
            I => \N__3622\
        );

    \I__665\ : Span12Mux_v
    port map (
            O => \N__3625\,
            I => \N__3617\
        );

    \I__664\ : Span12Mux_h
    port map (
            O => \N__3622\,
            I => \N__3617\
        );

    \I__663\ : Odrv12
    port map (
            O => \N__3617\,
            I => \D_LL_040_in_5\
        );

    \I__662\ : IoInMux
    port map (
            O => \N__3614\,
            I => \N__3611\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__3611\,
            I => \N__3608\
        );

    \I__660\ : IoSpan4Mux
    port map (
            O => \N__3608\,
            I => \N__3605\
        );

    \I__659\ : Sp12to4
    port map (
            O => \N__3605\,
            I => \N__3602\
        );

    \I__658\ : Span12Mux_s6_v
    port map (
            O => \N__3602\,
            I => \N__3599\
        );

    \I__657\ : Odrv12
    port map (
            O => \N__3599\,
            I => \un1_D_UM_040_5\
        );

    \I__656\ : CascadeMux
    port map (
            O => \N__3596\,
            I => \N__3593\
        );

    \I__655\ : InMux
    port map (
            O => \N__3593\,
            I => \N__3590\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__3590\,
            I => \N__3587\
        );

    \I__653\ : Span4Mux_v
    port map (
            O => \N__3587\,
            I => \N__3584\
        );

    \I__652\ : Sp12to4
    port map (
            O => \N__3584\,
            I => \N__3581\
        );

    \I__651\ : Odrv12
    port map (
            O => \N__3581\,
            I => \D_LL_AMIGA_in_6\
        );

    \I__650\ : IoInMux
    port map (
            O => \N__3578\,
            I => \N__3575\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__3575\,
            I => \N__3572\
        );

    \I__648\ : Span4Mux_s2_h
    port map (
            O => \N__3572\,
            I => \N__3569\
        );

    \I__647\ : Span4Mux_v
    port map (
            O => \N__3569\,
            I => \N__3566\
        );

    \I__646\ : Span4Mux_v
    port map (
            O => \N__3566\,
            I => \N__3563\
        );

    \I__645\ : Sp12to4
    port map (
            O => \N__3563\,
            I => \N__3560\
        );

    \I__644\ : Span12Mux_s11_h
    port map (
            O => \N__3560\,
            I => \N__3557\
        );

    \I__643\ : Odrv12
    port map (
            O => \N__3557\,
            I => \un1_D_LL_AMIGA_6\
        );

    \I__642\ : InMux
    port map (
            O => \N__3554\,
            I => \N__3551\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__3551\,
            I => \N__3548\
        );

    \I__640\ : Span4Mux_v
    port map (
            O => \N__3548\,
            I => \N__3545\
        );

    \I__639\ : Sp12to4
    port map (
            O => \N__3545\,
            I => \N__3542\
        );

    \I__638\ : Odrv12
    port map (
            O => \N__3542\,
            I => \D_LM_AMIGA_in_5\
        );

    \I__637\ : IoInMux
    port map (
            O => \N__3539\,
            I => \N__3536\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__3536\,
            I => \N__3533\
        );

    \I__635\ : IoSpan4Mux
    port map (
            O => \N__3533\,
            I => \N__3530\
        );

    \I__634\ : Sp12to4
    port map (
            O => \N__3530\,
            I => \N__3527\
        );

    \I__633\ : Span12Mux_s9_h
    port map (
            O => \N__3527\,
            I => \N__3524\
        );

    \I__632\ : Span12Mux_h
    port map (
            O => \N__3524\,
            I => \N__3521\
        );

    \I__631\ : Odrv12
    port map (
            O => \N__3521\,
            I => \un1_D_LM_AMIGA_5\
        );

    \I__630\ : CascadeMux
    port map (
            O => \N__3518\,
            I => \N__3515\
        );

    \I__629\ : InMux
    port map (
            O => \N__3515\,
            I => \N__3512\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__3512\,
            I => \N__3509\
        );

    \I__627\ : Span4Mux_v
    port map (
            O => \N__3509\,
            I => \N__3506\
        );

    \I__626\ : Sp12to4
    port map (
            O => \N__3506\,
            I => \N__3503\
        );

    \I__625\ : Odrv12
    port map (
            O => \N__3503\,
            I => \D_LM_AMIGA_in_7\
        );

    \I__624\ : IoInMux
    port map (
            O => \N__3500\,
            I => \N__3497\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3497\,
            I => \N__3494\
        );

    \I__622\ : Span12Mux_s4_h
    port map (
            O => \N__3494\,
            I => \N__3491\
        );

    \I__621\ : Span12Mux_h
    port map (
            O => \N__3491\,
            I => \N__3488\
        );

    \I__620\ : Odrv12
    port map (
            O => \N__3488\,
            I => \un1_D_LM_AMIGA_7\
        );

    \I__619\ : IoInMux
    port map (
            O => \N__3485\,
            I => \N__3482\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__3482\,
            I => \N__3479\
        );

    \I__617\ : Odrv12
    port map (
            O => \N__3479\,
            I => \TSn_c\
        );

    \I__616\ : InMux
    port map (
            O => \N__3476\,
            I => \N__3473\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__3473\,
            I => \N__3470\
        );

    \I__614\ : Span4Mux_v
    port map (
            O => \N__3470\,
            I => \N__3467\
        );

    \I__613\ : Span4Mux_h
    port map (
            O => \N__3467\,
            I => \N__3464\
        );

    \I__612\ : Span4Mux_h
    port map (
            O => \N__3464\,
            I => \N__3461\
        );

    \I__611\ : Odrv4
    port map (
            O => \N__3461\,
            I => \D_LL_AMIGA_in_0\
        );

    \I__610\ : IoInMux
    port map (
            O => \N__3458\,
            I => \N__3455\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__3455\,
            I => \N__3452\
        );

    \I__608\ : IoSpan4Mux
    port map (
            O => \N__3452\,
            I => \N__3449\
        );

    \I__607\ : IoSpan4Mux
    port map (
            O => \N__3449\,
            I => \N__3446\
        );

    \I__606\ : Sp12to4
    port map (
            O => \N__3446\,
            I => \N__3443\
        );

    \I__605\ : Span12Mux_s9_h
    port map (
            O => \N__3443\,
            I => \N__3440\
        );

    \I__604\ : Odrv12
    port map (
            O => \N__3440\,
            I => \un1_D_LL_AMIGA_0\
        );

    \I__603\ : InMux
    port map (
            O => \N__3437\,
            I => \N__3434\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__3434\,
            I => \N__3431\
        );

    \I__601\ : Span4Mux_v
    port map (
            O => \N__3431\,
            I => \N__3428\
        );

    \I__600\ : Sp12to4
    port map (
            O => \N__3428\,
            I => \N__3425\
        );

    \I__599\ : Span12Mux_h
    port map (
            O => \N__3425\,
            I => \N__3422\
        );

    \I__598\ : Odrv12
    port map (
            O => \N__3422\,
            I => \D_UU_040_in_4\
        );

    \I__597\ : IoInMux
    port map (
            O => \N__3419\,
            I => \N__3416\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3416\,
            I => \N__3413\
        );

    \I__595\ : Span4Mux_s1_h
    port map (
            O => \N__3413\,
            I => \N__3409\
        );

    \I__594\ : InMux
    port map (
            O => \N__3412\,
            I => \N__3406\
        );

    \I__593\ : Sp12to4
    port map (
            O => \N__3409\,
            I => \N__3403\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__3406\,
            I => \N__3400\
        );

    \I__591\ : Span12Mux_v
    port map (
            O => \N__3403\,
            I => \N__3397\
        );

    \I__590\ : Span12Mux_h
    port map (
            O => \N__3400\,
            I => \N__3394\
        );

    \I__589\ : Span12Mux_h
    port map (
            O => \N__3397\,
            I => \N__3391\
        );

    \I__588\ : Span12Mux_v
    port map (
            O => \N__3394\,
            I => \N__3388\
        );

    \I__587\ : Span12Mux_h
    port map (
            O => \N__3391\,
            I => \N__3385\
        );

    \I__586\ : Span12Mux_h
    port map (
            O => \N__3388\,
            I => \N__3382\
        );

    \I__585\ : Odrv12
    port map (
            O => \N__3385\,
            I => \D_LM_040_in_4\
        );

    \I__584\ : Odrv12
    port map (
            O => \N__3382\,
            I => \D_LM_040_in_4\
        );

    \I__583\ : IoInMux
    port map (
            O => \N__3377\,
            I => \N__3374\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__3374\,
            I => \N__3371\
        );

    \I__581\ : Span4Mux_s2_v
    port map (
            O => \N__3371\,
            I => \N__3368\
        );

    \I__580\ : Span4Mux_h
    port map (
            O => \N__3368\,
            I => \N__3365\
        );

    \I__579\ : Span4Mux_v
    port map (
            O => \N__3365\,
            I => \N__3362\
        );

    \I__578\ : Odrv4
    port map (
            O => \N__3362\,
            I => \un1_D_UU_040_4\
        );

    \I__577\ : InMux
    port map (
            O => \N__3359\,
            I => \N__3356\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__3356\,
            I => \N__3353\
        );

    \I__575\ : Span4Mux_v
    port map (
            O => \N__3353\,
            I => \N__3350\
        );

    \I__574\ : Sp12to4
    port map (
            O => \N__3350\,
            I => \N__3347\
        );

    \I__573\ : Span12Mux_h
    port map (
            O => \N__3347\,
            I => \N__3344\
        );

    \I__572\ : Odrv12
    port map (
            O => \N__3344\,
            I => \D_LL_AMIGA_in_1\
        );

    \I__571\ : IoInMux
    port map (
            O => \N__3341\,
            I => \N__3338\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3338\,
            I => \N__3335\
        );

    \I__569\ : IoSpan4Mux
    port map (
            O => \N__3335\,
            I => \N__3332\
        );

    \I__568\ : IoSpan4Mux
    port map (
            O => \N__3332\,
            I => \N__3329\
        );

    \I__567\ : Span4Mux_s2_h
    port map (
            O => \N__3329\,
            I => \N__3326\
        );

    \I__566\ : Sp12to4
    port map (
            O => \N__3326\,
            I => \N__3323\
        );

    \I__565\ : Span12Mux_s11_h
    port map (
            O => \N__3323\,
            I => \N__3320\
        );

    \I__564\ : Odrv12
    port map (
            O => \N__3320\,
            I => \un1_D_LL_AMIGA_1\
        );

    \I__563\ : InMux
    port map (
            O => \N__3317\,
            I => \N__3314\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3314\,
            I => \N__3311\
        );

    \I__561\ : Span4Mux_v
    port map (
            O => \N__3311\,
            I => \N__3308\
        );

    \I__560\ : Sp12to4
    port map (
            O => \N__3308\,
            I => \N__3305\
        );

    \I__559\ : Span12Mux_h
    port map (
            O => \N__3305\,
            I => \N__3302\
        );

    \I__558\ : Odrv12
    port map (
            O => \N__3302\,
            I => \D_LL_AMIGA_in_2\
        );

    \I__557\ : IoInMux
    port map (
            O => \N__3299\,
            I => \N__3296\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__3296\,
            I => \N__3293\
        );

    \I__555\ : IoSpan4Mux
    port map (
            O => \N__3293\,
            I => \N__3290\
        );

    \I__554\ : Sp12to4
    port map (
            O => \N__3290\,
            I => \N__3287\
        );

    \I__553\ : Span12Mux_s7_h
    port map (
            O => \N__3287\,
            I => \N__3284\
        );

    \I__552\ : Span12Mux_h
    port map (
            O => \N__3284\,
            I => \N__3281\
        );

    \I__551\ : Odrv12
    port map (
            O => \N__3281\,
            I => \un1_D_LL_AMIGA_2\
        );

    \I__550\ : InMux
    port map (
            O => \N__3278\,
            I => \N__3275\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3275\,
            I => \N__3272\
        );

    \I__548\ : Span4Mux_v
    port map (
            O => \N__3272\,
            I => \N__3269\
        );

    \I__547\ : Sp12to4
    port map (
            O => \N__3269\,
            I => \N__3266\
        );

    \I__546\ : Span12Mux_h
    port map (
            O => \N__3266\,
            I => \N__3263\
        );

    \I__545\ : Odrv12
    port map (
            O => \N__3263\,
            I => \D_LM_AMIGA_in_0\
        );

    \I__544\ : IoInMux
    port map (
            O => \N__3260\,
            I => \N__3257\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__3257\,
            I => \N__3254\
        );

    \I__542\ : Span12Mux_s7_h
    port map (
            O => \N__3254\,
            I => \N__3251\
        );

    \I__541\ : Span12Mux_h
    port map (
            O => \N__3251\,
            I => \N__3248\
        );

    \I__540\ : Odrv12
    port map (
            O => \N__3248\,
            I => \un1_D_LM_AMIGA_0\
        );

    \I__539\ : CascadeMux
    port map (
            O => \N__3245\,
            I => \N__3242\
        );

    \I__538\ : InMux
    port map (
            O => \N__3242\,
            I => \N__3239\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__3239\,
            I => \N__3236\
        );

    \I__536\ : Span12Mux_h
    port map (
            O => \N__3236\,
            I => \N__3233\
        );

    \I__535\ : Span12Mux_h
    port map (
            O => \N__3233\,
            I => \N__3230\
        );

    \I__534\ : Odrv12
    port map (
            O => \N__3230\,
            I => \D_UM_040_in_2\
        );

    \I__533\ : InMux
    port map (
            O => \N__3227\,
            I => \N__3223\
        );

    \I__532\ : IoInMux
    port map (
            O => \N__3226\,
            I => \N__3220\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__3223\,
            I => \N__3217\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__3220\,
            I => \N__3214\
        );

    \I__529\ : Span4Mux_v
    port map (
            O => \N__3217\,
            I => \N__3211\
        );

    \I__528\ : Span4Mux_s1_h
    port map (
            O => \N__3214\,
            I => \N__3208\
        );

    \I__527\ : Sp12to4
    port map (
            O => \N__3211\,
            I => \N__3205\
        );

    \I__526\ : Sp12to4
    port map (
            O => \N__3208\,
            I => \N__3202\
        );

    \I__525\ : Span12Mux_h
    port map (
            O => \N__3205\,
            I => \N__3199\
        );

    \I__524\ : Span12Mux_v
    port map (
            O => \N__3202\,
            I => \N__3196\
        );

    \I__523\ : Span12Mux_v
    port map (
            O => \N__3199\,
            I => \N__3193\
        );

    \I__522\ : Span12Mux_h
    port map (
            O => \N__3196\,
            I => \N__3190\
        );

    \I__521\ : Span12Mux_h
    port map (
            O => \N__3193\,
            I => \N__3187\
        );

    \I__520\ : Span12Mux_h
    port map (
            O => \N__3190\,
            I => \N__3184\
        );

    \I__519\ : Odrv12
    port map (
            O => \N__3187\,
            I => \D_LL_040_in_2\
        );

    \I__518\ : Odrv12
    port map (
            O => \N__3184\,
            I => \D_LL_040_in_2\
        );

    \I__517\ : IoInMux
    port map (
            O => \N__3179\,
            I => \N__3176\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__3176\,
            I => \N__3173\
        );

    \I__515\ : Span4Mux_s3_h
    port map (
            O => \N__3173\,
            I => \N__3170\
        );

    \I__514\ : Span4Mux_v
    port map (
            O => \N__3170\,
            I => \N__3167\
        );

    \I__513\ : Odrv4
    port map (
            O => \N__3167\,
            I => \un1_D_UM_040_2\
        );

    \I__512\ : InMux
    port map (
            O => \N__3164\,
            I => \N__3160\
        );

    \I__511\ : IoInMux
    port map (
            O => \N__3163\,
            I => \N__3157\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__3160\,
            I => \N__3154\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__3157\,
            I => \N__3151\
        );

    \I__508\ : Sp12to4
    port map (
            O => \N__3154\,
            I => \N__3148\
        );

    \I__507\ : Span4Mux_s3_h
    port map (
            O => \N__3151\,
            I => \N__3145\
        );

    \I__506\ : Span12Mux_v
    port map (
            O => \N__3148\,
            I => \N__3142\
        );

    \I__505\ : Sp12to4
    port map (
            O => \N__3145\,
            I => \N__3139\
        );

    \I__504\ : Span12Mux_v
    port map (
            O => \N__3142\,
            I => \N__3136\
        );

    \I__503\ : Span12Mux_v
    port map (
            O => \N__3139\,
            I => \N__3133\
        );

    \I__502\ : Span12Mux_h
    port map (
            O => \N__3136\,
            I => \N__3130\
        );

    \I__501\ : Span12Mux_h
    port map (
            O => \N__3133\,
            I => \N__3127\
        );

    \I__500\ : Span12Mux_h
    port map (
            O => \N__3130\,
            I => \N__3124\
        );

    \I__499\ : Span12Mux_h
    port map (
            O => \N__3127\,
            I => \N__3121\
        );

    \I__498\ : Odrv12
    port map (
            O => \N__3124\,
            I => \D_LL_040_in_1\
        );

    \I__497\ : Odrv12
    port map (
            O => \N__3121\,
            I => \D_LL_040_in_1\
        );

    \I__496\ : CascadeMux
    port map (
            O => \N__3116\,
            I => \N__3113\
        );

    \I__495\ : InMux
    port map (
            O => \N__3113\,
            I => \N__3110\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__3110\,
            I => \N__3107\
        );

    \I__493\ : Span4Mux_h
    port map (
            O => \N__3107\,
            I => \N__3104\
        );

    \I__492\ : Sp12to4
    port map (
            O => \N__3104\,
            I => \N__3101\
        );

    \I__491\ : Span12Mux_v
    port map (
            O => \N__3101\,
            I => \N__3098\
        );

    \I__490\ : Span12Mux_h
    port map (
            O => \N__3098\,
            I => \N__3095\
        );

    \I__489\ : Odrv12
    port map (
            O => \N__3095\,
            I => \D_UM_040_in_1\
        );

    \I__488\ : IoInMux
    port map (
            O => \N__3092\,
            I => \N__3089\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__3089\,
            I => \N__3086\
        );

    \I__486\ : Span4Mux_s2_h
    port map (
            O => \N__3086\,
            I => \N__3083\
        );

    \I__485\ : Span4Mux_h
    port map (
            O => \N__3083\,
            I => \N__3080\
        );

    \I__484\ : Odrv4
    port map (
            O => \N__3080\,
            I => \un1_D_UM_040_1\
        );

    \I__483\ : IoInMux
    port map (
            O => \N__3077\,
            I => \N__3073\
        );

    \I__482\ : InMux
    port map (
            O => \N__3076\,
            I => \N__3070\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__3073\,
            I => \N__3067\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3070\,
            I => \N__3064\
        );

    \I__479\ : IoSpan4Mux
    port map (
            O => \N__3067\,
            I => \N__3061\
        );

    \I__478\ : Sp12to4
    port map (
            O => \N__3064\,
            I => \N__3058\
        );

    \I__477\ : Span4Mux_s3_h
    port map (
            O => \N__3061\,
            I => \N__3055\
        );

    \I__476\ : Span12Mux_v
    port map (
            O => \N__3058\,
            I => \N__3052\
        );

    \I__475\ : Sp12to4
    port map (
            O => \N__3055\,
            I => \N__3049\
        );

    \I__474\ : Span12Mux_v
    port map (
            O => \N__3052\,
            I => \N__3046\
        );

    \I__473\ : Span12Mux_v
    port map (
            O => \N__3049\,
            I => \N__3043\
        );

    \I__472\ : Span12Mux_h
    port map (
            O => \N__3046\,
            I => \N__3040\
        );

    \I__471\ : Span12Mux_h
    port map (
            O => \N__3043\,
            I => \N__3037\
        );

    \I__470\ : Span12Mux_h
    port map (
            O => \N__3040\,
            I => \N__3034\
        );

    \I__469\ : Span12Mux_h
    port map (
            O => \N__3037\,
            I => \N__3031\
        );

    \I__468\ : Odrv12
    port map (
            O => \N__3034\,
            I => \D_LL_040_in_7\
        );

    \I__467\ : Odrv12
    port map (
            O => \N__3031\,
            I => \D_LL_040_in_7\
        );

    \I__466\ : CascadeMux
    port map (
            O => \N__3026\,
            I => \N__3023\
        );

    \I__465\ : InMux
    port map (
            O => \N__3023\,
            I => \N__3020\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__3020\,
            I => \N__3017\
        );

    \I__463\ : Span4Mux_v
    port map (
            O => \N__3017\,
            I => \N__3014\
        );

    \I__462\ : Span4Mux_v
    port map (
            O => \N__3014\,
            I => \N__3011\
        );

    \I__461\ : Sp12to4
    port map (
            O => \N__3011\,
            I => \N__3008\
        );

    \I__460\ : Span12Mux_h
    port map (
            O => \N__3008\,
            I => \N__3005\
        );

    \I__459\ : Span12Mux_h
    port map (
            O => \N__3005\,
            I => \N__3002\
        );

    \I__458\ : Odrv12
    port map (
            O => \N__3002\,
            I => \D_UM_040_in_7\
        );

    \I__457\ : IoInMux
    port map (
            O => \N__2999\,
            I => \N__2996\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__2996\,
            I => \N__2993\
        );

    \I__455\ : Span4Mux_s1_h
    port map (
            O => \N__2993\,
            I => \N__2990\
        );

    \I__454\ : Span4Mux_h
    port map (
            O => \N__2990\,
            I => \N__2987\
        );

    \I__453\ : Span4Mux_v
    port map (
            O => \N__2987\,
            I => \N__2984\
        );

    \I__452\ : Odrv4
    port map (
            O => \N__2984\,
            I => \un1_D_UM_040_7\
        );

    \I__451\ : InMux
    port map (
            O => \N__2981\,
            I => \N__2978\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__2978\,
            I => \N__2975\
        );

    \I__449\ : Sp12to4
    port map (
            O => \N__2975\,
            I => \N__2972\
        );

    \I__448\ : Span12Mux_v
    port map (
            O => \N__2972\,
            I => \N__2969\
        );

    \I__447\ : Span12Mux_h
    port map (
            O => \N__2969\,
            I => \N__2966\
        );

    \I__446\ : Span12Mux_h
    port map (
            O => \N__2966\,
            I => \N__2963\
        );

    \I__445\ : Odrv12
    port map (
            O => \N__2963\,
            I => \D_UU_040_in_1\
        );

    \I__444\ : CascadeMux
    port map (
            O => \N__2960\,
            I => \N__2957\
        );

    \I__443\ : InMux
    port map (
            O => \N__2957\,
            I => \N__2953\
        );

    \I__442\ : IoInMux
    port map (
            O => \N__2956\,
            I => \N__2950\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__2953\,
            I => \N__2947\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__2950\,
            I => \N__2944\
        );

    \I__439\ : Sp12to4
    port map (
            O => \N__2947\,
            I => \N__2941\
        );

    \I__438\ : Span4Mux_s3_h
    port map (
            O => \N__2944\,
            I => \N__2938\
        );

    \I__437\ : Span12Mux_v
    port map (
            O => \N__2941\,
            I => \N__2935\
        );

    \I__436\ : Sp12to4
    port map (
            O => \N__2938\,
            I => \N__2932\
        );

    \I__435\ : Span12Mux_v
    port map (
            O => \N__2935\,
            I => \N__2929\
        );

    \I__434\ : Span12Mux_v
    port map (
            O => \N__2932\,
            I => \N__2926\
        );

    \I__433\ : Span12Mux_h
    port map (
            O => \N__2929\,
            I => \N__2923\
        );

    \I__432\ : Span12Mux_h
    port map (
            O => \N__2926\,
            I => \N__2920\
        );

    \I__431\ : Span12Mux_h
    port map (
            O => \N__2923\,
            I => \N__2917\
        );

    \I__430\ : Span12Mux_h
    port map (
            O => \N__2920\,
            I => \N__2914\
        );

    \I__429\ : Odrv12
    port map (
            O => \N__2917\,
            I => \D_LM_040_in_1\
        );

    \I__428\ : Odrv12
    port map (
            O => \N__2914\,
            I => \D_LM_040_in_1\
        );

    \I__427\ : IoInMux
    port map (
            O => \N__2909\,
            I => \N__2906\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__2906\,
            I => \N__2903\
        );

    \I__425\ : Span4Mux_s2_h
    port map (
            O => \N__2903\,
            I => \N__2900\
        );

    \I__424\ : Span4Mux_h
    port map (
            O => \N__2900\,
            I => \N__2897\
        );

    \I__423\ : Odrv4
    port map (
            O => \N__2897\,
            I => \un1_D_UU_040_1\
        );

    \I__422\ : InMux
    port map (
            O => \N__2894\,
            I => \N__2891\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__2891\,
            I => \N__2888\
        );

    \I__420\ : Odrv12
    port map (
            O => \N__2888\,
            I => \D_LM_AMIGA_in_3\
        );

    \I__419\ : IoInMux
    port map (
            O => \N__2885\,
            I => \N__2882\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__2882\,
            I => \N__2879\
        );

    \I__417\ : Span4Mux_s2_h
    port map (
            O => \N__2879\,
            I => \N__2876\
        );

    \I__416\ : Sp12to4
    port map (
            O => \N__2876\,
            I => \N__2873\
        );

    \I__415\ : Span12Mux_v
    port map (
            O => \N__2873\,
            I => \N__2870\
        );

    \I__414\ : Span12Mux_h
    port map (
            O => \N__2870\,
            I => \N__2867\
        );

    \I__413\ : Odrv12
    port map (
            O => \N__2867\,
            I => \un1_D_LM_AMIGA_3\
        );

    \I__412\ : IoInMux
    port map (
            O => \N__2864\,
            I => \N__2861\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__2861\,
            I => \N__2858\
        );

    \I__410\ : IoSpan4Mux
    port map (
            O => \N__2858\,
            I => \N__2854\
        );

    \I__409\ : InMux
    port map (
            O => \N__2857\,
            I => \N__2851\
        );

    \I__408\ : Span4Mux_s2_h
    port map (
            O => \N__2854\,
            I => \N__2848\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__2851\,
            I => \N__2845\
        );

    \I__406\ : Sp12to4
    port map (
            O => \N__2848\,
            I => \N__2842\
        );

    \I__405\ : Span4Mux_v
    port map (
            O => \N__2845\,
            I => \N__2839\
        );

    \I__404\ : Span12Mux_h
    port map (
            O => \N__2842\,
            I => \N__2836\
        );

    \I__403\ : Sp12to4
    port map (
            O => \N__2839\,
            I => \N__2833\
        );

    \I__402\ : Span12Mux_h
    port map (
            O => \N__2836\,
            I => \N__2830\
        );

    \I__401\ : Span12Mux_h
    port map (
            O => \N__2833\,
            I => \N__2827\
        );

    \I__400\ : Odrv12
    port map (
            O => \N__2830\,
            I => \D_LM_040_in_7\
        );

    \I__399\ : Odrv12
    port map (
            O => \N__2827\,
            I => \D_LM_040_in_7\
        );

    \I__398\ : CascadeMux
    port map (
            O => \N__2822\,
            I => \N__2819\
        );

    \I__397\ : InMux
    port map (
            O => \N__2819\,
            I => \N__2816\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__2816\,
            I => \N__2813\
        );

    \I__395\ : Span4Mux_v
    port map (
            O => \N__2813\,
            I => \N__2810\
        );

    \I__394\ : Sp12to4
    port map (
            O => \N__2810\,
            I => \N__2807\
        );

    \I__393\ : Span12Mux_h
    port map (
            O => \N__2807\,
            I => \N__2804\
        );

    \I__392\ : Span12Mux_h
    port map (
            O => \N__2804\,
            I => \N__2801\
        );

    \I__391\ : Odrv12
    port map (
            O => \N__2801\,
            I => \D_UU_040_in_7\
        );

    \I__390\ : IoInMux
    port map (
            O => \N__2798\,
            I => \N__2795\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__2795\,
            I => \N__2792\
        );

    \I__388\ : Span4Mux_s2_v
    port map (
            O => \N__2792\,
            I => \N__2789\
        );

    \I__387\ : Span4Mux_h
    port map (
            O => \N__2789\,
            I => \N__2786\
        );

    \I__386\ : Span4Mux_v
    port map (
            O => \N__2786\,
            I => \N__2783\
        );

    \I__385\ : Odrv4
    port map (
            O => \N__2783\,
            I => \un1_D_UU_040_7\
        );

    \I__384\ : IoInMux
    port map (
            O => \N__2780\,
            I => \N__2777\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__2777\,
            I => \N__2773\
        );

    \I__382\ : InMux
    port map (
            O => \N__2776\,
            I => \N__2770\
        );

    \I__381\ : IoSpan4Mux
    port map (
            O => \N__2773\,
            I => \N__2767\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__2770\,
            I => \N__2764\
        );

    \I__379\ : IoSpan4Mux
    port map (
            O => \N__2767\,
            I => \N__2761\
        );

    \I__378\ : Span4Mux_v
    port map (
            O => \N__2764\,
            I => \N__2758\
        );

    \I__377\ : Span4Mux_s2_h
    port map (
            O => \N__2761\,
            I => \N__2755\
        );

    \I__376\ : Sp12to4
    port map (
            O => \N__2758\,
            I => \N__2752\
        );

    \I__375\ : Sp12to4
    port map (
            O => \N__2755\,
            I => \N__2749\
        );

    \I__374\ : Span12Mux_v
    port map (
            O => \N__2752\,
            I => \N__2746\
        );

    \I__373\ : Span12Mux_h
    port map (
            O => \N__2749\,
            I => \N__2743\
        );

    \I__372\ : Span12Mux_h
    port map (
            O => \N__2746\,
            I => \N__2740\
        );

    \I__371\ : Span12Mux_h
    port map (
            O => \N__2743\,
            I => \N__2737\
        );

    \I__370\ : Odrv12
    port map (
            O => \N__2740\,
            I => \D_LM_040_in_3\
        );

    \I__369\ : Odrv12
    port map (
            O => \N__2737\,
            I => \D_LM_040_in_3\
        );

    \I__368\ : CascadeMux
    port map (
            O => \N__2732\,
            I => \N__2729\
        );

    \I__367\ : InMux
    port map (
            O => \N__2729\,
            I => \N__2726\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__2726\,
            I => \N__2723\
        );

    \I__365\ : Span4Mux_v
    port map (
            O => \N__2723\,
            I => \N__2720\
        );

    \I__364\ : Sp12to4
    port map (
            O => \N__2720\,
            I => \N__2717\
        );

    \I__363\ : Span12Mux_h
    port map (
            O => \N__2717\,
            I => \N__2714\
        );

    \I__362\ : Span12Mux_h
    port map (
            O => \N__2714\,
            I => \N__2711\
        );

    \I__361\ : Odrv12
    port map (
            O => \N__2711\,
            I => \D_UU_040_in_3\
        );

    \I__360\ : IoInMux
    port map (
            O => \N__2708\,
            I => \N__2705\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__2705\,
            I => \N__2702\
        );

    \I__358\ : IoSpan4Mux
    port map (
            O => \N__2702\,
            I => \N__2699\
        );

    \I__357\ : Span4Mux_s2_v
    port map (
            O => \N__2699\,
            I => \N__2696\
        );

    \I__356\ : Span4Mux_v
    port map (
            O => \N__2696\,
            I => \N__2693\
        );

    \I__355\ : Odrv4
    port map (
            O => \N__2693\,
            I => \un1_D_UU_040_3\
        );

    \I__354\ : IoInMux
    port map (
            O => \N__2690\,
            I => \N__2686\
        );

    \I__353\ : IoInMux
    port map (
            O => \N__2689\,
            I => \N__2683\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__2686\,
            I => \N__2676\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__2683\,
            I => \N__2676\
        );

    \I__350\ : IoInMux
    port map (
            O => \N__2682\,
            I => \N__2673\
        );

    \I__349\ : IoInMux
    port map (
            O => \N__2681\,
            I => \N__2670\
        );

    \I__348\ : IoSpan4Mux
    port map (
            O => \N__2676\,
            I => \N__2661\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__2673\,
            I => \N__2661\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__2670\,
            I => \N__2661\
        );

    \I__345\ : IoInMux
    port map (
            O => \N__2669\,
            I => \N__2658\
        );

    \I__344\ : IoInMux
    port map (
            O => \N__2668\,
            I => \N__2655\
        );

    \I__343\ : IoSpan4Mux
    port map (
            O => \N__2661\,
            I => \N__2648\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2658\,
            I => \N__2648\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__2655\,
            I => \N__2648\
        );

    \I__340\ : IoSpan4Mux
    port map (
            O => \N__2648\,
            I => \N__2639\
        );

    \I__339\ : IoInMux
    port map (
            O => \N__2647\,
            I => \N__2636\
        );

    \I__338\ : IoInMux
    port map (
            O => \N__2646\,
            I => \N__2626\
        );

    \I__337\ : IoInMux
    port map (
            O => \N__2645\,
            I => \N__2623\
        );

    \I__336\ : IoInMux
    port map (
            O => \N__2644\,
            I => \N__2620\
        );

    \I__335\ : IoInMux
    port map (
            O => \N__2643\,
            I => \N__2617\
        );

    \I__334\ : IoInMux
    port map (
            O => \N__2642\,
            I => \N__2614\
        );

    \I__333\ : IoSpan4Mux
    port map (
            O => \N__2639\,
            I => \N__2609\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__2636\,
            I => \N__2609\
        );

    \I__331\ : IoInMux
    port map (
            O => \N__2635\,
            I => \N__2606\
        );

    \I__330\ : IoInMux
    port map (
            O => \N__2634\,
            I => \N__2603\
        );

    \I__329\ : IoInMux
    port map (
            O => \N__2633\,
            I => \N__2600\
        );

    \I__328\ : IoInMux
    port map (
            O => \N__2632\,
            I => \N__2597\
        );

    \I__327\ : IoInMux
    port map (
            O => \N__2631\,
            I => \N__2590\
        );

    \I__326\ : IoInMux
    port map (
            O => \N__2630\,
            I => \N__2587\
        );

    \I__325\ : IoInMux
    port map (
            O => \N__2629\,
            I => \N__2584\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__2626\,
            I => \N__2575\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__2623\,
            I => \N__2575\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__2620\,
            I => \N__2575\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__2617\,
            I => \N__2575\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__2614\,
            I => \N__2570\
        );

    \I__319\ : IoSpan4Mux
    port map (
            O => \N__2609\,
            I => \N__2556\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__2606\,
            I => \N__2556\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__2603\,
            I => \N__2556\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__2600\,
            I => \N__2556\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__2597\,
            I => \N__2556\
        );

    \I__314\ : IoInMux
    port map (
            O => \N__2596\,
            I => \N__2553\
        );

    \I__313\ : IoInMux
    port map (
            O => \N__2595\,
            I => \N__2550\
        );

    \I__312\ : IoInMux
    port map (
            O => \N__2594\,
            I => \N__2547\
        );

    \I__311\ : IoInMux
    port map (
            O => \N__2593\,
            I => \N__2544\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__2590\,
            I => \N__2535\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__2587\,
            I => \N__2535\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__2584\,
            I => \N__2535\
        );

    \I__307\ : IoSpan4Mux
    port map (
            O => \N__2575\,
            I => \N__2535\
        );

    \I__306\ : IoInMux
    port map (
            O => \N__2574\,
            I => \N__2532\
        );

    \I__305\ : IoInMux
    port map (
            O => \N__2573\,
            I => \N__2529\
        );

    \I__304\ : IoSpan4Mux
    port map (
            O => \N__2570\,
            I => \N__2526\
        );

    \I__303\ : IoInMux
    port map (
            O => \N__2569\,
            I => \N__2522\
        );

    \I__302\ : IoInMux
    port map (
            O => \N__2568\,
            I => \N__2519\
        );

    \I__301\ : IoInMux
    port map (
            O => \N__2567\,
            I => \N__2516\
        );

    \I__300\ : IoSpan4Mux
    port map (
            O => \N__2556\,
            I => \N__2508\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__2553\,
            I => \N__2508\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__2550\,
            I => \N__2508\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__2547\,
            I => \N__2497\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__2544\,
            I => \N__2497\
        );

    \I__295\ : IoSpan4Mux
    port map (
            O => \N__2535\,
            I => \N__2497\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__2532\,
            I => \N__2497\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__2529\,
            I => \N__2497\
        );

    \I__292\ : Span4Mux_s3_v
    port map (
            O => \N__2526\,
            I => \N__2494\
        );

    \I__291\ : IoInMux
    port map (
            O => \N__2525\,
            I => \N__2491\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__2522\,
            I => \N__2484\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__2519\,
            I => \N__2484\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__2516\,
            I => \N__2481\
        );

    \I__287\ : IoInMux
    port map (
            O => \N__2515\,
            I => \N__2478\
        );

    \I__286\ : IoSpan4Mux
    port map (
            O => \N__2508\,
            I => \N__2473\
        );

    \I__285\ : IoSpan4Mux
    port map (
            O => \N__2497\,
            I => \N__2473\
        );

    \I__284\ : Span4Mux_v
    port map (
            O => \N__2494\,
            I => \N__2468\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__2491\,
            I => \N__2468\
        );

    \I__282\ : IoInMux
    port map (
            O => \N__2490\,
            I => \N__2465\
        );

    \I__281\ : IoInMux
    port map (
            O => \N__2489\,
            I => \N__2462\
        );

    \I__280\ : Span12Mux_s9_h
    port map (
            O => \N__2484\,
            I => \N__2459\
        );

    \I__279\ : Span12Mux_s9_h
    port map (
            O => \N__2481\,
            I => \N__2456\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__2478\,
            I => \N__2453\
        );

    \I__277\ : Span4Mux_s2_h
    port map (
            O => \N__2473\,
            I => \N__2450\
        );

    \I__276\ : Span4Mux_s3_v
    port map (
            O => \N__2468\,
            I => \N__2447\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2465\,
            I => \N__2442\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__2462\,
            I => \N__2442\
        );

    \I__273\ : Span12Mux_v
    port map (
            O => \N__2459\,
            I => \N__2439\
        );

    \I__272\ : Span12Mux_v
    port map (
            O => \N__2456\,
            I => \N__2434\
        );

    \I__271\ : Span12Mux_s9_h
    port map (
            O => \N__2453\,
            I => \N__2434\
        );

    \I__270\ : Span4Mux_h
    port map (
            O => \N__2450\,
            I => \N__2429\
        );

    \I__269\ : Span4Mux_v
    port map (
            O => \N__2447\,
            I => \N__2429\
        );

    \I__268\ : Span12Mux_s2_h
    port map (
            O => \N__2442\,
            I => \N__2426\
        );

    \I__267\ : Odrv12
    port map (
            O => \N__2439\,
            I => \RnW_c_i_0\
        );

    \I__266\ : Odrv12
    port map (
            O => \N__2434\,
            I => \RnW_c_i_0\
        );

    \I__265\ : Odrv4
    port map (
            O => \N__2429\,
            I => \RnW_c_i_0\
        );

    \I__264\ : Odrv12
    port map (
            O => \N__2426\,
            I => \RnW_c_i_0\
        );

    \I__263\ : InMux
    port map (
            O => \N__2417\,
            I => \N__2414\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__2414\,
            I => \N__2411\
        );

    \I__261\ : Span4Mux_h
    port map (
            O => \N__2411\,
            I => \N__2408\
        );

    \I__260\ : Span4Mux_v
    port map (
            O => \N__2408\,
            I => \N__2405\
        );

    \I__259\ : Odrv4
    port map (
            O => \N__2405\,
            I => \A_040_c_0\
        );

    \I__258\ : IoInMux
    port map (
            O => \N__2402\,
            I => \N__2399\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__2399\,
            I => \N__2396\
        );

    \I__256\ : Span4Mux_s2_v
    port map (
            O => \N__2396\,
            I => \N__2393\
        );

    \I__255\ : Span4Mux_v
    port map (
            O => \N__2393\,
            I => \N__2390\
        );

    \I__254\ : Odrv4
    port map (
            O => \N__2390\,
            I => \A_AMIGA_c_0\
        );

    \I__253\ : InMux
    port map (
            O => \N__2387\,
            I => \N__2384\
        );

    \I__252\ : LocalMux
    port map (
            O => \N__2384\,
            I => \N__2381\
        );

    \I__251\ : Span12Mux_h
    port map (
            O => \N__2381\,
            I => \N__2378\
        );

    \I__250\ : Odrv12
    port map (
            O => \N__2378\,
            I => \A_040_c_1\
        );

    \I__249\ : CascadeMux
    port map (
            O => \N__2375\,
            I => \A_AMIGA_c_1_cascade_\
        );

    \I__248\ : InMux
    port map (
            O => \N__2372\,
            I => \N__2369\
        );

    \I__247\ : LocalMux
    port map (
            O => \N__2369\,
            I => \N__2366\
        );

    \I__246\ : Span4Mux_v
    port map (
            O => \N__2366\,
            I => \N__2363\
        );

    \I__245\ : Sp12to4
    port map (
            O => \N__2363\,
            I => \N__2360\
        );

    \I__244\ : Odrv12
    port map (
            O => \N__2360\,
            I => \D_LL_AMIGA_in_3\
        );

    \I__243\ : IoInMux
    port map (
            O => \N__2357\,
            I => \N__2354\
        );

    \I__242\ : LocalMux
    port map (
            O => \N__2354\,
            I => \N__2351\
        );

    \I__241\ : Span4Mux_s1_h
    port map (
            O => \N__2351\,
            I => \N__2348\
        );

    \I__240\ : Sp12to4
    port map (
            O => \N__2348\,
            I => \N__2345\
        );

    \I__239\ : Span12Mux_s6_v
    port map (
            O => \N__2345\,
            I => \N__2342\
        );

    \I__238\ : Span12Mux_h
    port map (
            O => \N__2342\,
            I => \N__2339\
        );

    \I__237\ : Odrv12
    port map (
            O => \N__2339\,
            I => \un1_D_LL_AMIGA_3\
        );

    \I__236\ : CascadeMux
    port map (
            O => \N__2336\,
            I => \N__2333\
        );

    \I__235\ : InMux
    port map (
            O => \N__2333\,
            I => \N__2330\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__2330\,
            I => \N__2327\
        );

    \I__233\ : Span4Mux_v
    port map (
            O => \N__2327\,
            I => \N__2324\
        );

    \I__232\ : Span4Mux_h
    port map (
            O => \N__2324\,
            I => \N__2321\
        );

    \I__231\ : Odrv4
    port map (
            O => \N__2321\,
            I => \D_LL_AMIGA_in_4\
        );

    \I__230\ : IoInMux
    port map (
            O => \N__2318\,
            I => \N__2315\
        );

    \I__229\ : LocalMux
    port map (
            O => \N__2315\,
            I => \N__2312\
        );

    \I__228\ : Sp12to4
    port map (
            O => \N__2312\,
            I => \N__2309\
        );

    \I__227\ : Span12Mux_h
    port map (
            O => \N__2309\,
            I => \N__2306\
        );

    \I__226\ : Span12Mux_h
    port map (
            O => \N__2306\,
            I => \N__2303\
        );

    \I__225\ : Odrv12
    port map (
            O => \N__2303\,
            I => \un1_D_LL_AMIGA_4\
        );

    \I__224\ : InMux
    port map (
            O => \N__2300\,
            I => \N__2297\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__2297\,
            I => \N__2294\
        );

    \I__222\ : Sp12to4
    port map (
            O => \N__2294\,
            I => \N__2291\
        );

    \I__221\ : Span12Mux_v
    port map (
            O => \N__2291\,
            I => \N__2288\
        );

    \I__220\ : Span12Mux_h
    port map (
            O => \N__2288\,
            I => \N__2285\
        );

    \I__219\ : Span12Mux_h
    port map (
            O => \N__2285\,
            I => \N__2282\
        );

    \I__218\ : Odrv12
    port map (
            O => \N__2282\,
            I => \D_UM_040_in_0\
        );

    \I__217\ : CascadeMux
    port map (
            O => \N__2279\,
            I => \N__2276\
        );

    \I__216\ : InMux
    port map (
            O => \N__2276\,
            I => \N__2272\
        );

    \I__215\ : IoInMux
    port map (
            O => \N__2275\,
            I => \N__2269\
        );

    \I__214\ : LocalMux
    port map (
            O => \N__2272\,
            I => \N__2266\
        );

    \I__213\ : LocalMux
    port map (
            O => \N__2269\,
            I => \N__2263\
        );

    \I__212\ : Span4Mux_v
    port map (
            O => \N__2266\,
            I => \N__2260\
        );

    \I__211\ : IoSpan4Mux
    port map (
            O => \N__2263\,
            I => \N__2257\
        );

    \I__210\ : Sp12to4
    port map (
            O => \N__2260\,
            I => \N__2254\
        );

    \I__209\ : Span4Mux_s2_h
    port map (
            O => \N__2257\,
            I => \N__2251\
        );

    \I__208\ : Span12Mux_h
    port map (
            O => \N__2254\,
            I => \N__2248\
        );

    \I__207\ : Sp12to4
    port map (
            O => \N__2251\,
            I => \N__2245\
        );

    \I__206\ : Span12Mux_v
    port map (
            O => \N__2248\,
            I => \N__2242\
        );

    \I__205\ : Span12Mux_h
    port map (
            O => \N__2245\,
            I => \N__2239\
        );

    \I__204\ : Span12Mux_h
    port map (
            O => \N__2242\,
            I => \N__2236\
        );

    \I__203\ : Span12Mux_h
    port map (
            O => \N__2239\,
            I => \N__2233\
        );

    \I__202\ : Odrv12
    port map (
            O => \N__2236\,
            I => \D_LL_040_in_0\
        );

    \I__201\ : Odrv12
    port map (
            O => \N__2233\,
            I => \D_LL_040_in_0\
        );

    \I__200\ : IoInMux
    port map (
            O => \N__2228\,
            I => \N__2225\
        );

    \I__199\ : LocalMux
    port map (
            O => \N__2225\,
            I => \N__2222\
        );

    \I__198\ : IoSpan4Mux
    port map (
            O => \N__2222\,
            I => \N__2219\
        );

    \I__197\ : Span4Mux_s1_h
    port map (
            O => \N__2219\,
            I => \N__2216\
        );

    \I__196\ : Span4Mux_h
    port map (
            O => \N__2216\,
            I => \N__2213\
        );

    \I__195\ : Odrv4
    port map (
            O => \N__2213\,
            I => \un1_D_UM_040_0\
        );

    \INVU111_CYCLE_SM.UU_LATCHED_nesr_5C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UU_LATCHED_nesr_5C_net\,
            I => \N__5626\
        );

    \INVU111_CYCLE_SM.UM_LATCHED_nesr_1C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UM_LATCHED_nesr_1C_net\,
            I => \N__5629\
        );

    \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net\,
            I => \N__5631\
        );

    \INVU111_CYCLE_SM.UU_LATCHED_nesr_4C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net\,
            I => \N__5623\
        );

    \INVU111_CYCLE_SM.CYCLE_STATE_0C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.CYCLE_STATE_0C_net\,
            I => \N__5624\
        );

    \INVU111_CYCLE_SM.LW_CYCLEC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.LW_CYCLEC_net\,
            I => \N__5627\
        );

    \INVU111_CYCLE_SM.UU_LATCHED_nesr_6C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UU_LATCHED_nesr_6C_net\,
            I => \N__5625\
        );

    \INVU111_CYCLE_SM.LW_CYCLE_STARTC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.LW_CYCLE_STARTC_net\,
            I => \N__5628\
        );

    \INVU111_CYCLE_SM.UM_LATCHED_nesr_2C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UM_LATCHED_nesr_2C_net\,
            I => \N__5630\
        );

    \INVU111_CYCLE_SM.TA_ENC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.TA_ENC_net\,
            I => \N__5632\
        );

    \INVU111_CYCLE_SM.TSnC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.TSnC_net\,
            I => \N__5531\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7346\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2417\,
            lcout => \A_AMIGA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__2387\,
            in1 => \N__5474\,
            in2 => \_gnd_net_\,
            in3 => \N__7345\,
            lcout => \A_AMIGA_c_1\,
            ltout => \A_AMIGA_c_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIGCUI2_LC_3_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__7082\,
            in1 => \N__6328\,
            in2 => \N__2375\,
            in3 => \N__2372\,
            lcout => \un1_D_LL_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIIEUI2_LC_3_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__6329\,
            in1 => \N__6842\,
            in2 => \N__2336\,
            in3 => \N__5795\,
            lcout => \un1_D_LL_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIKNOB2_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__6326\,
            in1 => \N__2300\,
            in2 => \N__2279\,
            in3 => \N__5796\,
            lcout => \un1_D_UM_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIOROB2_LC_3_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__5797\,
            in1 => \N__6327\,
            in2 => \N__3245\,
            in3 => \N__3227\,
            lcout => \un1_D_UM_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIMPOB2_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__3164\,
            in1 => \N__6284\,
            in2 => \N__3116\,
            in3 => \N__5851\,
            lcout => \un1_D_UM_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI26PB2_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__3076\,
            in1 => \N__6266\,
            in2 => \N__3026\,
            in3 => \N__5852\,
            lcout => \un1_D_UM_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIVEQV1_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__2981\,
            in1 => \N__6267\,
            in2 => \N__2960\,
            in3 => \N__5853\,
            lcout => \un1_D_UU_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIPJJF2_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__5883\,
            in1 => \N__6316\,
            in2 => \N__4403\,
            in3 => \N__2894\,
            lcout => \un1_D_LM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIBRQV1_LC_5_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__6292\,
            in1 => \N__2857\,
            in2 => \N__2822\,
            in3 => \N__5957\,
            lcout => \un1_D_UU_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI3JQV1_LC_5_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__6291\,
            in1 => \N__2776\,
            in2 => \N__2732\,
            in3 => \N__5956\,
            lcout => \un1_D_UU_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RnW_c_sbtinv_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5165\,
            lcout => \RnW_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIMIUI2_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__6268\,
            in1 => \N__6586\,
            in2 => \N__3596\,
            in3 => \N__5913\,
            lcout => \un1_D_LL_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNITNJF2_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__3554\,
            in1 => \N__6237\,
            in2 => \N__7393\,
            in3 => \N__5919\,
            lcout => \un1_D_LM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI1SJF2_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__6681\,
            in1 => \N__6184\,
            in2 => \N__3518\,
            in3 => \N__5949\,
            lcout => \un1_D_LM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TSn_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__5266\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4577\,
            lcout => \TSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TSnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIA6UI2_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__6317\,
            in1 => \N__3476\,
            in2 => \N__6530\,
            in3 => \N__5864\,
            lcout => \un1_D_LL_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI5LQV1_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__3437\,
            in1 => \N__3412\,
            in2 => \N__6288\,
            in3 => \N__5970\,
            lcout => \un1_D_UU_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIC8UI2_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__6998\,
            in1 => \N__6321\,
            in2 => \N__5940\,
            in3 => \N__3359\,
            lcout => \un1_D_LL_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIEAUI2_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__6322\,
            in1 => \N__4238\,
            in2 => \N__5941\,
            in3 => \N__3317\,
            lcout => \un1_D_LL_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIJDJF2_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__6302\,
            in1 => \N__6464\,
            in2 => \N__5966\,
            in3 => \N__3278\,
            lcout => \un1_D_LM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI1HQV1_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__6245\,
            in1 => \N__4166\,
            in2 => \N__4148\,
            in3 => \N__5983\,
            lcout => \un1_D_UU_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNITCQV1_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__5985\,
            in1 => \N__6247\,
            in2 => \N__4094\,
            in3 => \N__4066\,
            lcout => \un1_D_UU_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNISVOB2_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__6246\,
            in1 => \N__4000\,
            in2 => \N__3962\,
            in3 => \N__5984\,
            lcout => \un1_D_UM_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNINHJF2_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__5859\,
            in1 => \N__6230\,
            in2 => \N__4874\,
            in3 => \N__3917\,
            lcout => \un1_D_LM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIVPJF2_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__6109\,
            in1 => \N__4945\,
            in2 => \N__3890\,
            in3 => \N__5912\,
            lcout => \un1_D_LM_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIQTOB2_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__5969\,
            in1 => \N__6164\,
            in2 => \N__3854\,
            in3 => \N__3826\,
            lcout => \un1_D_UM_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI7NQV1_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__5968\,
            in1 => \N__6163\,
            in2 => \N__3767\,
            in3 => \N__3730\,
            lcout => \un1_D_UU_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIU1PB2_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__5992\,
            in1 => \N__6229\,
            in2 => \N__3686\,
            in3 => \N__3661\,
            lcout => \un1_D_UM_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIKGUI2_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__4337\,
            in1 => \N__6269\,
            in2 => \N__6392\,
            in3 => \N__5945\,
            lcout => \un1_D_LL_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIOKUI2_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__6270\,
            in1 => \N__6770\,
            in2 => \N__5967\,
            in3 => \N__4295\,
            lcout => \un1_D_LL_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_EN_RNO_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5287\,
            lcout => \U111_CYCLE_SM.RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4196\,
            in1 => \N__4237\,
            in2 => \_gnd_net_\,
            in3 => \N__7304\,
            lcout => \un1_D_UM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_EN_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000011011100"
        )
    port map (
            in0 => \N__5507\,
            in1 => \N__5363\,
            in2 => \N__4667\,
            in3 => \N__5405\,
            lcout => \U111_CYCLE_SM.TA_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TA_ENC_net\,
            ce => 'H',
            sr => \N__4247\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4224\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_2C_net\,
            ce => \N__7190\,
            sr => \N__7143\
        );

    \U111_CYCLE_SM.LW_CYCLE_START_RNO_0_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000000000"
        )
    port map (
            in0 => \N__4496\,
            in1 => \N__4523\,
            in2 => \N__4573\,
            in3 => \N__4543\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.un3_LW_CYCLE_START_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_START_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001010100000"
        )
    port map (
            in0 => \N__5309\,
            in1 => \N__7252\,
            in2 => \N__4187\,
            in3 => \N__5503\,
            lcout => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.LW_CYCLE_STARTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_1_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011001110"
        )
    port map (
            in0 => \N__5544\,
            in1 => \N__5355\,
            in2 => \N__4184\,
            in3 => \N__5400\,
            lcout => \U111_CYCLE_SM.TS_EN_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111011"
        )
    port map (
            in0 => \N__5543\,
            in1 => \N__5354\,
            in2 => \_gnd_net_\,
            in3 => \N__5401\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.N_69_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__5310\,
            in1 => \N__4569\,
            in2 => \N__4586\,
            in3 => \N__4583\,
            lcout => \U111_CYCLE_SM.TS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.LW_CYCLE_STARTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4946\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_6C_net\,
            ce => \N__7191\,
            sr => \N__7139\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4867\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_6C_net\,
            ce => \N__7191\,
            sr => \N__7139\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4393\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_6C_net\,
            ce => \N__7191\,
            sr => \N__7139\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI2RET_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011010111"
        )
    port map (
            in0 => \N__4550\,
            in1 => \N__4519\,
            in2 => \N__4495\,
            in3 => \N__7331\,
            lcout => \U111_CYCLE_SM.un1_LW_TRANS_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7333\,
            in1 => \N__4412\,
            in2 => \_gnd_net_\,
            in3 => \N__4392\,
            lcout => \un1_D_UU_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7334\,
            in1 => \N__4955\,
            in2 => \_gnd_net_\,
            in3 => \N__4944\,
            lcout => \un1_D_UU_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7332\,
            in1 => \N__4883\,
            in2 => \_gnd_net_\,
            in3 => \N__4866\,
            lcout => \un1_D_UU_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK40_THRU_LUT4_0_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5546\,
            lcout => \GB_BUFFER_CLK40_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNILFJF2_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__5926\,
            in1 => \N__6290\,
            in2 => \N__4790\,
            in3 => \N__6909\,
            lcout => \un1_D_LM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI04PB2_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__4754\,
            in1 => \N__6289\,
            in2 => \N__4732\,
            in3 => \N__5860\,
            lcout => \un1_D_UM_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_EN_RNI1DSB_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4666\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5425\,
            lcout => \U111_CYCLE_SM_TAn_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIRLJF2_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__4631\,
            in1 => \N__6265\,
            in2 => \N__5708\,
            in3 => \N__5955\,
            lcout => \un1_D_LM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__5357\,
            in1 => \N__4592\,
            in2 => \N__5315\,
            in3 => \N__5552\,
            lcout => \U111_CYCLE_SM.LW_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.LW_CYCLEC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNO_1_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010101010"
        )
    port map (
            in0 => \N__7251\,
            in1 => \N__5356\,
            in2 => \N__5447\,
            in3 => \N__5399\,
            lcout => \U111_CYCLE_SM.LW_CYCLE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5500\,
            in2 => \_gnd_net_\,
            in3 => \N__5398\,
            lcout => \U111_CYCLE_SM.A_OUT_0_sqmuxa_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__5350\,
            in1 => \N__5502\,
            in2 => \_gnd_net_\,
            in3 => \N__5545\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.N_91_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__5444\,
            in1 => \N__5312\,
            in2 => \N__5510\,
            in3 => \N__5397\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.CYCLE_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A_OUT_RNO_0_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101101010000"
        )
    port map (
            in0 => \N__5395\,
            in1 => \N__5501\,
            in2 => \N__5361\,
            in3 => \N__5458\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.A_OUT_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A_OUT_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5477\,
            in3 => \N__5311\,
            lcout => \U111_CYCLE_SM.A_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.CYCLE_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_1_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101001000000000"
        )
    port map (
            in0 => \N__5396\,
            in1 => \N__5445\,
            in2 => \N__5362\,
            in3 => \N__5314\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.CYCLE_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIFCLM_0_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__5446\,
            in1 => \N__5394\,
            in2 => \_gnd_net_\,
            in3 => \N__5346\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa\,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1_0_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111110101"
        )
    port map (
            in0 => \N__5313\,
            in1 => \_gnd_net_\,
            in2 => \N__5249\,
            in3 => \N__5098\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0\,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIGG4C2_0_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4958\,
            in3 => \N__6479\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5701\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net\,
            ce => \N__7188\,
            sr => \N__7138\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6463\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net\,
            ce => \N__7188\,
            sr => \N__7138\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6385\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net\,
            ce => \N__7188\,
            sr => \N__7138\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7316\,
            in1 => \N__6473\,
            in2 => \_gnd_net_\,
            in3 => \N__6456\,
            lcout => \un1_D_UU_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7315\,
            in1 => \N__6401\,
            in2 => \_gnd_net_\,
            in3 => \N__6384\,
            lcout => \un1_D_UM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI9PQV1_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__6244\,
            in1 => \N__6059\,
            in2 => \N__6040\,
            in3 => \N__5993\,
            lcout => \un1_D_UU_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5700\,
            in1 => \N__5669\,
            in2 => \_gnd_net_\,
            in3 => \N__7317\,
            lcout => \un1_D_UU_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK80_THRU_LUT4_0_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5639\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_CLK80_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6488\,
            in1 => \N__6507\,
            in2 => \_gnd_net_\,
            in3 => \N__7286\,
            lcout => \un1_D_UM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7287\,
            in1 => \N__6539\,
            in2 => \_gnd_net_\,
            in3 => \N__6582\,
            lcout => \un1_D_UM_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6587\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net\,
            ce => \N__7192\,
            sr => \N__7144\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6520\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net\,
            ce => \N__7192\,
            sr => \N__7144\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6996\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_1C_net\,
            ce => \N__7189\,
            sr => \N__7125\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6769\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_1C_net\,
            ce => \N__7189\,
            sr => \N__7125\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7394\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_5C_net\,
            ce => \N__7193\,
            sr => \N__7145\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7081\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_5C_net\,
            ce => \N__7193\,
            sr => \N__7145\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6838\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_5C_net\,
            ce => \N__7193\,
            sr => \N__7145\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6683\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_5C_net\,
            ce => \N__7193\,
            sr => \N__7145\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6914\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_5C_net\,
            ce => \N__7193\,
            sr => \N__7145\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7322\,
            in1 => \N__7088\,
            in2 => \_gnd_net_\,
            in3 => \N__7080\,
            lcout => \un1_D_UM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6997\,
            in1 => \N__6953\,
            in2 => \_gnd_net_\,
            in3 => \N__7321\,
            lcout => \un1_D_UM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7323\,
            in1 => \N__6923\,
            in2 => \_gnd_net_\,
            in3 => \N__6910\,
            lcout => \un1_D_UU_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7324\,
            in1 => \N__6851\,
            in2 => \_gnd_net_\,
            in3 => \N__6831\,
            lcout => \un1_D_UM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6762\,
            in1 => \N__6722\,
            in2 => \_gnd_net_\,
            in3 => \N__7325\,
            lcout => \un1_D_UM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7339\,
            in1 => \N__6692\,
            in2 => \_gnd_net_\,
            in3 => \N__6682\,
            lcout => \un1_D_UU_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7403\,
            in1 => \N__7389\,
            in2 => \_gnd_net_\,
            in3 => \N__7338\,
            lcout => \un1_D_UU_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     May 31 2025 14:22:48

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U111_TOP" view "INTERFACE"

module U111_TOP (
    D_UU_AMIGA,
    D_LL_AMIGA,
    D_UM_AMIGA,
    D_LM_AMIGA,
    D_UU_040,
    D_LM_040,
    D_UM_040,
    D_LL_040,
    A_AMIGA,
    A_040,
    SIZ,
    TEAn,
    TSn,
    RESETn,
    CLKRAMA,
    PORTSIZE,
    TEA_CPUn,
    LBENn,
    CLK40B,
    TBI_CPUn,
    TAn,
    CPUBGn,
    BUFENn,
    RnW,
    CLK80_CPU,
    BUFDIR,
    TCI_CPUn,
    TS_CPUn,
    CLKRAMB,
    CLK40A,
    TCIn,
    TBIn,
    DMAn,
    CLK40C,
    CLK40_IN,
    TACKn,
    BGn);

    inout [7:0] D_UU_AMIGA;
    inout [7:0] D_LL_AMIGA;
    inout [7:0] D_UM_AMIGA;
    inout [7:0] D_LM_AMIGA;
    inout [7:0] D_UU_040;
    inout [7:0] D_LM_040;
    inout [7:0] D_UM_040;
    inout [7:0] D_LL_040;
    output [1:0] A_AMIGA;
    input [1:0] A_040;
    input [1:0] SIZ;
    input TEAn;
    output TSn;
    input RESETn;
    output CLKRAMA;
    input PORTSIZE;
    output TEA_CPUn;
    input LBENn;
    output CLK40B;
    output TBI_CPUn;
    inout TAn;
    output CPUBGn;
    output BUFENn;
    input RnW;
    output CLK80_CPU;
    output BUFDIR;
    output TCI_CPUn;
    input TS_CPUn;
    output CLKRAMB;
    output CLK40A;
    input TCIn;
    input TBIn;
    output DMAn;
    output CLK40C;
    input CLK40_IN;
    inout TACKn;
    input BGn;

    wire N__13729;
    wire N__13713;
    wire N__13712;
    wire N__13711;
    wire N__13704;
    wire N__13703;
    wire N__13702;
    wire N__13695;
    wire N__13694;
    wire N__13693;
    wire N__13686;
    wire N__13685;
    wire N__13684;
    wire N__13677;
    wire N__13676;
    wire N__13675;
    wire N__13668;
    wire N__13667;
    wire N__13666;
    wire N__13659;
    wire N__13658;
    wire N__13657;
    wire N__13650;
    wire N__13649;
    wire N__13648;
    wire N__13641;
    wire N__13640;
    wire N__13639;
    wire N__13632;
    wire N__13631;
    wire N__13630;
    wire N__13623;
    wire N__13622;
    wire N__13621;
    wire N__13614;
    wire N__13613;
    wire N__13612;
    wire N__13605;
    wire N__13604;
    wire N__13603;
    wire N__13596;
    wire N__13595;
    wire N__13594;
    wire N__13587;
    wire N__13586;
    wire N__13585;
    wire N__13578;
    wire N__13577;
    wire N__13576;
    wire N__13569;
    wire N__13568;
    wire N__13567;
    wire N__13560;
    wire N__13559;
    wire N__13558;
    wire N__13551;
    wire N__13550;
    wire N__13549;
    wire N__13542;
    wire N__13541;
    wire N__13540;
    wire N__13533;
    wire N__13532;
    wire N__13531;
    wire N__13524;
    wire N__13523;
    wire N__13522;
    wire N__13515;
    wire N__13514;
    wire N__13513;
    wire N__13506;
    wire N__13505;
    wire N__13504;
    wire N__13497;
    wire N__13496;
    wire N__13495;
    wire N__13488;
    wire N__13487;
    wire N__13486;
    wire N__13479;
    wire N__13478;
    wire N__13477;
    wire N__13470;
    wire N__13469;
    wire N__13468;
    wire N__13461;
    wire N__13460;
    wire N__13459;
    wire N__13452;
    wire N__13451;
    wire N__13450;
    wire N__13443;
    wire N__13442;
    wire N__13441;
    wire N__13434;
    wire N__13433;
    wire N__13432;
    wire N__13425;
    wire N__13424;
    wire N__13423;
    wire N__13416;
    wire N__13415;
    wire N__13414;
    wire N__13407;
    wire N__13406;
    wire N__13405;
    wire N__13398;
    wire N__13397;
    wire N__13396;
    wire N__13389;
    wire N__13388;
    wire N__13387;
    wire N__13380;
    wire N__13379;
    wire N__13378;
    wire N__13371;
    wire N__13370;
    wire N__13369;
    wire N__13362;
    wire N__13361;
    wire N__13360;
    wire N__13353;
    wire N__13352;
    wire N__13351;
    wire N__13344;
    wire N__13343;
    wire N__13342;
    wire N__13335;
    wire N__13334;
    wire N__13333;
    wire N__13326;
    wire N__13325;
    wire N__13324;
    wire N__13317;
    wire N__13316;
    wire N__13315;
    wire N__13308;
    wire N__13307;
    wire N__13306;
    wire N__13299;
    wire N__13298;
    wire N__13297;
    wire N__13290;
    wire N__13289;
    wire N__13288;
    wire N__13281;
    wire N__13280;
    wire N__13279;
    wire N__13272;
    wire N__13271;
    wire N__13270;
    wire N__13263;
    wire N__13262;
    wire N__13261;
    wire N__13254;
    wire N__13253;
    wire N__13252;
    wire N__13245;
    wire N__13244;
    wire N__13243;
    wire N__13236;
    wire N__13235;
    wire N__13234;
    wire N__13227;
    wire N__13226;
    wire N__13225;
    wire N__13218;
    wire N__13217;
    wire N__13216;
    wire N__13209;
    wire N__13208;
    wire N__13207;
    wire N__13200;
    wire N__13199;
    wire N__13198;
    wire N__13191;
    wire N__13190;
    wire N__13189;
    wire N__13182;
    wire N__13181;
    wire N__13180;
    wire N__13173;
    wire N__13172;
    wire N__13171;
    wire N__13164;
    wire N__13163;
    wire N__13162;
    wire N__13155;
    wire N__13154;
    wire N__13153;
    wire N__13146;
    wire N__13145;
    wire N__13144;
    wire N__13137;
    wire N__13136;
    wire N__13135;
    wire N__13128;
    wire N__13127;
    wire N__13126;
    wire N__13119;
    wire N__13118;
    wire N__13117;
    wire N__13110;
    wire N__13109;
    wire N__13108;
    wire N__13101;
    wire N__13100;
    wire N__13099;
    wire N__13092;
    wire N__13091;
    wire N__13090;
    wire N__13083;
    wire N__13082;
    wire N__13081;
    wire N__13074;
    wire N__13073;
    wire N__13072;
    wire N__13065;
    wire N__13064;
    wire N__13063;
    wire N__13056;
    wire N__13055;
    wire N__13054;
    wire N__13047;
    wire N__13046;
    wire N__13045;
    wire N__13038;
    wire N__13037;
    wire N__13036;
    wire N__13029;
    wire N__13028;
    wire N__13027;
    wire N__13020;
    wire N__13019;
    wire N__13018;
    wire N__13011;
    wire N__13010;
    wire N__13009;
    wire N__13002;
    wire N__13001;
    wire N__13000;
    wire N__12993;
    wire N__12992;
    wire N__12991;
    wire N__12984;
    wire N__12983;
    wire N__12982;
    wire N__12975;
    wire N__12974;
    wire N__12973;
    wire N__12966;
    wire N__12965;
    wire N__12964;
    wire N__12957;
    wire N__12956;
    wire N__12955;
    wire N__12948;
    wire N__12947;
    wire N__12946;
    wire N__12939;
    wire N__12938;
    wire N__12937;
    wire N__12930;
    wire N__12929;
    wire N__12928;
    wire N__12921;
    wire N__12920;
    wire N__12919;
    wire N__12912;
    wire N__12911;
    wire N__12910;
    wire N__12903;
    wire N__12902;
    wire N__12901;
    wire N__12894;
    wire N__12893;
    wire N__12892;
    wire N__12885;
    wire N__12884;
    wire N__12883;
    wire N__12876;
    wire N__12875;
    wire N__12874;
    wire N__12867;
    wire N__12866;
    wire N__12865;
    wire N__12848;
    wire N__12845;
    wire N__12844;
    wire N__12843;
    wire N__12842;
    wire N__12841;
    wire N__12840;
    wire N__12839;
    wire N__12838;
    wire N__12837;
    wire N__12836;
    wire N__12835;
    wire N__12834;
    wire N__12833;
    wire N__12832;
    wire N__12831;
    wire N__12828;
    wire N__12827;
    wire N__12826;
    wire N__12825;
    wire N__12824;
    wire N__12823;
    wire N__12822;
    wire N__12821;
    wire N__12820;
    wire N__12819;
    wire N__12818;
    wire N__12817;
    wire N__12816;
    wire N__12815;
    wire N__12814;
    wire N__12813;
    wire N__12812;
    wire N__12811;
    wire N__12810;
    wire N__12809;
    wire N__12808;
    wire N__12807;
    wire N__12806;
    wire N__12805;
    wire N__12804;
    wire N__12803;
    wire N__12802;
    wire N__12801;
    wire N__12800;
    wire N__12799;
    wire N__12798;
    wire N__12797;
    wire N__12796;
    wire N__12795;
    wire N__12794;
    wire N__12793;
    wire N__12792;
    wire N__12791;
    wire N__12790;
    wire N__12789;
    wire N__12788;
    wire N__12787;
    wire N__12786;
    wire N__12785;
    wire N__12784;
    wire N__12783;
    wire N__12782;
    wire N__12659;
    wire N__12656;
    wire N__12655;
    wire N__12654;
    wire N__12653;
    wire N__12652;
    wire N__12651;
    wire N__12650;
    wire N__12649;
    wire N__12648;
    wire N__12647;
    wire N__12646;
    wire N__12645;
    wire N__12644;
    wire N__12643;
    wire N__12642;
    wire N__12641;
    wire N__12640;
    wire N__12639;
    wire N__12638;
    wire N__12637;
    wire N__12636;
    wire N__12635;
    wire N__12634;
    wire N__12633;
    wire N__12632;
    wire N__12631;
    wire N__12630;
    wire N__12629;
    wire N__12628;
    wire N__12627;
    wire N__12626;
    wire N__12625;
    wire N__12624;
    wire N__12623;
    wire N__12622;
    wire N__12621;
    wire N__12620;
    wire N__12619;
    wire N__12618;
    wire N__12617;
    wire N__12616;
    wire N__12615;
    wire N__12614;
    wire N__12613;
    wire N__12612;
    wire N__12521;
    wire N__12518;
    wire N__12515;
    wire N__12512;
    wire N__12511;
    wire N__12510;
    wire N__12509;
    wire N__12508;
    wire N__12507;
    wire N__12506;
    wire N__12505;
    wire N__12504;
    wire N__12503;
    wire N__12502;
    wire N__12501;
    wire N__12500;
    wire N__12499;
    wire N__12498;
    wire N__12497;
    wire N__12496;
    wire N__12495;
    wire N__12494;
    wire N__12493;
    wire N__12492;
    wire N__12491;
    wire N__12490;
    wire N__12489;
    wire N__12488;
    wire N__12487;
    wire N__12486;
    wire N__12485;
    wire N__12484;
    wire N__12483;
    wire N__12482;
    wire N__12481;
    wire N__12480;
    wire N__12479;
    wire N__12478;
    wire N__12477;
    wire N__12476;
    wire N__12475;
    wire N__12474;
    wire N__12473;
    wire N__12472;
    wire N__12471;
    wire N__12470;
    wire N__12469;
    wire N__12468;
    wire N__12467;
    wire N__12466;
    wire N__12465;
    wire N__12464;
    wire N__12463;
    wire N__12462;
    wire N__12459;
    wire N__12356;
    wire N__12353;
    wire N__12350;
    wire N__12347;
    wire N__12344;
    wire N__12341;
    wire N__12338;
    wire N__12335;
    wire N__12332;
    wire N__12329;
    wire N__12326;
    wire N__12323;
    wire N__12320;
    wire N__12317;
    wire N__12314;
    wire N__12311;
    wire N__12308;
    wire N__12305;
    wire N__12302;
    wire N__12299;
    wire N__12296;
    wire N__12293;
    wire N__12290;
    wire N__12287;
    wire N__12284;
    wire N__12281;
    wire N__12278;
    wire N__12275;
    wire N__12272;
    wire N__12269;
    wire N__12266;
    wire N__12263;
    wire N__12260;
    wire N__12259;
    wire N__12258;
    wire N__12257;
    wire N__12256;
    wire N__12253;
    wire N__12252;
    wire N__12251;
    wire N__12248;
    wire N__12245;
    wire N__12244;
    wire N__12243;
    wire N__12242;
    wire N__12239;
    wire N__12236;
    wire N__12231;
    wire N__12230;
    wire N__12229;
    wire N__12228;
    wire N__12227;
    wire N__12226;
    wire N__12223;
    wire N__12218;
    wire N__12217;
    wire N__12216;
    wire N__12213;
    wire N__12210;
    wire N__12207;
    wire N__12206;
    wire N__12205;
    wire N__12204;
    wire N__12203;
    wire N__12202;
    wire N__12197;
    wire N__12194;
    wire N__12189;
    wire N__12186;
    wire N__12183;
    wire N__12180;
    wire N__12175;
    wire N__12172;
    wire N__12171;
    wire N__12168;
    wire N__12167;
    wire N__12166;
    wire N__12159;
    wire N__12156;
    wire N__12153;
    wire N__12150;
    wire N__12147;
    wire N__12144;
    wire N__12127;
    wire N__12124;
    wire N__12121;
    wire N__12118;
    wire N__12117;
    wire N__12116;
    wire N__12113;
    wire N__12106;
    wire N__12095;
    wire N__12094;
    wire N__12093;
    wire N__12092;
    wire N__12091;
    wire N__12090;
    wire N__12089;
    wire N__12084;
    wire N__12081;
    wire N__12078;
    wire N__12075;
    wire N__12074;
    wire N__12073;
    wire N__12068;
    wire N__12065;
    wire N__12062;
    wire N__12059;
    wire N__12056;
    wire N__12053;
    wire N__12052;
    wire N__12051;
    wire N__12050;
    wire N__12049;
    wire N__12048;
    wire N__12047;
    wire N__12046;
    wire N__12045;
    wire N__12044;
    wire N__12043;
    wire N__12042;
    wire N__12039;
    wire N__12032;
    wire N__12029;
    wire N__12024;
    wire N__12023;
    wire N__12022;
    wire N__12017;
    wire N__12014;
    wire N__12013;
    wire N__12008;
    wire N__12005;
    wire N__11998;
    wire N__11995;
    wire N__11994;
    wire N__11993;
    wire N__11986;
    wire N__11981;
    wire N__11976;
    wire N__11975;
    wire N__11974;
    wire N__11973;
    wire N__11972;
    wire N__11971;
    wire N__11966;
    wire N__11961;
    wire N__11956;
    wire N__11951;
    wire N__11948;
    wire N__11945;
    wire N__11942;
    wire N__11939;
    wire N__11938;
    wire N__11937;
    wire N__11934;
    wire N__11929;
    wire N__11928;
    wire N__11927;
    wire N__11926;
    wire N__11925;
    wire N__11920;
    wire N__11917;
    wire N__11908;
    wire N__11905;
    wire N__11904;
    wire N__11903;
    wire N__11902;
    wire N__11901;
    wire N__11900;
    wire N__11897;
    wire N__11894;
    wire N__11891;
    wire N__11888;
    wire N__11885;
    wire N__11882;
    wire N__11877;
    wire N__11874;
    wire N__11871;
    wire N__11868;
    wire N__11865;
    wire N__11858;
    wire N__11855;
    wire N__11848;
    wire N__11845;
    wire N__11840;
    wire N__11833;
    wire N__11830;
    wire N__11825;
    wire N__11820;
    wire N__11815;
    wire N__11810;
    wire N__11801;
    wire N__11792;
    wire N__11789;
    wire N__11786;
    wire N__11779;
    wire N__11774;
    wire N__11765;
    wire N__11764;
    wire N__11761;
    wire N__11760;
    wire N__11759;
    wire N__11758;
    wire N__11755;
    wire N__11752;
    wire N__11749;
    wire N__11748;
    wire N__11745;
    wire N__11744;
    wire N__11741;
    wire N__11740;
    wire N__11739;
    wire N__11734;
    wire N__11731;
    wire N__11726;
    wire N__11723;
    wire N__11720;
    wire N__11717;
    wire N__11716;
    wire N__11715;
    wire N__11712;
    wire N__11711;
    wire N__11710;
    wire N__11709;
    wire N__11708;
    wire N__11707;
    wire N__11706;
    wire N__11705;
    wire N__11704;
    wire N__11703;
    wire N__11692;
    wire N__11689;
    wire N__11688;
    wire N__11685;
    wire N__11684;
    wire N__11677;
    wire N__11674;
    wire N__11671;
    wire N__11668;
    wire N__11667;
    wire N__11666;
    wire N__11663;
    wire N__11662;
    wire N__11659;
    wire N__11656;
    wire N__11655;
    wire N__11654;
    wire N__11651;
    wire N__11650;
    wire N__11649;
    wire N__11646;
    wire N__11641;
    wire N__11636;
    wire N__11633;
    wire N__11632;
    wire N__11631;
    wire N__11630;
    wire N__11623;
    wire N__11618;
    wire N__11609;
    wire N__11608;
    wire N__11607;
    wire N__11606;
    wire N__11605;
    wire N__11602;
    wire N__11601;
    wire N__11598;
    wire N__11597;
    wire N__11596;
    wire N__11595;
    wire N__11594;
    wire N__11593;
    wire N__11590;
    wire N__11589;
    wire N__11588;
    wire N__11587;
    wire N__11586;
    wire N__11585;
    wire N__11584;
    wire N__11581;
    wire N__11576;
    wire N__11573;
    wire N__11566;
    wire N__11561;
    wire N__11560;
    wire N__11559;
    wire N__11558;
    wire N__11555;
    wire N__11554;
    wire N__11547;
    wire N__11544;
    wire N__11539;
    wire N__11538;
    wire N__11537;
    wire N__11536;
    wire N__11535;
    wire N__11532;
    wire N__11529;
    wire N__11526;
    wire N__11523;
    wire N__11522;
    wire N__11515;
    wire N__11514;
    wire N__11513;
    wire N__11508;
    wire N__11507;
    wire N__11506;
    wire N__11505;
    wire N__11502;
    wire N__11499;
    wire N__11496;
    wire N__11493;
    wire N__11490;
    wire N__11489;
    wire N__11488;
    wire N__11485;
    wire N__11482;
    wire N__11479;
    wire N__11474;
    wire N__11469;
    wire N__11466;
    wire N__11461;
    wire N__11458;
    wire N__11457;
    wire N__11454;
    wire N__11453;
    wire N__11448;
    wire N__11445;
    wire N__11442;
    wire N__11435;
    wire N__11432;
    wire N__11425;
    wire N__11422;
    wire N__11419;
    wire N__11416;
    wire N__11413;
    wire N__11410;
    wire N__11407;
    wire N__11404;
    wire N__11401;
    wire N__11396;
    wire N__11393;
    wire N__11390;
    wire N__11383;
    wire N__11380;
    wire N__11377;
    wire N__11374;
    wire N__11371;
    wire N__11364;
    wire N__11361;
    wire N__11356;
    wire N__11353;
    wire N__11346;
    wire N__11343;
    wire N__11342;
    wire N__11339;
    wire N__11334;
    wire N__11327;
    wire N__11324;
    wire N__11321;
    wire N__11316;
    wire N__11309;
    wire N__11306;
    wire N__11303;
    wire N__11300;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11284;
    wire N__11279;
    wire N__11276;
    wire N__11271;
    wire N__11268;
    wire N__11265;
    wire N__11262;
    wire N__11259;
    wire N__11254;
    wire N__11251;
    wire N__11246;
    wire N__11241;
    wire N__11238;
    wire N__11233;
    wire N__11230;
    wire N__11227;
    wire N__11224;
    wire N__11221;
    wire N__11216;
    wire N__11211;
    wire N__11204;
    wire N__11199;
    wire N__11194;
    wire N__11183;
    wire N__11182;
    wire N__11181;
    wire N__11178;
    wire N__11175;
    wire N__11174;
    wire N__11169;
    wire N__11168;
    wire N__11167;
    wire N__11166;
    wire N__11163;
    wire N__11162;
    wire N__11161;
    wire N__11158;
    wire N__11157;
    wire N__11154;
    wire N__11151;
    wire N__11150;
    wire N__11149;
    wire N__11148;
    wire N__11145;
    wire N__11144;
    wire N__11143;
    wire N__11142;
    wire N__11139;
    wire N__11138;
    wire N__11137;
    wire N__11134;
    wire N__11133;
    wire N__11132;
    wire N__11131;
    wire N__11130;
    wire N__11127;
    wire N__11126;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11114;
    wire N__11113;
    wire N__11110;
    wire N__11109;
    wire N__11104;
    wire N__11101;
    wire N__11098;
    wire N__11095;
    wire N__11092;
    wire N__11087;
    wire N__11084;
    wire N__11083;
    wire N__11080;
    wire N__11079;
    wire N__11078;
    wire N__11077;
    wire N__11076;
    wire N__11073;
    wire N__11070;
    wire N__11069;
    wire N__11068;
    wire N__11067;
    wire N__11066;
    wire N__11065;
    wire N__11064;
    wire N__11061;
    wire N__11058;
    wire N__11055;
    wire N__11054;
    wire N__11053;
    wire N__11050;
    wire N__11047;
    wire N__11044;
    wire N__11039;
    wire N__11038;
    wire N__11037;
    wire N__11034;
    wire N__11031;
    wire N__11028;
    wire N__11025;
    wire N__11024;
    wire N__11023;
    wire N__11016;
    wire N__11007;
    wire N__11004;
    wire N__11001;
    wire N__10998;
    wire N__10995;
    wire N__10994;
    wire N__10993;
    wire N__10992;
    wire N__10989;
    wire N__10986;
    wire N__10983;
    wire N__10980;
    wire N__10977;
    wire N__10974;
    wire N__10973;
    wire N__10970;
    wire N__10969;
    wire N__10968;
    wire N__10967;
    wire N__10966;
    wire N__10965;
    wire N__10962;
    wire N__10961;
    wire N__10958;
    wire N__10955;
    wire N__10954;
    wire N__10953;
    wire N__10946;
    wire N__10943;
    wire N__10940;
    wire N__10935;
    wire N__10932;
    wire N__10929;
    wire N__10926;
    wire N__10923;
    wire N__10918;
    wire N__10913;
    wire N__10908;
    wire N__10905;
    wire N__10894;
    wire N__10891;
    wire N__10888;
    wire N__10885;
    wire N__10884;
    wire N__10883;
    wire N__10880;
    wire N__10877;
    wire N__10876;
    wire N__10871;
    wire N__10866;
    wire N__10859;
    wire N__10856;
    wire N__10855;
    wire N__10854;
    wire N__10853;
    wire N__10852;
    wire N__10851;
    wire N__10848;
    wire N__10847;
    wire N__10844;
    wire N__10843;
    wire N__10840;
    wire N__10839;
    wire N__10836;
    wire N__10831;
    wire N__10828;
    wire N__10825;
    wire N__10824;
    wire N__10821;
    wire N__10820;
    wire N__10813;
    wire N__10810;
    wire N__10801;
    wire N__10794;
    wire N__10785;
    wire N__10782;
    wire N__10779;
    wire N__10776;
    wire N__10771;
    wire N__10768;
    wire N__10765;
    wire N__10758;
    wire N__10751;
    wire N__10746;
    wire N__10737;
    wire N__10732;
    wire N__10725;
    wire N__10718;
    wire N__10715;
    wire N__10712;
    wire N__10707;
    wire N__10704;
    wire N__10703;
    wire N__10694;
    wire N__10693;
    wire N__10690;
    wire N__10687;
    wire N__10686;
    wire N__10683;
    wire N__10672;
    wire N__10669;
    wire N__10666;
    wire N__10663;
    wire N__10658;
    wire N__10655;
    wire N__10652;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10640;
    wire N__10637;
    wire N__10634;
    wire N__10625;
    wire N__10622;
    wire N__10613;
    wire N__10606;
    wire N__10603;
    wire N__10596;
    wire N__10593;
    wire N__10586;
    wire N__10585;
    wire N__10584;
    wire N__10583;
    wire N__10582;
    wire N__10581;
    wire N__10580;
    wire N__10577;
    wire N__10574;
    wire N__10573;
    wire N__10572;
    wire N__10571;
    wire N__10570;
    wire N__10569;
    wire N__10568;
    wire N__10567;
    wire N__10564;
    wire N__10561;
    wire N__10558;
    wire N__10555;
    wire N__10554;
    wire N__10551;
    wire N__10550;
    wire N__10549;
    wire N__10548;
    wire N__10545;
    wire N__10542;
    wire N__10539;
    wire N__10536;
    wire N__10535;
    wire N__10532;
    wire N__10529;
    wire N__10528;
    wire N__10527;
    wire N__10524;
    wire N__10521;
    wire N__10518;
    wire N__10511;
    wire N__10508;
    wire N__10505;
    wire N__10504;
    wire N__10503;
    wire N__10502;
    wire N__10499;
    wire N__10498;
    wire N__10495;
    wire N__10494;
    wire N__10493;
    wire N__10490;
    wire N__10487;
    wire N__10486;
    wire N__10485;
    wire N__10478;
    wire N__10473;
    wire N__10470;
    wire N__10465;
    wire N__10462;
    wire N__10461;
    wire N__10458;
    wire N__10455;
    wire N__10454;
    wire N__10451;
    wire N__10450;
    wire N__10449;
    wire N__10448;
    wire N__10447;
    wire N__10446;
    wire N__10445;
    wire N__10444;
    wire N__10443;
    wire N__10442;
    wire N__10441;
    wire N__10434;
    wire N__10431;
    wire N__10428;
    wire N__10425;
    wire N__10422;
    wire N__10419;
    wire N__10416;
    wire N__10411;
    wire N__10406;
    wire N__10403;
    wire N__10400;
    wire N__10395;
    wire N__10392;
    wire N__10389;
    wire N__10386;
    wire N__10383;
    wire N__10382;
    wire N__10381;
    wire N__10376;
    wire N__10373;
    wire N__10372;
    wire N__10369;
    wire N__10366;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10351;
    wire N__10350;
    wire N__10347;
    wire N__10340;
    wire N__10339;
    wire N__10338;
    wire N__10337;
    wire N__10336;
    wire N__10327;
    wire N__10312;
    wire N__10309;
    wire N__10300;
    wire N__10297;
    wire N__10294;
    wire N__10291;
    wire N__10288;
    wire N__10285;
    wire N__10282;
    wire N__10277;
    wire N__10274;
    wire N__10271;
    wire N__10268;
    wire N__10265;
    wire N__10262;
    wire N__10257;
    wire N__10252;
    wire N__10251;
    wire N__10250;
    wire N__10249;
    wire N__10248;
    wire N__10245;
    wire N__10242;
    wire N__10241;
    wire N__10240;
    wire N__10239;
    wire N__10238;
    wire N__10237;
    wire N__10236;
    wire N__10235;
    wire N__10234;
    wire N__10233;
    wire N__10232;
    wire N__10227;
    wire N__10222;
    wire N__10217;
    wire N__10212;
    wire N__10209;
    wire N__10206;
    wire N__10201;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10185;
    wire N__10176;
    wire N__10171;
    wire N__10170;
    wire N__10167;
    wire N__10164;
    wire N__10157;
    wire N__10152;
    wire N__10149;
    wire N__10148;
    wire N__10145;
    wire N__10142;
    wire N__10137;
    wire N__10134;
    wire N__10131;
    wire N__10128;
    wire N__10123;
    wire N__10116;
    wire N__10111;
    wire N__10108;
    wire N__10101;
    wire N__10098;
    wire N__10095;
    wire N__10088;
    wire N__10085;
    wire N__10082;
    wire N__10079;
    wire N__10074;
    wire N__10069;
    wire N__10062;
    wire N__10053;
    wire N__10050;
    wire N__10045;
    wire N__10042;
    wire N__10037;
    wire N__10028;
    wire N__10025;
    wire N__10022;
    wire N__10019;
    wire N__10016;
    wire N__10013;
    wire N__10010;
    wire N__10007;
    wire N__10004;
    wire N__10001;
    wire N__9998;
    wire N__9995;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9983;
    wire N__9980;
    wire N__9977;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9965;
    wire N__9962;
    wire N__9959;
    wire N__9956;
    wire N__9953;
    wire N__9950;
    wire N__9947;
    wire N__9944;
    wire N__9941;
    wire N__9938;
    wire N__9935;
    wire N__9932;
    wire N__9929;
    wire N__9926;
    wire N__9923;
    wire N__9920;
    wire N__9917;
    wire N__9914;
    wire N__9911;
    wire N__9908;
    wire N__9905;
    wire N__9902;
    wire N__9899;
    wire N__9896;
    wire N__9893;
    wire N__9890;
    wire N__9887;
    wire N__9884;
    wire N__9881;
    wire N__9878;
    wire N__9875;
    wire N__9872;
    wire N__9869;
    wire N__9866;
    wire N__9863;
    wire N__9860;
    wire N__9857;
    wire N__9854;
    wire N__9851;
    wire N__9848;
    wire N__9845;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9830;
    wire N__9827;
    wire N__9824;
    wire N__9821;
    wire N__9818;
    wire N__9815;
    wire N__9812;
    wire N__9809;
    wire N__9806;
    wire N__9803;
    wire N__9800;
    wire N__9797;
    wire N__9794;
    wire N__9791;
    wire N__9788;
    wire N__9785;
    wire N__9782;
    wire N__9779;
    wire N__9776;
    wire N__9773;
    wire N__9770;
    wire N__9767;
    wire N__9764;
    wire N__9761;
    wire N__9758;
    wire N__9755;
    wire N__9752;
    wire N__9749;
    wire N__9746;
    wire N__9743;
    wire N__9740;
    wire N__9737;
    wire N__9734;
    wire N__9731;
    wire N__9728;
    wire N__9725;
    wire N__9722;
    wire N__9719;
    wire N__9716;
    wire N__9713;
    wire N__9710;
    wire N__9707;
    wire N__9704;
    wire N__9701;
    wire N__9698;
    wire N__9695;
    wire N__9692;
    wire N__9689;
    wire N__9686;
    wire N__9683;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9671;
    wire N__9668;
    wire N__9665;
    wire N__9662;
    wire N__9659;
    wire N__9656;
    wire N__9653;
    wire N__9650;
    wire N__9647;
    wire N__9644;
    wire N__9641;
    wire N__9638;
    wire N__9635;
    wire N__9632;
    wire N__9629;
    wire N__9626;
    wire N__9623;
    wire N__9620;
    wire N__9617;
    wire N__9616;
    wire N__9613;
    wire N__9610;
    wire N__9607;
    wire N__9606;
    wire N__9603;
    wire N__9600;
    wire N__9597;
    wire N__9596;
    wire N__9593;
    wire N__9588;
    wire N__9585;
    wire N__9582;
    wire N__9579;
    wire N__9576;
    wire N__9573;
    wire N__9570;
    wire N__9567;
    wire N__9564;
    wire N__9561;
    wire N__9558;
    wire N__9551;
    wire N__9548;
    wire N__9545;
    wire N__9542;
    wire N__9539;
    wire N__9536;
    wire N__9533;
    wire N__9530;
    wire N__9527;
    wire N__9524;
    wire N__9521;
    wire N__9518;
    wire N__9515;
    wire N__9512;
    wire N__9509;
    wire N__9506;
    wire N__9503;
    wire N__9500;
    wire N__9497;
    wire N__9494;
    wire N__9491;
    wire N__9488;
    wire N__9485;
    wire N__9482;
    wire N__9479;
    wire N__9476;
    wire N__9473;
    wire N__9470;
    wire N__9467;
    wire N__9464;
    wire N__9461;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9422;
    wire N__9419;
    wire N__9416;
    wire N__9413;
    wire N__9410;
    wire N__9407;
    wire N__9404;
    wire N__9401;
    wire N__9398;
    wire N__9395;
    wire N__9392;
    wire N__9391;
    wire N__9388;
    wire N__9385;
    wire N__9384;
    wire N__9381;
    wire N__9378;
    wire N__9375;
    wire N__9372;
    wire N__9367;
    wire N__9362;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9350;
    wire N__9347;
    wire N__9344;
    wire N__9341;
    wire N__9338;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9328;
    wire N__9325;
    wire N__9322;
    wire N__9321;
    wire N__9318;
    wire N__9315;
    wire N__9312;
    wire N__9309;
    wire N__9306;
    wire N__9303;
    wire N__9296;
    wire N__9293;
    wire N__9290;
    wire N__9287;
    wire N__9284;
    wire N__9281;
    wire N__9278;
    wire N__9275;
    wire N__9272;
    wire N__9269;
    wire N__9268;
    wire N__9265;
    wire N__9262;
    wire N__9259;
    wire N__9256;
    wire N__9253;
    wire N__9250;
    wire N__9247;
    wire N__9244;
    wire N__9241;
    wire N__9238;
    wire N__9235;
    wire N__9232;
    wire N__9229;
    wire N__9224;
    wire N__9221;
    wire N__9218;
    wire N__9215;
    wire N__9212;
    wire N__9209;
    wire N__9206;
    wire N__9203;
    wire N__9200;
    wire N__9197;
    wire N__9194;
    wire N__9191;
    wire N__9188;
    wire N__9185;
    wire N__9182;
    wire N__9179;
    wire N__9176;
    wire N__9173;
    wire N__9170;
    wire N__9167;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9155;
    wire N__9154;
    wire N__9151;
    wire N__9148;
    wire N__9145;
    wire N__9142;
    wire N__9139;
    wire N__9136;
    wire N__9131;
    wire N__9128;
    wire N__9125;
    wire N__9122;
    wire N__9119;
    wire N__9116;
    wire N__9113;
    wire N__9110;
    wire N__9109;
    wire N__9108;
    wire N__9107;
    wire N__9106;
    wire N__9105;
    wire N__9104;
    wire N__9097;
    wire N__9096;
    wire N__9095;
    wire N__9092;
    wire N__9091;
    wire N__9090;
    wire N__9089;
    wire N__9086;
    wire N__9085;
    wire N__9080;
    wire N__9077;
    wire N__9074;
    wire N__9071;
    wire N__9068;
    wire N__9063;
    wire N__9056;
    wire N__9053;
    wire N__9052;
    wire N__9051;
    wire N__9046;
    wire N__9043;
    wire N__9038;
    wire N__9033;
    wire N__9030;
    wire N__9027;
    wire N__9026;
    wire N__9025;
    wire N__9022;
    wire N__9011;
    wire N__9008;
    wire N__9005;
    wire N__9002;
    wire N__8999;
    wire N__8996;
    wire N__8993;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8971;
    wire N__8968;
    wire N__8967;
    wire N__8964;
    wire N__8961;
    wire N__8958;
    wire N__8955;
    wire N__8952;
    wire N__8949;
    wire N__8946;
    wire N__8943;
    wire N__8940;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8924;
    wire N__8921;
    wire N__8918;
    wire N__8915;
    wire N__8912;
    wire N__8909;
    wire N__8906;
    wire N__8903;
    wire N__8900;
    wire N__8897;
    wire N__8894;
    wire N__8891;
    wire N__8890;
    wire N__8887;
    wire N__8884;
    wire N__8881;
    wire N__8878;
    wire N__8875;
    wire N__8872;
    wire N__8869;
    wire N__8866;
    wire N__8863;
    wire N__8860;
    wire N__8857;
    wire N__8854;
    wire N__8851;
    wire N__8848;
    wire N__8843;
    wire N__8840;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8828;
    wire N__8827;
    wire N__8824;
    wire N__8823;
    wire N__8822;
    wire N__8821;
    wire N__8818;
    wire N__8817;
    wire N__8816;
    wire N__8815;
    wire N__8812;
    wire N__8809;
    wire N__8808;
    wire N__8807;
    wire N__8804;
    wire N__8801;
    wire N__8800;
    wire N__8799;
    wire N__8798;
    wire N__8797;
    wire N__8796;
    wire N__8793;
    wire N__8792;
    wire N__8791;
    wire N__8788;
    wire N__8785;
    wire N__8782;
    wire N__8781;
    wire N__8776;
    wire N__8773;
    wire N__8770;
    wire N__8769;
    wire N__8768;
    wire N__8763;
    wire N__8758;
    wire N__8757;
    wire N__8756;
    wire N__8751;
    wire N__8748;
    wire N__8747;
    wire N__8746;
    wire N__8745;
    wire N__8742;
    wire N__8741;
    wire N__8736;
    wire N__8735;
    wire N__8734;
    wire N__8731;
    wire N__8728;
    wire N__8725;
    wire N__8722;
    wire N__8721;
    wire N__8714;
    wire N__8711;
    wire N__8710;
    wire N__8707;
    wire N__8702;
    wire N__8699;
    wire N__8696;
    wire N__8691;
    wire N__8688;
    wire N__8685;
    wire N__8682;
    wire N__8679;
    wire N__8676;
    wire N__8673;
    wire N__8670;
    wire N__8667;
    wire N__8666;
    wire N__8657;
    wire N__8654;
    wire N__8649;
    wire N__8646;
    wire N__8645;
    wire N__8642;
    wire N__8637;
    wire N__8634;
    wire N__8625;
    wire N__8616;
    wire N__8613;
    wire N__8610;
    wire N__8605;
    wire N__8600;
    wire N__8597;
    wire N__8596;
    wire N__8593;
    wire N__8588;
    wire N__8583;
    wire N__8578;
    wire N__8571;
    wire N__8568;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8543;
    wire N__8540;
    wire N__8537;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8527;
    wire N__8524;
    wire N__8521;
    wire N__8518;
    wire N__8515;
    wire N__8512;
    wire N__8509;
    wire N__8506;
    wire N__8503;
    wire N__8498;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8464;
    wire N__8461;
    wire N__8458;
    wire N__8457;
    wire N__8454;
    wire N__8451;
    wire N__8448;
    wire N__8445;
    wire N__8440;
    wire N__8437;
    wire N__8434;
    wire N__8431;
    wire N__8428;
    wire N__8425;
    wire N__8422;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire N__8402;
    wire N__8399;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8384;
    wire N__8381;
    wire N__8378;
    wire N__8375;
    wire N__8372;
    wire N__8371;
    wire N__8370;
    wire N__8367;
    wire N__8364;
    wire N__8361;
    wire N__8358;
    wire N__8353;
    wire N__8350;
    wire N__8347;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8333;
    wire N__8330;
    wire N__8327;
    wire N__8324;
    wire N__8321;
    wire N__8318;
    wire N__8315;
    wire N__8312;
    wire N__8311;
    wire N__8310;
    wire N__8307;
    wire N__8304;
    wire N__8301;
    wire N__8296;
    wire N__8293;
    wire N__8290;
    wire N__8287;
    wire N__8284;
    wire N__8281;
    wire N__8276;
    wire N__8273;
    wire N__8270;
    wire N__8267;
    wire N__8264;
    wire N__8261;
    wire N__8260;
    wire N__8257;
    wire N__8256;
    wire N__8253;
    wire N__8250;
    wire N__8247;
    wire N__8244;
    wire N__8241;
    wire N__8238;
    wire N__8235;
    wire N__8232;
    wire N__8229;
    wire N__8226;
    wire N__8223;
    wire N__8218;
    wire N__8213;
    wire N__8210;
    wire N__8207;
    wire N__8204;
    wire N__8201;
    wire N__8198;
    wire N__8195;
    wire N__8192;
    wire N__8189;
    wire N__8186;
    wire N__8183;
    wire N__8180;
    wire N__8177;
    wire N__8174;
    wire N__8171;
    wire N__8168;
    wire N__8165;
    wire N__8162;
    wire N__8159;
    wire N__8156;
    wire N__8155;
    wire N__8152;
    wire N__8149;
    wire N__8146;
    wire N__8143;
    wire N__8140;
    wire N__8137;
    wire N__8134;
    wire N__8131;
    wire N__8128;
    wire N__8125;
    wire N__8122;
    wire N__8117;
    wire N__8114;
    wire N__8111;
    wire N__8108;
    wire N__8105;
    wire N__8102;
    wire N__8099;
    wire N__8096;
    wire N__8093;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8081;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8069;
    wire N__8068;
    wire N__8065;
    wire N__8062;
    wire N__8059;
    wire N__8056;
    wire N__8053;
    wire N__8050;
    wire N__8047;
    wire N__8044;
    wire N__8041;
    wire N__8038;
    wire N__8035;
    wire N__8032;
    wire N__8027;
    wire N__8024;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8012;
    wire N__8009;
    wire N__8006;
    wire N__8005;
    wire N__8002;
    wire N__7999;
    wire N__7996;
    wire N__7993;
    wire N__7992;
    wire N__7989;
    wire N__7986;
    wire N__7983;
    wire N__7980;
    wire N__7975;
    wire N__7970;
    wire N__7967;
    wire N__7964;
    wire N__7961;
    wire N__7958;
    wire N__7955;
    wire N__7952;
    wire N__7949;
    wire N__7946;
    wire N__7943;
    wire N__7940;
    wire N__7937;
    wire N__7934;
    wire N__7931;
    wire N__7928;
    wire N__7927;
    wire N__7924;
    wire N__7921;
    wire N__7920;
    wire N__7917;
    wire N__7914;
    wire N__7911;
    wire N__7904;
    wire N__7901;
    wire N__7898;
    wire N__7895;
    wire N__7892;
    wire N__7889;
    wire N__7886;
    wire N__7883;
    wire N__7880;
    wire N__7877;
    wire N__7874;
    wire N__7871;
    wire N__7868;
    wire N__7867;
    wire N__7866;
    wire N__7865;
    wire N__7862;
    wire N__7859;
    wire N__7858;
    wire N__7857;
    wire N__7854;
    wire N__7851;
    wire N__7848;
    wire N__7845;
    wire N__7842;
    wire N__7839;
    wire N__7836;
    wire N__7833;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7814;
    wire N__7805;
    wire N__7802;
    wire N__7799;
    wire N__7798;
    wire N__7797;
    wire N__7796;
    wire N__7795;
    wire N__7794;
    wire N__7791;
    wire N__7788;
    wire N__7785;
    wire N__7782;
    wire N__7779;
    wire N__7776;
    wire N__7763;
    wire N__7760;
    wire N__7757;
    wire N__7754;
    wire N__7751;
    wire N__7750;
    wire N__7747;
    wire N__7744;
    wire N__7741;
    wire N__7738;
    wire N__7735;
    wire N__7732;
    wire N__7729;
    wire N__7726;
    wire N__7723;
    wire N__7720;
    wire N__7717;
    wire N__7714;
    wire N__7709;
    wire N__7706;
    wire N__7703;
    wire N__7700;
    wire N__7699;
    wire N__7698;
    wire N__7695;
    wire N__7692;
    wire N__7689;
    wire N__7684;
    wire N__7681;
    wire N__7678;
    wire N__7675;
    wire N__7672;
    wire N__7669;
    wire N__7664;
    wire N__7661;
    wire N__7658;
    wire N__7655;
    wire N__7652;
    wire N__7649;
    wire N__7646;
    wire N__7643;
    wire N__7640;
    wire N__7637;
    wire N__7634;
    wire N__7631;
    wire N__7628;
    wire N__7625;
    wire N__7622;
    wire N__7619;
    wire N__7616;
    wire N__7613;
    wire N__7610;
    wire N__7607;
    wire N__7604;
    wire N__7601;
    wire N__7600;
    wire N__7599;
    wire N__7596;
    wire N__7593;
    wire N__7590;
    wire N__7585;
    wire N__7582;
    wire N__7579;
    wire N__7576;
    wire N__7573;
    wire N__7570;
    wire N__7567;
    wire N__7562;
    wire N__7559;
    wire N__7556;
    wire N__7553;
    wire N__7550;
    wire N__7547;
    wire N__7544;
    wire N__7541;
    wire N__7540;
    wire N__7537;
    wire N__7536;
    wire N__7533;
    wire N__7530;
    wire N__7527;
    wire N__7524;
    wire N__7519;
    wire N__7516;
    wire N__7513;
    wire N__7510;
    wire N__7507;
    wire N__7504;
    wire N__7501;
    wire N__7498;
    wire N__7495;
    wire N__7490;
    wire N__7487;
    wire N__7484;
    wire N__7481;
    wire N__7478;
    wire N__7475;
    wire N__7472;
    wire N__7469;
    wire N__7466;
    wire N__7463;
    wire N__7460;
    wire N__7457;
    wire N__7454;
    wire N__7451;
    wire N__7448;
    wire N__7445;
    wire N__7442;
    wire N__7439;
    wire N__7436;
    wire N__7433;
    wire N__7430;
    wire N__7427;
    wire N__7424;
    wire N__7421;
    wire N__7418;
    wire N__7415;
    wire N__7414;
    wire N__7411;
    wire N__7410;
    wire N__7409;
    wire N__7406;
    wire N__7405;
    wire N__7402;
    wire N__7399;
    wire N__7396;
    wire N__7391;
    wire N__7388;
    wire N__7387;
    wire N__7386;
    wire N__7383;
    wire N__7378;
    wire N__7375;
    wire N__7372;
    wire N__7369;
    wire N__7368;
    wire N__7363;
    wire N__7356;
    wire N__7353;
    wire N__7346;
    wire N__7343;
    wire N__7340;
    wire N__7337;
    wire N__7334;
    wire N__7333;
    wire N__7332;
    wire N__7331;
    wire N__7330;
    wire N__7329;
    wire N__7326;
    wire N__7323;
    wire N__7320;
    wire N__7317;
    wire N__7312;
    wire N__7311;
    wire N__7308;
    wire N__7299;
    wire N__7296;
    wire N__7293;
    wire N__7288;
    wire N__7285;
    wire N__7282;
    wire N__7279;
    wire N__7276;
    wire N__7271;
    wire N__7268;
    wire N__7267;
    wire N__7264;
    wire N__7261;
    wire N__7256;
    wire N__7255;
    wire N__7254;
    wire N__7253;
    wire N__7250;
    wire N__7247;
    wire N__7246;
    wire N__7243;
    wire N__7242;
    wire N__7241;
    wire N__7240;
    wire N__7237;
    wire N__7232;
    wire N__7227;
    wire N__7224;
    wire N__7221;
    wire N__7218;
    wire N__7207;
    wire N__7204;
    wire N__7201;
    wire N__7198;
    wire N__7195;
    wire N__7190;
    wire N__7187;
    wire N__7186;
    wire N__7183;
    wire N__7180;
    wire N__7177;
    wire N__7174;
    wire N__7169;
    wire N__7166;
    wire N__7165;
    wire N__7162;
    wire N__7161;
    wire N__7158;
    wire N__7155;
    wire N__7154;
    wire N__7151;
    wire N__7150;
    wire N__7145;
    wire N__7142;
    wire N__7139;
    wire N__7136;
    wire N__7127;
    wire N__7124;
    wire N__7123;
    wire N__7120;
    wire N__7117;
    wire N__7114;
    wire N__7111;
    wire N__7106;
    wire N__7103;
    wire N__7100;
    wire N__7097;
    wire N__7094;
    wire N__7091;
    wire N__7088;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7076;
    wire N__7073;
    wire N__7070;
    wire N__7067;
    wire N__7064;
    wire N__7061;
    wire N__7058;
    wire N__7055;
    wire N__7052;
    wire N__7049;
    wire N__7046;
    wire N__7043;
    wire N__7040;
    wire N__7037;
    wire N__7034;
    wire N__7031;
    wire N__7030;
    wire N__7029;
    wire N__7026;
    wire N__7023;
    wire N__7020;
    wire N__7017;
    wire N__7014;
    wire N__7011;
    wire N__7006;
    wire N__7003;
    wire N__6998;
    wire N__6995;
    wire N__6992;
    wire N__6989;
    wire N__6986;
    wire N__6983;
    wire N__6980;
    wire N__6977;
    wire N__6974;
    wire N__6971;
    wire N__6968;
    wire N__6965;
    wire N__6964;
    wire N__6963;
    wire N__6960;
    wire N__6957;
    wire N__6954;
    wire N__6949;
    wire N__6946;
    wire N__6943;
    wire N__6940;
    wire N__6937;
    wire N__6934;
    wire N__6931;
    wire N__6926;
    wire N__6923;
    wire N__6920;
    wire N__6917;
    wire N__6914;
    wire N__6911;
    wire N__6908;
    wire N__6905;
    wire N__6902;
    wire N__6899;
    wire N__6896;
    wire N__6893;
    wire N__6890;
    wire N__6887;
    wire N__6886;
    wire N__6883;
    wire N__6880;
    wire N__6877;
    wire N__6874;
    wire N__6871;
    wire N__6868;
    wire N__6867;
    wire N__6864;
    wire N__6861;
    wire N__6858;
    wire N__6855;
    wire N__6850;
    wire N__6847;
    wire N__6844;
    wire N__6839;
    wire N__6836;
    wire N__6833;
    wire N__6830;
    wire N__6827;
    wire N__6824;
    wire N__6821;
    wire N__6818;
    wire N__6815;
    wire N__6812;
    wire N__6809;
    wire N__6806;
    wire N__6803;
    wire N__6800;
    wire N__6797;
    wire N__6794;
    wire N__6791;
    wire N__6788;
    wire N__6785;
    wire N__6782;
    wire N__6779;
    wire N__6776;
    wire N__6773;
    wire N__6770;
    wire N__6767;
    wire N__6766;
    wire N__6765;
    wire N__6764;
    wire N__6761;
    wire N__6760;
    wire N__6757;
    wire N__6754;
    wire N__6751;
    wire N__6748;
    wire N__6745;
    wire N__6734;
    wire N__6731;
    wire N__6728;
    wire N__6725;
    wire N__6722;
    wire N__6719;
    wire N__6716;
    wire N__6713;
    wire N__6712;
    wire N__6711;
    wire N__6710;
    wire N__6709;
    wire N__6702;
    wire N__6697;
    wire N__6692;
    wire N__6689;
    wire N__6686;
    wire N__6685;
    wire N__6682;
    wire N__6679;
    wire N__6674;
    wire N__6671;
    wire N__6668;
    wire N__6665;
    wire N__6664;
    wire N__6663;
    wire N__6662;
    wire N__6659;
    wire N__6656;
    wire N__6653;
    wire N__6650;
    wire N__6641;
    wire N__6640;
    wire N__6639;
    wire N__6638;
    wire N__6637;
    wire N__6634;
    wire N__6627;
    wire N__6624;
    wire N__6617;
    wire N__6616;
    wire N__6615;
    wire N__6612;
    wire N__6609;
    wire N__6606;
    wire N__6599;
    wire N__6598;
    wire N__6597;
    wire N__6596;
    wire N__6595;
    wire N__6592;
    wire N__6589;
    wire N__6584;
    wire N__6581;
    wire N__6572;
    wire N__6569;
    wire N__6566;
    wire N__6563;
    wire N__6560;
    wire N__6557;
    wire N__6554;
    wire N__6553;
    wire N__6550;
    wire N__6547;
    wire N__6542;
    wire N__6539;
    wire N__6536;
    wire N__6533;
    wire N__6530;
    wire N__6527;
    wire N__6524;
    wire N__6523;
    wire N__6522;
    wire N__6519;
    wire N__6516;
    wire N__6513;
    wire N__6510;
    wire N__6507;
    wire N__6504;
    wire N__6501;
    wire N__6498;
    wire N__6495;
    wire N__6490;
    wire N__6485;
    wire N__6482;
    wire N__6479;
    wire N__6476;
    wire N__6473;
    wire N__6470;
    wire N__6467;
    wire N__6464;
    wire N__6461;
    wire N__6458;
    wire N__6455;
    wire N__6452;
    wire N__6449;
    wire N__6446;
    wire N__6445;
    wire N__6442;
    wire N__6439;
    wire N__6436;
    wire N__6433;
    wire N__6430;
    wire N__6427;
    wire N__6424;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6412;
    wire N__6409;
    wire N__6404;
    wire N__6401;
    wire N__6398;
    wire N__6395;
    wire N__6392;
    wire N__6389;
    wire N__6386;
    wire N__6383;
    wire N__6380;
    wire N__6377;
    wire N__6374;
    wire N__6373;
    wire N__6370;
    wire N__6367;
    wire N__6364;
    wire N__6361;
    wire N__6358;
    wire N__6355;
    wire N__6350;
    wire N__6347;
    wire N__6344;
    wire N__6341;
    wire N__6338;
    wire N__6335;
    wire N__6332;
    wire N__6329;
    wire N__6326;
    wire N__6323;
    wire N__6320;
    wire N__6317;
    wire N__6314;
    wire N__6311;
    wire N__6308;
    wire N__6305;
    wire N__6302;
    wire N__6299;
    wire N__6298;
    wire N__6295;
    wire N__6292;
    wire N__6287;
    wire N__6284;
    wire N__6281;
    wire N__6278;
    wire N__6275;
    wire N__6274;
    wire N__6271;
    wire N__6268;
    wire N__6265;
    wire N__6262;
    wire N__6259;
    wire N__6256;
    wire N__6251;
    wire N__6248;
    wire N__6245;
    wire N__6242;
    wire N__6239;
    wire N__6238;
    wire N__6237;
    wire N__6236;
    wire N__6229;
    wire N__6228;
    wire N__6225;
    wire N__6222;
    wire N__6219;
    wire N__6212;
    wire N__6209;
    wire N__6208;
    wire N__6207;
    wire N__6206;
    wire N__6203;
    wire N__6198;
    wire N__6195;
    wire N__6188;
    wire N__6185;
    wire N__6184;
    wire N__6183;
    wire N__6182;
    wire N__6181;
    wire N__6180;
    wire N__6177;
    wire N__6174;
    wire N__6171;
    wire N__6164;
    wire N__6155;
    wire N__6154;
    wire N__6149;
    wire N__6146;
    wire N__6143;
    wire N__6140;
    wire N__6137;
    wire N__6134;
    wire N__6133;
    wire N__6130;
    wire N__6127;
    wire N__6122;
    wire N__6119;
    wire N__6116;
    wire N__6113;
    wire N__6110;
    wire N__6107;
    wire N__6104;
    wire N__6101;
    wire N__6098;
    wire N__6095;
    wire N__6092;
    wire N__6089;
    wire N__6088;
    wire N__6085;
    wire N__6084;
    wire N__6081;
    wire N__6078;
    wire N__6075;
    wire N__6072;
    wire N__6067;
    wire N__6064;
    wire N__6061;
    wire N__6058;
    wire N__6055;
    wire N__6052;
    wire N__6047;
    wire N__6046;
    wire N__6045;
    wire N__6040;
    wire N__6037;
    wire N__6032;
    wire N__6029;
    wire N__6026;
    wire N__6025;
    wire N__6020;
    wire N__6017;
    wire N__6014;
    wire N__6011;
    wire N__6010;
    wire N__6007;
    wire N__6004;
    wire N__5999;
    wire N__5996;
    wire N__5993;
    wire N__5990;
    wire N__5987;
    wire N__5984;
    wire N__5981;
    wire N__5978;
    wire N__5975;
    wire N__5972;
    wire N__5969;
    wire N__5966;
    wire N__5963;
    wire N__5960;
    wire N__5959;
    wire N__5956;
    wire N__5953;
    wire N__5950;
    wire N__5947;
    wire N__5944;
    wire N__5941;
    wire N__5938;
    wire N__5935;
    wire N__5932;
    wire N__5929;
    wire N__5926;
    wire N__5923;
    wire N__5920;
    wire N__5915;
    wire N__5912;
    wire N__5909;
    wire N__5906;
    wire N__5903;
    wire N__5900;
    wire N__5897;
    wire N__5894;
    wire N__5891;
    wire N__5888;
    wire N__5885;
    wire N__5882;
    wire N__5879;
    wire N__5876;
    wire N__5873;
    wire N__5870;
    wire N__5867;
    wire N__5864;
    wire N__5861;
    wire N__5858;
    wire N__5855;
    wire N__5852;
    wire N__5849;
    wire N__5846;
    wire N__5843;
    wire N__5840;
    wire N__5837;
    wire N__5834;
    wire N__5831;
    wire N__5828;
    wire N__5825;
    wire N__5822;
    wire N__5819;
    wire N__5816;
    wire N__5815;
    wire N__5812;
    wire N__5809;
    wire N__5806;
    wire N__5803;
    wire N__5800;
    wire N__5797;
    wire N__5794;
    wire N__5791;
    wire N__5786;
    wire N__5783;
    wire N__5780;
    wire N__5777;
    wire N__5774;
    wire N__5771;
    wire N__5768;
    wire N__5765;
    wire N__5762;
    wire N__5759;
    wire N__5756;
    wire N__5753;
    wire N__5750;
    wire N__5747;
    wire N__5744;
    wire N__5741;
    wire N__5738;
    wire N__5735;
    wire N__5732;
    wire N__5729;
    wire N__5728;
    wire N__5725;
    wire N__5722;
    wire N__5717;
    wire N__5714;
    wire N__5711;
    wire N__5708;
    wire N__5707;
    wire N__5704;
    wire N__5701;
    wire N__5698;
    wire N__5695;
    wire N__5690;
    wire N__5687;
    wire N__5684;
    wire N__5681;
    wire N__5678;
    wire N__5675;
    wire N__5672;
    wire N__5669;
    wire N__5666;
    wire N__5663;
    wire N__5660;
    wire N__5657;
    wire N__5654;
    wire N__5651;
    wire N__5648;
    wire N__5645;
    wire N__5642;
    wire N__5639;
    wire N__5636;
    wire N__5633;
    wire N__5630;
    wire N__5627;
    wire N__5624;
    wire N__5621;
    wire N__5618;
    wire N__5615;
    wire N__5612;
    wire N__5609;
    wire N__5606;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5594;
    wire N__5593;
    wire N__5590;
    wire N__5587;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5570;
    wire N__5567;
    wire N__5564;
    wire N__5561;
    wire N__5558;
    wire N__5557;
    wire N__5554;
    wire N__5551;
    wire N__5548;
    wire N__5545;
    wire N__5542;
    wire N__5539;
    wire N__5536;
    wire N__5533;
    wire N__5530;
    wire N__5527;
    wire N__5524;
    wire N__5519;
    wire N__5516;
    wire N__5513;
    wire N__5510;
    wire N__5507;
    wire N__5504;
    wire N__5501;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5489;
    wire N__5486;
    wire N__5483;
    wire N__5480;
    wire N__5477;
    wire N__5474;
    wire N__5471;
    wire N__5468;
    wire N__5465;
    wire N__5462;
    wire N__5459;
    wire N__5456;
    wire N__5455;
    wire N__5452;
    wire N__5449;
    wire N__5446;
    wire N__5443;
    wire N__5438;
    wire N__5435;
    wire N__5432;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5396;
    wire N__5395;
    wire N__5392;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5362;
    wire N__5359;
    wire N__5356;
    wire N__5353;
    wire N__5350;
    wire N__5345;
    wire N__5342;
    wire N__5339;
    wire N__5336;
    wire N__5333;
    wire N__5330;
    wire N__5327;
    wire N__5324;
    wire N__5321;
    wire N__5318;
    wire N__5315;
    wire N__5312;
    wire N__5309;
    wire N__5306;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5294;
    wire N__5291;
    wire N__5288;
    wire N__5285;
    wire N__5282;
    wire N__5279;
    wire N__5276;
    wire N__5273;
    wire N__5270;
    wire N__5267;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5255;
    wire N__5252;
    wire N__5249;
    wire N__5246;
    wire N__5243;
    wire N__5240;
    wire N__5239;
    wire N__5236;
    wire N__5233;
    wire N__5230;
    wire N__5227;
    wire N__5224;
    wire N__5221;
    wire N__5218;
    wire N__5215;
    wire N__5212;
    wire N__5209;
    wire N__5206;
    wire N__5203;
    wire N__5200;
    wire N__5195;
    wire N__5192;
    wire N__5189;
    wire N__5186;
    wire N__5183;
    wire N__5180;
    wire N__5177;
    wire N__5174;
    wire N__5171;
    wire N__5168;
    wire N__5165;
    wire N__5162;
    wire N__5159;
    wire N__5156;
    wire N__5153;
    wire N__5150;
    wire N__5147;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5135;
    wire N__5132;
    wire N__5129;
    wire N__5126;
    wire N__5123;
    wire N__5120;
    wire N__5117;
    wire N__5114;
    wire N__5111;
    wire N__5108;
    wire N__5105;
    wire N__5102;
    wire N__5099;
    wire N__5096;
    wire N__5093;
    wire N__5090;
    wire N__5087;
    wire N__5084;
    wire N__5081;
    wire N__5078;
    wire N__5075;
    wire N__5072;
    wire N__5069;
    wire N__5066;
    wire N__5063;
    wire N__5060;
    wire N__5057;
    wire N__5054;
    wire N__5053;
    wire N__5050;
    wire N__5047;
    wire N__5044;
    wire N__5041;
    wire N__5036;
    wire N__5033;
    wire N__5030;
    wire N__5027;
    wire N__5024;
    wire N__5021;
    wire N__5018;
    wire N__5015;
    wire N__5012;
    wire N__5009;
    wire N__5006;
    wire N__5003;
    wire N__5000;
    wire N__4997;
    wire N__4994;
    wire N__4991;
    wire N__4988;
    wire N__4985;
    wire N__4982;
    wire N__4979;
    wire N__4976;
    wire N__4973;
    wire N__4970;
    wire N__4967;
    wire N__4964;
    wire N__4961;
    wire N__4958;
    wire N__4955;
    wire N__4952;
    wire N__4949;
    wire N__4946;
    wire N__4943;
    wire N__4940;
    wire N__4937;
    wire N__4934;
    wire N__4931;
    wire N__4928;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4916;
    wire N__4913;
    wire N__4910;
    wire N__4907;
    wire N__4904;
    wire N__4901;
    wire N__4898;
    wire N__4895;
    wire N__4892;
    wire N__4891;
    wire N__4888;
    wire N__4885;
    wire N__4880;
    wire N__4877;
    wire N__4874;
    wire N__4871;
    wire N__4868;
    wire N__4865;
    wire N__4862;
    wire N__4859;
    wire N__4856;
    wire N__4853;
    wire N__4850;
    wire N__4847;
    wire N__4844;
    wire N__4841;
    wire N__4838;
    wire N__4835;
    wire N__4832;
    wire N__4829;
    wire N__4826;
    wire N__4823;
    wire N__4820;
    wire N__4817;
    wire N__4814;
    wire N__4811;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4799;
    wire N__4796;
    wire N__4793;
    wire N__4790;
    wire N__4787;
    wire N__4784;
    wire N__4781;
    wire N__4778;
    wire N__4775;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4748;
    wire N__4745;
    wire N__4742;
    wire N__4739;
    wire N__4736;
    wire N__4733;
    wire N__4730;
    wire N__4729;
    wire N__4726;
    wire N__4723;
    wire N__4720;
    wire N__4717;
    wire N__4714;
    wire N__4711;
    wire N__4708;
    wire N__4705;
    wire N__4702;
    wire N__4699;
    wire N__4696;
    wire N__4693;
    wire N__4690;
    wire N__4685;
    wire N__4682;
    wire N__4679;
    wire N__4676;
    wire N__4673;
    wire N__4670;
    wire N__4667;
    wire N__4664;
    wire N__4661;
    wire N__4658;
    wire N__4655;
    wire N__4652;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4640;
    wire N__4637;
    wire N__4634;
    wire N__4631;
    wire N__4628;
    wire N__4625;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4613;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4601;
    wire N__4598;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4586;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4565;
    wire N__4562;
    wire N__4559;
    wire N__4556;
    wire N__4553;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4541;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4523;
    wire N__4520;
    wire N__4517;
    wire N__4514;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4484;
    wire N__4481;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4463;
    wire N__4460;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4448;
    wire N__4445;
    wire N__4442;
    wire N__4439;
    wire N__4436;
    wire N__4433;
    wire N__4430;
    wire N__4427;
    wire N__4424;
    wire N__4421;
    wire N__4418;
    wire N__4415;
    wire N__4412;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4400;
    wire N__4397;
    wire N__4394;
    wire N__4391;
    wire N__4388;
    wire N__4385;
    wire N__4382;
    wire N__4379;
    wire N__4376;
    wire N__4373;
    wire N__4370;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4346;
    wire N__4343;
    wire N__4340;
    wire N__4337;
    wire N__4334;
    wire N__4331;
    wire N__4328;
    wire N__4325;
    wire N__4322;
    wire N__4319;
    wire N__4316;
    wire N__4313;
    wire N__4310;
    wire N__4307;
    wire N__4304;
    wire N__4301;
    wire N__4298;
    wire N__4295;
    wire N__4292;
    wire N__4289;
    wire N__4286;
    wire N__4283;
    wire N__4280;
    wire N__4277;
    wire N__4274;
    wire N__4271;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4256;
    wire N__4253;
    wire N__4250;
    wire N__4247;
    wire N__4244;
    wire N__4241;
    wire N__4238;
    wire N__4235;
    wire N__4232;
    wire N__4229;
    wire N__4226;
    wire N__4223;
    wire N__4220;
    wire N__4217;
    wire N__4214;
    wire N__4211;
    wire N__4208;
    wire N__4205;
    wire N__4202;
    wire N__4199;
    wire N__4196;
    wire N__4193;
    wire N__4190;
    wire N__4187;
    wire N__4184;
    wire N__4181;
    wire N__4178;
    wire N__4175;
    wire N__4172;
    wire N__4169;
    wire N__4166;
    wire N__4163;
    wire N__4160;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4148;
    wire N__4145;
    wire N__4142;
    wire N__4139;
    wire N__4136;
    wire N__4133;
    wire N__4130;
    wire N__4127;
    wire N__4124;
    wire N__4121;
    wire N__4118;
    wire N__4115;
    wire N__4112;
    wire N__4109;
    wire N__4106;
    wire N__4103;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4088;
    wire N__4085;
    wire N__4082;
    wire N__4079;
    wire N__4076;
    wire N__4073;
    wire N__4070;
    wire N__4067;
    wire N__4064;
    wire N__4061;
    wire N__4058;
    wire N__4055;
    wire N__4052;
    wire N__4049;
    wire N__4046;
    wire N__4043;
    wire N__4040;
    wire N__4037;
    wire TCIn_c;
    wire VCCG0;
    wire GNDG0;
    wire TAn_in;
    wire N_240_i;
    wire N_237_i;
    wire N_239_i;
    wire WRITE_CYCLE_ACTIVE_rep26_i_ess;
    wire N_238_i;
    wire WRITE_CYCLE_ACTIVE_rep24_i_ess;
    wire N_242_i;
    wire N_243_i;
    wire N_229_i;
    wire N_244_i;
    wire WRITE_CYCLE_ACTIVE_rep29_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep17_i_ess;
    wire N_230_i;
    wire RESETn_c_i;
    wire \U111_CYCLE_SM.CYCLE_STATE_0_0 ;
    wire N_221_i;
    wire N_223_i;
    wire N_233_i;
    wire WRITE_CYCLE_ACTIVE_rep10_i_ess;
    wire N_234_i;
    wire WRITE_CYCLE_ACTIVE_rep9_i_ess;
    wire N_222_i;
    wire N_236_i;
    wire N_235_i;
    wire N_224_i;
    wire N_227_i;
    wire N_214_i;
    wire N_228_i;
    wire N_225_i;
    wire WRITE_CYCLE_ACTIVE_rep15_i_ess;
    wire N_241_i;
    wire WRITE_CYCLE_ACTIVE_rep25_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep30_i_ess;
    wire WRITE_CYCLE_ACTIVE_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep16_i_ess;
    wire N_232_i;
    wire WRITE_CYCLE_ACTIVE_rep8_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep20_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep11_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep22_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep14_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep1_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep12_i_ess;
    wire N_216_i;
    wire WRITE_CYCLE_ACTIVE_rep5_i_ess;
    wire N_218_i;
    wire A_040_c_0;
    wire A_AMIGA_c_0;
    wire U111_CYCLE_SM_A_AMIGA_0_i_1;
    wire WRITE_CYCLE_ACTIVE_rep28_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep27_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep19_i_ess;
    wire N_231_i;
    wire WRITE_CYCLE_ACTIVE_rep18_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep21_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep23_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep7_i_ess;
    wire N_220_i;
    wire WRITE_CYCLE_ACTIVE_rep3_i_ess;
    wire N_219_i;
    wire D_LL_AMIGA_in_0;
    wire un2_D_LL_AMIGA_0;
    wire D_LM_AMIGA_in_1;
    wire un2_D_LM_AMIGA_1;
    wire D_UM_040_in_2;
    wire D_LL_040_in_2;
    wire un1_D_UM_040_2;
    wire D_UM_040_in_6;
    wire D_LL_040_in_6;
    wire un1_D_UM_040_6;
    wire D_LM_AMIGA_in_2;
    wire un2_D_LM_AMIGA_2;
    wire WRITE_CYCLE_ACTIVE_rep0_i_ess;
    wire N_213_i;
    wire N_226_i;
    wire WRITE_CYCLE_ACTIVE_rep6_i_ess;
    wire D_LL_AMIGA_in_1;
    wire un2_D_LL_AMIGA_1;
    wire A_040_c_1;
    wire WRITE_CYCLE_ACTIVE_rep13_i_ess;
    wire WRITE_CYCLE_ACTIVE_rep4_i_ess;
    wire N_217_i;
    wire D_LL_AMIGA_in_4;
    wire un2_D_LL_AMIGA_4;
    wire D_LL_040_in_0;
    wire D_UM_040_in_0;
    wire un1_D_UM_040_0;
    wire D_LM_AMIGA_in_3;
    wire un2_D_LM_AMIGA_3;
    wire LBENn_c_i;
    wire WRITE_CYCLE_ACTIVE_rep2_i_ess;
    wire N_215_i;
    wire CONSTANT_ONE_NET;
    wire D_LL_AMIGA_in_2;
    wire un2_D_LL_AMIGA_2;
    wire D_LM_AMIGA_in_0;
    wire un2_D_LM_AMIGA_0;
    wire TSn_c;
    wire \INVU111_CYCLE_SM.TSnC_net ;
    wire \U111_CYCLE_SM.TS_ENZ0 ;
    wire D_UM_040_in_1;
    wire D_LL_040_in_1;
    wire un1_D_UM_040_1;
    wire D_LM_AMIGA_in_6;
    wire un2_D_LM_AMIGA_6;
    wire D_LM_040_in_1;
    wire D_UU_040_in_1;
    wire un1_D_UU_040_1;
    wire D_LL_040_in_5;
    wire D_UM_040_in_5;
    wire un1_D_UM_040_5;
    wire D_UU_040_in_6;
    wire D_LM_040_in_6;
    wire un1_D_UU_040_6;
    wire D_LL_AMIGA_in_3;
    wire un2_D_LL_AMIGA_3;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa_cascade_ ;
    wire \U111_CYCLE_SM.un1_CYCLE_STATE_0 ;
    wire \U111_CYCLE_SM.TS_EN_6 ;
    wire SIZ_c_1;
    wire SIZ_c_0;
    wire \U111_CYCLE_SM.FLIP_WORD_2 ;
    wire PORTSIZE_c;
    wire \U111_CYCLE_SM.LW_TRANSZ0 ;
    wire \U111_CYCLE_SM.PORT_MISMATCH_2 ;
    wire \U111_CYCLE_SM.A2_ENZ0 ;
    wire D_LM_AMIGA_in_5;
    wire un2_D_LM_AMIGA_5;
    wire D_LM_040_in_0;
    wire D_UU_040_in_0;
    wire un1_D_UU_040_0;
    wire D_LL_AMIGA_in_6;
    wire un2_D_LL_AMIGA_6;
    wire \U111_CYCLE_SM.N_124_0 ;
    wire \U111_CYCLE_SM.N_132_cascade_ ;
    wire \U111_CYCLE_SM.BURST_COUNTZ0Z_1 ;
    wire TBIn_c;
    wire \U111_CYCLE_SM.un7_CYCLE_STATE_0 ;
    wire \U111_CYCLE_SM.un7_CYCLE_STATE_0_cascade_ ;
    wire \U111_CYCLE_SM.CYCLE_STATE_srsts_i_1_2_cascade_ ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ;
    wire \U111_CYCLE_SM.PORT_MISMATCHZ0 ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ;
    wire \U111_CYCLE_SM.BURST_COUNTZ0Z_0 ;
    wire \U111_CYCLE_SM.BURSTZ0 ;
    wire \U111_CYCLE_SM.N_131_cascade_ ;
    wire \U111_CYCLE_SM.CYCLE_STATE_srsts_0_1_0 ;
    wire \U111_CYCLE_SM.TS_EN6 ;
    wire \U111_CYCLE_SM.N_144 ;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ;
    wire D_UU_AMIGA_in_1;
    wire un1_D_UU_AMIGA_1;
    wire D_UM_040_in_3;
    wire D_LL_040_in_3;
    wire un1_D_UM_040_3;
    wire D_LM_040_in_3;
    wire D_UU_040_in_3;
    wire un1_D_UU_040_3;
    wire LBENn_c_i_0;
    wire D_LL_AMIGA_in_7;
    wire un2_D_LL_AMIGA_7;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ;
    wire \U111_CYCLE_SM.N_119_0 ;
    wire \U111_CYCLE_SM.N_117_0 ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ;
    wire \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_cascade_ ;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1_cascade_ ;
    wire \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa ;
    wire TACKn_in;
    wire TEAn_c;
    wire RESETn_c;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ;
    wire \U111_CYCLE_SM.CYCLE_STATE_srsts_i_o2_0_5_cascade_ ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ;
    wire \U111_CYCLE_SM.TA_DISZ0 ;
    wire TAn_1_i;
    wire D_LM_AMIGA_in_4;
    wire un2_D_LM_AMIGA_4;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ;
    wire D_UU_AMIGA_in_5;
    wire un1_D_UU_AMIGA_5;
    wire D_UM_AMIGA_in_1;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ;
    wire un1_D_UM_AMIGA_1;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ;
    wire D_UU_AMIGA_in_0;
    wire un1_D_UU_AMIGA_0;
    wire D_LL_AMIGA_in_5;
    wire un2_D_LL_AMIGA_5;
    wire \U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0 ;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1 ;
    wire CLK80;
    wire GB_BUFFER_CLK80_THRU_CO;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ;
    wire D_UU_AMIGA_in_2;
    wire un1_D_UU_AMIGA_2;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ;
    wire un1_D_UU_AMIGA_7;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ;
    wire D_UU_AMIGA_in_4;
    wire un1_D_UU_AMIGA_4;
    wire D_UM_AMIGA_in_3;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ;
    wire un1_D_UM_AMIGA_3;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ;
    wire D_UM_AMIGA_in_4;
    wire un1_D_UM_AMIGA_4;
    wire D_LM_AMIGA_in_7;
    wire D_UU_AMIGA_in_7;
    wire un2_D_LM_AMIGA_7;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ;
    wire D_UM_AMIGA_in_7;
    wire un1_D_UM_AMIGA_7;
    wire D_UM_AMIGA_in_5;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ;
    wire un1_D_UM_AMIGA_5;
    wire D_UU_040_in_2;
    wire D_LM_040_in_2;
    wire un1_D_UU_040_2;
    wire D_UU_040_in_5;
    wire D_LM_040_in_5;
    wire un1_D_UU_040_5;
    wire D_UU_AMIGA_in_3;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ;
    wire un1_D_UU_AMIGA_3;
    wire D_UU_AMIGA_in_6;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ;
    wire un1_D_UU_AMIGA_6;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ;
    wire D_UM_AMIGA_in_2;
    wire un1_D_UM_AMIGA_2;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ;
    wire D_UM_AMIGA_in_6;
    wire un1_D_UM_AMIGA_6;
    wire D_LL_040_in_4;
    wire D_UM_040_in_4;
    wire un1_D_UM_040_4;
    wire D_UU_040_in_4;
    wire D_LM_040_in_4;
    wire un1_D_UU_040_4;
    wire \U111_CYCLE_SM.LATCH_ENZ0 ;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ;
    wire D_UM_AMIGA_in_0;
    wire un1_D_UM_AMIGA_0;
    wire D_UM_040_in_7;
    wire D_LL_040_in_7;
    wire un1_D_UM_040_7;
    wire \U111_CYCLE_SM.FLIP_WORDZ0 ;
    wire D_UU_040_in_7;
    wire D_LM_040_in_7;
    wire un1_D_UU_040_7;
    wire READ_CYCLE_ACTIVE_rep4_i_ess;
    wire N_185_i;
    wire READ_CYCLE_ACTIVE_rep2_i_ess;
    wire N_183_i;
    wire READ_CYCLE_ACTIVE_rep0_i_ess;
    wire N_181_i;
    wire READ_CYCLE_ACTIVE_rep7_i_ess;
    wire N_188_i;
    wire N_209_i;
    wire READ_CYCLE_ACTIVE_rep28_i_ess;
    wire GB_BUFFER_CLK40_THRU_CO;
    wire READ_CYCLE_ACTIVE_rep5_i_ess;
    wire N_186_i;
    wire READ_CYCLE_ACTIVE_rep6_i_ess;
    wire N_187_i;
    wire N_193_i;
    wire N_194_i;
    wire N_205_i;
    wire N_206_i;
    wire N_208_i;
    wire READ_CYCLE_ACTIVE_rep25_i_ess;
    wire READ_CYCLE_ACTIVE_rep24_i_ess;
    wire READ_CYCLE_ACTIVE_rep27_i_ess;
    wire N_211_i;
    wire READ_CYCLE_ACTIVE_rep26_i_ess;
    wire N_207_i;
    wire READ_CYCLE_ACTIVE_rep30_i_ess;
    wire READ_CYCLE_ACTIVE_rep17_i_ess;
    wire N_198_i;
    wire READ_CYCLE_ACTIVE_rep18_i_ess;
    wire N_199_i;
    wire READ_CYCLE_ACTIVE_rep31_i_ess;
    wire N_212_i;
    wire N_197_i;
    wire N_200_i;
    wire READ_CYCLE_ACTIVE_rep19_i_ess;
    wire READ_CYCLE_ACTIVE_rep16_i_ess;
    wire READ_CYCLE_ACTIVE_rep20_i_ess;
    wire N_201_i;
    wire READ_CYCLE_ACTIVE_rep8_i_ess;
    wire N_189_i;
    wire READ_CYCLE_ACTIVE_rep21_i_ess;
    wire N_202_i;
    wire N_210_i;
    wire N_191_i;
    wire READ_CYCLE_ACTIVE_rep10_i_ess;
    wire READ_CYCLE_ACTIVE_rep29_i_ess;
    wire N_195_i;
    wire READ_CYCLE_ACTIVE_rep14_i_ess;
    wire READ_CYCLE_ACTIVE_rep22_i_ess;
    wire N_203_i;
    wire READ_CYCLE_ACTIVE_rep23_i_ess;
    wire N_204_i;
    wire READ_CYCLE_ACTIVE_rep9_i_ess;
    wire N_190_i;
    wire READ_CYCLE_ACTIVE_rep11_i_ess;
    wire N_192_i;
    wire READ_CYCLE_ACTIVE_rep3_i_ess;
    wire N_184_i;
    wire READ_CYCLE_ACTIVE_rep15_i_ess;
    wire N_196_i;
    wire READ_CYCLE_ACTIVE_rep1_i_ess;
    wire N_182_i;
    wire READ_CYCLE_ACTIVE_rep13_i_ess;
    wire BGn_c;
    wire TS_CPUn_c;
    wire LBENn_c;
    wire RnW_c;
    wire READ_CYCLE_ACTIVE_rep12_i_ess;
    wire _gnd_net_;
    wire CLK40;
    wire \U111_CYCLE_SM.CYCLE_STATE_0_g_0 ;
    wire RESETn_c_i_g;

    defparam pll_pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll_pll.TEST_MODE=1'b0;
    defparam pll_pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll_pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll_pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll_pll.FILTER_RANGE=3'b011;
    defparam pll_pll.FEEDBACK_PATH="SIMPLE";
    defparam pll_pll.FDA_RELATIVE=4'b0000;
    defparam pll_pll.FDA_FEEDBACK=4'b0000;
    defparam pll_pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll_pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll_pll.DIVR=4'b0000;
    defparam pll_pll.DIVQ=3'b011;
    defparam pll_pll.DIVF=7'b0001111;
    defparam pll_pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40_2F pll_pll (
            .SCLK(),
            .PLLOUTGLOBALA(CLK80),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALB(CLK40),
            .SDI(),
            .PLLOUTCOREA(),
            .BYPASS(),
            .RESETB(N__5708),
            .PLLOUTCOREB(),
            .LOCK(),
            .SDO(),
            .EXTFEEDBACK(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__13729));
    IO_PAD pll_iopad (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__13729),
            .PACKAGEPIN(CLK40_IN));
    IO_PAD LBENn_ibuf_iopad (
            .OE(N__13713),
            .DIN(N__13712),
            .DOUT(N__13711),
            .PACKAGEPIN(LBENn));
    defparam LBENn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam LBENn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO LBENn_ibuf_preio (
            .PADOEN(N__13713),
            .PADOUT(N__13712),
            .PADIN(N__13711),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(LBENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TAn_iobuf_iopad (
            .OE(N__13704),
            .DIN(N__13703),
            .DOUT(N__13702),
            .PACKAGEPIN(TAn));
    defparam TAn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TAn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TAn_iobuf_preio (
            .PADOEN(N__13704),
            .PADOUT(N__13703),
            .PADIN(N__13702),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7106),
            .DIN0(TAn_in),
            .DOUT0(N__7418),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_1_iopad (
            .OE(N__13695),
            .DIN(N__13694),
            .DOUT(N__13693),
            .PACKAGEPIN(D_LL_AMIGA[1]));
    defparam D_LL_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_1_preio (
            .PADOEN(N__13695),
            .PADOUT(N__13694),
            .PADIN(N__13693),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4103),
            .DIN0(D_LL_AMIGA_in_1),
            .DOUT0(N__5561),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_6_iopad (
            .OE(N__13686),
            .DIN(N__13685),
            .DOUT(N__13684),
            .PACKAGEPIN(D_UU_040[6]));
    defparam D_UU_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_6_preio (
            .PADOEN(N__13686),
            .PADOUT(N__13685),
            .PADIN(N__13684),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9524),
            .DIN0(D_UU_040_in_6),
            .DOUT0(N__7886),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam CPUBGn_obuf_iopad.PULLUP=1'b1;
    IO_PAD CPUBGn_obuf_iopad (
            .OE(N__13677),
            .DIN(N__13676),
            .DOUT(N__13675),
            .PACKAGEPIN(CPUBGn));
    defparam CPUBGn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CPUBGn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CPUBGn_obuf_preio (
            .PADOEN(N__13677),
            .PADOUT(N__13676),
            .PADIN(N__13675),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_3_iopad (
            .OE(N__13668),
            .DIN(N__13667),
            .DOUT(N__13666),
            .PACKAGEPIN(D_UM_AMIGA[3]));
    defparam D_UM_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_3_preio (
            .PADOEN(N__13668),
            .PADOUT(N__13667),
            .PADIN(N__13666),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4310),
            .DIN0(D_UM_AMIGA_in_3),
            .DOUT0(N__6401),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_040_ibuf_1_iopad.PULLUP=1'b1;
    IO_PAD A_040_ibuf_1_iopad (
            .OE(N__13659),
            .DIN(N__13658),
            .DOUT(N__13657),
            .PACKAGEPIN(A_040[1]));
    defparam A_040_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_040_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_040_ibuf_1_preio (
            .PADOEN(N__13659),
            .PADOUT(N__13658),
            .PADIN(N__13657),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_040_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_4_iopad (
            .OE(N__13650),
            .DIN(N__13649),
            .DOUT(N__13648),
            .PACKAGEPIN(D_LM_AMIGA[4]));
    defparam D_LM_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_4_preio (
            .PADOEN(N__13650),
            .PADOUT(N__13649),
            .PADIN(N__13648),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4394),
            .DIN0(D_LM_AMIGA_in_4),
            .DOUT0(N__9164),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_7_iopad (
            .OE(N__13641),
            .DIN(N__13640),
            .DOUT(N__13639),
            .PACKAGEPIN(D_LM_040[7]));
    defparam D_LM_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_7_preio (
            .PADOEN(N__13641),
            .PADOUT(N__13640),
            .PADIN(N__13639),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9971),
            .DIN0(D_LM_040_in_7),
            .DOUT0(N__8339),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_obuf_iopad (
            .OE(N__13632),
            .DIN(N__13631),
            .DOUT(N__13630),
            .PACKAGEPIN(CLK40B));
    defparam CLK40B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_obuf_preio (
            .PADOEN(N__13632),
            .PADOUT(N__13631),
            .PADIN(N__13630),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9617),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_1_iopad (
            .OE(N__13623),
            .DIN(N__13622),
            .DOUT(N__13621),
            .PACKAGEPIN(D_UM_040[1]));
    defparam D_UM_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_1_preio (
            .PADOEN(N__13623),
            .PADOUT(N__13622),
            .PADIN(N__13621),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9950),
            .DIN0(D_UM_040_in_1),
            .DOUT0(N__6917),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_ibuf_iopad (
            .OE(N__13614),
            .DIN(N__13613),
            .DOUT(N__13612),
            .PACKAGEPIN(TBIn));
    defparam TBIn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TBIn_ibuf_preio (
            .PADOEN(N__13614),
            .PADOUT(N__13613),
            .PADIN(N__13612),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TBIn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_7_iopad (
            .OE(N__13605),
            .DIN(N__13604),
            .DOUT(N__13603),
            .PACKAGEPIN(D_UU_AMIGA[7]));
    defparam D_UU_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_7_preio (
            .PADOEN(N__13605),
            .PADOUT(N__13604),
            .PADIN(N__13603),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4847),
            .DIN0(D_UU_AMIGA_in_7),
            .DOUT0(N__8498),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFDIR_obuf_iopad (
            .OE(N__13596),
            .DIN(N__13595),
            .DOUT(N__13594),
            .PACKAGEPIN(BUFDIR));
    defparam BUFDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFDIR_obuf_preio (
            .PADOEN(N__13596),
            .PADOUT(N__13595),
            .PADIN(N__13594),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10580),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__13587),
            .DIN(N__13586),
            .DOUT(N__13585),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__13587),
            .PADOUT(N__13586),
            .PADIN(N__13585),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TS_CPUn_ibuf_iopad (
            .OE(N__13578),
            .DIN(N__13577),
            .DOUT(N__13576),
            .PACKAGEPIN(TS_CPUn));
    defparam TS_CPUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TS_CPUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TS_CPUn_ibuf_preio (
            .PADOEN(N__13578),
            .PADOUT(N__13577),
            .PADIN(N__13576),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TS_CPUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_1_iopad (
            .OE(N__13569),
            .DIN(N__13568),
            .DOUT(N__13567),
            .PACKAGEPIN(D_LL_040[1]));
    defparam D_LL_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_1_preio (
            .PADOEN(N__13569),
            .PADOUT(N__13568),
            .PADIN(N__13567),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9680),
            .DIN0(D_LL_040_in_1),
            .DOUT0(N__4922),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_1_iopad (
            .OE(N__13560),
            .DIN(N__13559),
            .DOUT(N__13558),
            .PACKAGEPIN(D_UU_040[1]));
    defparam D_UU_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_1_preio (
            .PADOEN(N__13560),
            .PADOUT(N__13559),
            .PADIN(N__13558),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__12278),
            .DIN0(D_UU_040_in_1),
            .DOUT0(N__6482),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_1_iopad (
            .OE(N__13551),
            .DIN(N__13550),
            .DOUT(N__13549),
            .PACKAGEPIN(D_LM_AMIGA[1]));
    defparam D_LM_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_1_preio (
            .PADOEN(N__13551),
            .PADOUT(N__13550),
            .PADIN(N__13549),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4226),
            .DIN0(D_LM_AMIGA_in_1),
            .DOUT0(N__5465),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_2_iopad (
            .OE(N__13542),
            .DIN(N__13541),
            .DOUT(N__13540),
            .PACKAGEPIN(D_LM_040[2]));
    defparam D_LM_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_2_preio (
            .PADOEN(N__13542),
            .PADOUT(N__13541),
            .PADIN(N__13540),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9791),
            .DIN0(D_LM_040_in_2),
            .DOUT0(N__5000),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TACKn_iobuf_iopad.PULLUP=1'b1;
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__13533),
            .DIN(N__13532),
            .DOUT(N__13531),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__13533),
            .PADOUT(N__13532),
            .PADIN(N__13531),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6818),
            .DIN0(TACKn_in),
            .DOUT0(N__4178),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_2_iopad (
            .OE(N__13524),
            .DIN(N__13523),
            .DOUT(N__13522),
            .PACKAGEPIN(D_UM_040[2]));
    defparam D_UM_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_2_preio (
            .PADOEN(N__13524),
            .PADOUT(N__13523),
            .PADIN(N__13522),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9860),
            .DIN0(D_UM_040_in_2),
            .DOUT0(N__9350),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAMB_obuf_iopad (
            .OE(N__13515),
            .DIN(N__13514),
            .DOUT(N__13513),
            .PACKAGEPIN(CLKRAMB));
    defparam CLKRAMB_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAMB_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAMB_obuf_preio (
            .PADOEN(N__13515),
            .PADOUT(N__13514),
            .PADIN(N__13513),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7751),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_2_iopad (
            .OE(N__13506),
            .DIN(N__13505),
            .DOUT(N__13504),
            .PACKAGEPIN(D_LL_AMIGA[2]));
    defparam D_LL_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_2_preio (
            .PADOEN(N__13506),
            .PADOUT(N__13505),
            .PADIN(N__13504),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4124),
            .DIN0(D_LL_AMIGA_in_2),
            .DOUT0(N__4730),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_2_iopad (
            .OE(N__13497),
            .DIN(N__13496),
            .DOUT(N__13495),
            .PACKAGEPIN(D_UU_AMIGA[2]));
    defparam D_UU_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_2_preio (
            .PADOEN(N__13497),
            .PADOUT(N__13496),
            .PADIN(N__13495),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5099),
            .DIN0(D_UU_AMIGA_in_2),
            .DOUT0(N__8117),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TEAn_ibuf_iopad.PULLUP=1'b1;
    IO_PAD TEAn_ibuf_iopad (
            .OE(N__13488),
            .DIN(N__13487),
            .DOUT(N__13486),
            .PACKAGEPIN(TEAn));
    defparam TEAn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TEAn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TEAn_ibuf_preio (
            .PADOEN(N__13488),
            .PADOUT(N__13487),
            .PADIN(N__13486),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TEAn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__13479),
            .DIN(N__13478),
            .DOUT(N__13477),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__13479),
            .PADOUT(N__13478),
            .PADIN(N__13477),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5123),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMAn_obuf_iopad (
            .OE(N__13470),
            .DIN(N__13469),
            .DOUT(N__13468),
            .PACKAGEPIN(DMAn));
    defparam DMAn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMAn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMAn_obuf_preio (
            .PADOEN(N__13470),
            .PADOUT(N__13469),
            .PADIN(N__13468),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5707),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_6_iopad (
            .OE(N__13461),
            .DIN(N__13460),
            .DOUT(N__13459),
            .PACKAGEPIN(D_LL_040[6]));
    defparam D_LL_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_6_preio (
            .PADOEN(N__13461),
            .PADOUT(N__13460),
            .PADIN(N__13459),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9632),
            .DIN0(D_LL_040_in_6),
            .DOUT0(N__5864),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_5_iopad (
            .OE(N__13452),
            .DIN(N__13451),
            .DOUT(N__13450),
            .PACKAGEPIN(D_LL_AMIGA[5]));
    defparam D_LL_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_5_preio (
            .PADOEN(N__13452),
            .PADOUT(N__13451),
            .PADIN(N__13450),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4079),
            .DIN0(D_LL_AMIGA_in_5),
            .DOUT0(N__5396),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_0_iopad (
            .OE(N__13443),
            .DIN(N__13442),
            .DOUT(N__13441),
            .PACKAGEPIN(D_UM_AMIGA[0]));
    defparam D_UM_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_0_preio (
            .PADOEN(N__13443),
            .PADOUT(N__13442),
            .PADIN(N__13441),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4187),
            .DIN0(D_UM_AMIGA_in_0),
            .DOUT0(N__5180),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_2_iopad (
            .OE(N__13434),
            .DIN(N__13433),
            .DOUT(N__13432),
            .PACKAGEPIN(D_UU_040[2]));
    defparam D_UU_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_2_preio (
            .PADOEN(N__13434),
            .PADOUT(N__13433),
            .PADIN(N__13432),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9482),
            .DIN0(D_UU_040_in_2),
            .DOUT0(N__7661),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_2_iopad (
            .OE(N__13425),
            .DIN(N__13424),
            .DOUT(N__13423),
            .PACKAGEPIN(D_LM_AMIGA[2]));
    defparam D_LM_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_2_preio (
            .PADOEN(N__13425),
            .PADOUT(N__13424),
            .PADIN(N__13423),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4565),
            .DIN0(D_LM_AMIGA_in_2),
            .DOUT0(N__8155),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK80_CPU_obuf_iopad (
            .OE(N__13416),
            .DIN(N__13415),
            .DOUT(N__13414),
            .PACKAGEPIN(CLK80_CPU));
    defparam CLK80_CPU_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK80_CPU_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK80_CPU_obuf_preio (
            .PADOEN(N__13416),
            .PADOUT(N__13415),
            .PADIN(N__13414),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7750),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_3_iopad (
            .OE(N__13407),
            .DIN(N__13406),
            .DOUT(N__13405),
            .PACKAGEPIN(D_LL_040[3]));
    defparam D_LL_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_3_preio (
            .PADOEN(N__13407),
            .PADOUT(N__13406),
            .PADIN(N__13405),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9665),
            .DIN0(D_LL_040_in_3),
            .DOUT0(N__5747),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_1_iopad (
            .OE(N__13398),
            .DIN(N__13397),
            .DOUT(N__13396),
            .PACKAGEPIN(D_LM_040[1]));
    defparam D_LM_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_1_preio (
            .PADOEN(N__13398),
            .PADOUT(N__13397),
            .PADIN(N__13396),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9812),
            .DIN0(D_LM_040_in_1),
            .DOUT0(N__4769),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_obuf_iopad (
            .OE(N__13389),
            .DIN(N__13388),
            .DOUT(N__13387),
            .PACKAGEPIN(TSn));
    defparam TSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TSn_obuf_preio (
            .PADOEN(N__13389),
            .PADOUT(N__13388),
            .PADIN(N__13387),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5606),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_7_iopad (
            .OE(N__13380),
            .DIN(N__13379),
            .DOUT(N__13378),
            .PACKAGEPIN(D_UM_AMIGA[7]));
    defparam D_UM_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_7_preio (
            .PADOEN(N__13380),
            .PADOUT(N__13379),
            .PADIN(N__13378),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4484),
            .DIN0(D_UM_AMIGA_in_7),
            .DOUT0(N__8843),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_7_iopad (
            .OE(N__13371),
            .DIN(N__13370),
            .DOUT(N__13369),
            .PACKAGEPIN(D_LM_AMIGA[7]));
    defparam D_LM_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_7_preio (
            .PADOEN(N__13371),
            .PADOUT(N__13370),
            .PADIN(N__13369),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4340),
            .DIN0(D_LM_AMIGA_in_7),
            .DOUT0(N__8537),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PORTSIZE_ibuf_iopad (
            .OE(N__13362),
            .DIN(N__13361),
            .DOUT(N__13360),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO PORTSIZE_ibuf_preio (
            .PADOEN(N__13362),
            .PADOUT(N__13361),
            .PADIN(N__13360),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(PORTSIZE_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_AMIGA_obuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_AMIGA_obuf_0_iopad (
            .OE(N__13353),
            .DIN(N__13352),
            .DOUT(N__13351),
            .PACKAGEPIN(A_AMIGA[0]));
    defparam A_AMIGA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_AMIGA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO A_AMIGA_obuf_0_preio (
            .PADOEN(N__13353),
            .PADOUT(N__13352),
            .PADIN(N__13351),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4613),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_4_iopad (
            .OE(N__13344),
            .DIN(N__13343),
            .DOUT(N__13342),
            .PACKAGEPIN(D_LM_040[4]));
    defparam D_LM_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_4_preio (
            .PADOEN(N__13344),
            .PADOUT(N__13343),
            .PADIN(N__13342),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9923),
            .DIN0(D_LM_040_in_4),
            .DOUT0(N__7067),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_7_iopad (
            .OE(N__13335),
            .DIN(N__13334),
            .DOUT(N__13333),
            .PACKAGEPIN(D_UM_040[7]));
    defparam D_UM_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_7_preio (
            .PADOEN(N__13335),
            .PADOUT(N__13334),
            .PADIN(N__13333),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__12299),
            .DIN0(D_UM_040_in_7),
            .DOUT0(N__8276),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__13326),
            .DIN(N__13325),
            .DOUT(N__13324),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__13326),
            .PADOUT(N__13325),
            .PADIN(N__13324),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_1_iopad (
            .OE(N__13317),
            .DIN(N__13316),
            .DOUT(N__13315),
            .PACKAGEPIN(D_UU_AMIGA[1]));
    defparam D_UU_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_1_preio (
            .PADOEN(N__13317),
            .PADOUT(N__13316),
            .PADIN(N__13315),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4499),
            .DIN0(D_UU_AMIGA_in_1),
            .DOUT0(N__5414),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_obuf_iopad (
            .OE(N__13308),
            .DIN(N__13307),
            .DOUT(N__13306),
            .PACKAGEPIN(CLK40C));
    defparam CLK40C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_obuf_preio (
            .PADOEN(N__13308),
            .PADOUT(N__13307),
            .PADIN(N__13306),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9616),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_0_iopad (
            .OE(N__13299),
            .DIN(N__13298),
            .DOUT(N__13297),
            .PACKAGEPIN(D_UM_040[0]));
    defparam D_UM_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_0_preio (
            .PADOEN(N__13299),
            .PADOUT(N__13298),
            .PADIN(N__13297),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9905),
            .DIN0(D_UM_040_in_0),
            .DOUT0(N__8927),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_0_iopad (
            .OE(N__13290),
            .DIN(N__13289),
            .DOUT(N__13288),
            .PACKAGEPIN(D_LL_AMIGA[0]));
    defparam D_LL_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_0_preio (
            .PADOEN(N__13290),
            .PADOUT(N__13289),
            .PADIN(N__13288),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4139),
            .DIN0(D_LL_AMIGA_in_0),
            .DOUT0(N__5240),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_4_iopad (
            .OE(N__13281),
            .DIN(N__13280),
            .DOUT(N__13279),
            .PACKAGEPIN(D_UU_AMIGA[4]));
    defparam D_UU_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_4_preio (
            .PADOEN(N__13281),
            .PADOUT(N__13280),
            .PADIN(N__13279),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5291),
            .DIN0(D_UU_AMIGA_in_4),
            .DOUT0(N__9128),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_7_iopad (
            .OE(N__13272),
            .DIN(N__13271),
            .DOUT(N__13270),
            .PACKAGEPIN(D_UU_040[7]));
    defparam D_UU_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_7_preio (
            .PADOEN(N__13272),
            .PADOUT(N__13271),
            .PADIN(N__13270),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9437),
            .DIN0(D_UU_040_in_7),
            .DOUT0(N__7631),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__13263),
            .DIN(N__13262),
            .DOUT(N__13261),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__13263),
            .PADOUT(N__13262),
            .PADIN(N__13261),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam BGn_ibuf_iopad.PULLUP=1'b1;
    IO_PAD BGn_ibuf_iopad (
            .OE(N__13254),
            .DIN(N__13253),
            .DOUT(N__13252),
            .PACKAGEPIN(BGn));
    defparam BGn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam BGn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO BGn_ibuf_preio (
            .PADOEN(N__13254),
            .PADOUT(N__13253),
            .PADIN(N__13252),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(BGn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_0_iopad (
            .OE(N__13245),
            .DIN(N__13244),
            .DOUT(N__13243),
            .PACKAGEPIN(D_LL_040[0]));
    defparam D_LL_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_0_preio (
            .PADOEN(N__13245),
            .PADOUT(N__13244),
            .PADIN(N__13243),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9695),
            .DIN0(D_LL_040_in_0),
            .DOUT0(N__4793),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_2_iopad (
            .OE(N__13236),
            .DIN(N__13235),
            .DOUT(N__13234),
            .PACKAGEPIN(D_UM_AMIGA[2]));
    defparam D_UM_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_2_preio (
            .PADOEN(N__13236),
            .PADOUT(N__13235),
            .PADIN(N__13234),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4406),
            .DIN0(D_UM_AMIGA_in_2),
            .DOUT0(N__4685),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_0_iopad (
            .OE(N__13227),
            .DIN(N__13226),
            .DOUT(N__13225),
            .PACKAGEPIN(D_UU_040[0]));
    defparam D_UU_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_0_preio (
            .PADOEN(N__13227),
            .PADOUT(N__13226),
            .PADIN(N__13225),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9461),
            .DIN0(D_UU_040_in_0),
            .DOUT0(N__6839),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_ibuf_iopad (
            .OE(N__13218),
            .DIN(N__13217),
            .DOUT(N__13216),
            .PACKAGEPIN(TCIn));
    defparam TCIn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TCIn_ibuf_preio (
            .PADOEN(N__13218),
            .PADOUT(N__13217),
            .PADIN(N__13216),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TCIn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_040_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_040_ibuf_0_iopad (
            .OE(N__13209),
            .DIN(N__13208),
            .DOUT(N__13207),
            .PACKAGEPIN(A_040[0]));
    defparam A_040_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_040_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_040_ibuf_0_preio (
            .PADOEN(N__13209),
            .PADOUT(N__13208),
            .PADIN(N__13207),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_040_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_0_iopad (
            .OE(N__13200),
            .DIN(N__13199),
            .DOUT(N__13198),
            .PACKAGEPIN(D_LM_AMIGA[0]));
    defparam D_LM_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_0_preio (
            .PADOEN(N__13200),
            .PADOUT(N__13199),
            .PADIN(N__13198),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4268),
            .DIN0(D_LM_AMIGA_in_0),
            .DOUT0(N__5963),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBI_CPUn_obuf_iopad (
            .OE(N__13191),
            .DIN(N__13190),
            .DOUT(N__13189),
            .PACKAGEPIN(TBI_CPUn));
    defparam TBI_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TBI_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TBI_CPUn_obuf_preio (
            .PADOEN(N__13191),
            .PADOUT(N__13190),
            .PADIN(N__13189),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6274),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40A_obuf_iopad (
            .OE(N__13182),
            .DIN(N__13181),
            .DOUT(N__13180),
            .PACKAGEPIN(CLK40A));
    defparam CLK40A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40A_obuf_preio (
            .PADOEN(N__13182),
            .PADOUT(N__13181),
            .PADIN(N__13180),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9596),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_3_iopad (
            .OE(N__13173),
            .DIN(N__13172),
            .DOUT(N__13171),
            .PACKAGEPIN(D_LM_040[3]));
    defparam D_LM_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_3_preio (
            .PADOEN(N__13173),
            .PADOUT(N__13172),
            .PADIN(N__13171),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9743),
            .DIN0(D_LM_040_in_3),
            .DOUT0(N__5147),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_5_iopad (
            .OE(N__13164),
            .DIN(N__13163),
            .DOUT(N__13162),
            .PACKAGEPIN(D_LM_AMIGA[5]));
    defparam D_LM_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_5_preio (
            .PADOEN(N__13164),
            .PADOUT(N__13163),
            .PADIN(N__13162),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4373),
            .DIN0(D_LM_AMIGA_in_5),
            .DOUT0(N__8075),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_6_iopad (
            .OE(N__13155),
            .DIN(N__13154),
            .DOUT(N__13153),
            .PACKAGEPIN(D_LM_040[6]));
    defparam D_LM_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_6_preio (
            .PADOEN(N__13155),
            .PADOUT(N__13154),
            .PADIN(N__13153),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9992),
            .DIN0(D_LM_040_in_6),
            .DOUT0(N__5483),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_5_iopad (
            .OE(N__13146),
            .DIN(N__13145),
            .DOUT(N__13144),
            .PACKAGEPIN(D_UM_040[5]));
    defparam D_UM_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_5_preio (
            .PADOEN(N__13146),
            .PADOUT(N__13145),
            .PADIN(N__13144),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9710),
            .DIN0(D_UM_040_in_5),
            .DOUT0(N__8201),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_3_iopad (
            .OE(N__13137),
            .DIN(N__13136),
            .DOUT(N__13135),
            .PACKAGEPIN(D_LL_AMIGA[3]));
    defparam D_LL_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_3_preio (
            .PADOEN(N__13137),
            .PADOUT(N__13136),
            .PADIN(N__13135),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4154),
            .DIN0(D_LL_AMIGA_in_3),
            .DOUT0(N__6445),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_3_iopad (
            .OE(N__13128),
            .DIN(N__13127),
            .DOUT(N__13126),
            .PACKAGEPIN(D_UU_AMIGA[3]));
    defparam D_UU_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_3_preio (
            .PADOEN(N__13128),
            .PADOUT(N__13127),
            .PADIN(N__13126),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4667),
            .DIN0(D_UU_AMIGA_in_3),
            .DOUT0(N__6323),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_5_iopad (
            .OE(N__13119),
            .DIN(N__13118),
            .DOUT(N__13117),
            .PACKAGEPIN(D_LL_040[5]));
    defparam D_LL_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_5_preio (
            .PADOEN(N__13119),
            .PADOUT(N__13118),
            .PADIN(N__13117),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9875),
            .DIN0(D_LL_040_in_5),
            .DOUT0(N__7439),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_6_iopad (
            .OE(N__13110),
            .DIN(N__13109),
            .DOUT(N__13108),
            .PACKAGEPIN(D_LL_AMIGA[6]));
    defparam D_LL_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_6_preio (
            .PADOEN(N__13110),
            .PADOUT(N__13109),
            .PADIN(N__13108),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4283),
            .DIN0(D_LL_AMIGA_in_6),
            .DOUT0(N__5063),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_6_iopad (
            .OE(N__13101),
            .DIN(N__13100),
            .DOUT(N__13099),
            .PACKAGEPIN(D_UU_AMIGA[6]));
    defparam D_UU_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_6_preio (
            .PADOEN(N__13101),
            .PADOUT(N__13100),
            .PADIN(N__13099),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4823),
            .DIN0(D_UU_AMIGA_in_6),
            .DOUT0(N__5780),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_1_iopad (
            .OE(N__13092),
            .DIN(N__13091),
            .DOUT(N__13090),
            .PACKAGEPIN(D_UM_AMIGA[1]));
    defparam D_UM_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_1_preio (
            .PADOEN(N__13092),
            .PADOUT(N__13091),
            .PADIN(N__13090),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4355),
            .DIN0(D_UM_AMIGA_in_1),
            .DOUT0(N__5519),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_5_iopad (
            .OE(N__13083),
            .DIN(N__13082),
            .DOUT(N__13081),
            .PACKAGEPIN(D_UU_040[5]));
    defparam D_UU_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_5_preio (
            .PADOEN(N__13083),
            .PADOUT(N__13082),
            .PADIN(N__13081),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9545),
            .DIN0(D_UU_040_in_5),
            .DOUT0(N__6989),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAMA_obuf_iopad (
            .OE(N__13074),
            .DIN(N__13073),
            .DOUT(N__13072),
            .PACKAGEPIN(CLKRAMA));
    defparam CLKRAMA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAMA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAMA_obuf_preio (
            .PADOEN(N__13074),
            .PADOUT(N__13073),
            .PADIN(N__13072),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9606),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_2_iopad (
            .OE(N__13065),
            .DIN(N__13064),
            .DOUT(N__13063),
            .PACKAGEPIN(D_LL_040[2]));
    defparam D_LL_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_2_preio (
            .PADOEN(N__13065),
            .PADOUT(N__13064),
            .PADIN(N__13063),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9839),
            .DIN0(D_LL_040_in_2),
            .DOUT0(N__5669),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCI_CPUn_obuf_iopad (
            .OE(N__13056),
            .DIN(N__13055),
            .DOUT(N__13054),
            .PACKAGEPIN(TCI_CPUn));
    defparam TCI_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TCI_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TCI_CPUn_obuf_preio (
            .PADOEN(N__13056),
            .PADOUT(N__13055),
            .PADIN(N__13054),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4064),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_4_iopad (
            .OE(N__13047),
            .DIN(N__13046),
            .DOUT(N__13045),
            .PACKAGEPIN(D_UM_AMIGA[4]));
    defparam D_UM_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_4_preio (
            .PADOEN(N__13047),
            .PADOUT(N__13046),
            .PADIN(N__13045),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4469),
            .DIN0(D_UM_AMIGA_in_4),
            .DOUT0(N__9206),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_6_iopad (
            .OE(N__13038),
            .DIN(N__13037),
            .DOUT(N__13036),
            .PACKAGEPIN(D_LM_AMIGA[6]));
    defparam D_LM_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_6_preio (
            .PADOEN(N__13038),
            .PADOUT(N__13037),
            .PADIN(N__13036),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4325),
            .DIN0(D_LM_AMIGA_in_6),
            .DOUT0(N__5819),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__13029),
            .DIN(N__13028),
            .DOUT(N__13027),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__13029),
            .PADOUT(N__13028),
            .PADIN(N__13027),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_5_iopad (
            .OE(N__13020),
            .DIN(N__13019),
            .DOUT(N__13018),
            .PACKAGEPIN(D_LM_040[5]));
    defparam D_LM_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_5_preio (
            .PADOEN(N__13020),
            .PADOUT(N__13019),
            .PADIN(N__13018),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9890),
            .DIN0(D_LM_040_in_5),
            .DOUT0(N__5984),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_6_iopad (
            .OE(N__13011),
            .DIN(N__13010),
            .DOUT(N__13009),
            .PACKAGEPIN(D_UM_040[6]));
    defparam D_UM_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_6_preio (
            .PADOEN(N__13011),
            .PADOUT(N__13010),
            .PADIN(N__13009),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10016),
            .DIN0(D_UM_040_in_6),
            .DOUT0(N__9287),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_3_iopad (
            .OE(N__13002),
            .DIN(N__13001),
            .DOUT(N__13000),
            .PACKAGEPIN(D_UM_040[3]));
    defparam D_UM_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_3_preio (
            .PADOEN(N__13002),
            .PADOUT(N__13001),
            .PADIN(N__13000),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__12344),
            .DIN0(D_UM_040_in_3),
            .DOUT0(N__7478),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_5_iopad (
            .OE(N__12993),
            .DIN(N__12992),
            .DOUT(N__12991),
            .PACKAGEPIN(D_UU_AMIGA[5]));
    defparam D_UU_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_5_preio (
            .PADOEN(N__12993),
            .PADOUT(N__12992),
            .PADIN(N__12991),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4643),
            .DIN0(D_UU_AMIGA_in_5),
            .DOUT0(N__8027),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_7_iopad (
            .OE(N__12984),
            .DIN(N__12983),
            .DOUT(N__12982),
            .PACKAGEPIN(D_LL_040[7]));
    defparam D_LL_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_7_preio (
            .PADOEN(N__12984),
            .PADOUT(N__12983),
            .PADIN(N__12982),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9773),
            .DIN0(D_LL_040_in_7),
            .DOUT0(N__6791),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_4_iopad (
            .OE(N__12975),
            .DIN(N__12974),
            .DOUT(N__12973),
            .PACKAGEPIN(D_LL_AMIGA[4]));
    defparam D_LL_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_4_preio (
            .PADOEN(N__12975),
            .PADOUT(N__12974),
            .PADIN(N__12973),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4448),
            .DIN0(D_LL_AMIGA_in_4),
            .DOUT0(N__9269),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_3_iopad (
            .OE(N__12966),
            .DIN(N__12965),
            .DOUT(N__12964),
            .PACKAGEPIN(D_UU_040[3]));
    defparam D_UU_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_3_preio (
            .PADOEN(N__12966),
            .PADOUT(N__12965),
            .PADIN(N__12964),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__12323),
            .DIN0(D_UU_040_in_3),
            .DOUT0(N__7949),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TEA_CPUn_obuf_iopad (
            .OE(N__12957),
            .DIN(N__12956),
            .DOUT(N__12955),
            .PACKAGEPIN(TEA_CPUn));
    defparam TEA_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TEA_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TEA_CPUn_obuf_preio (
            .PADOEN(N__12957),
            .PADOUT(N__12956),
            .PADIN(N__12955),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7340),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_3_iopad (
            .OE(N__12948),
            .DIN(N__12947),
            .DOUT(N__12946),
            .PACKAGEPIN(D_LM_AMIGA[3]));
    defparam D_LM_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_3_preio (
            .PADOEN(N__12948),
            .PADOUT(N__12947),
            .PADIN(N__12946),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4550),
            .DIN0(D_LM_AMIGA_in_3),
            .DOUT0(N__6383),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_0_iopad (
            .OE(N__12939),
            .DIN(N__12938),
            .DOUT(N__12937),
            .PACKAGEPIN(D_LM_040[0]));
    defparam D_LM_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_0_preio (
            .PADOEN(N__12939),
            .PADOUT(N__12938),
            .PADIN(N__12937),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9758),
            .DIN0(D_LM_040_in_0),
            .DOUT0(N__5630),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_6_iopad (
            .OE(N__12930),
            .DIN(N__12929),
            .DOUT(N__12928),
            .PACKAGEPIN(D_UM_AMIGA[6]));
    defparam D_UM_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_6_preio (
            .PADOEN(N__12930),
            .PADOUT(N__12929),
            .PADIN(N__12928),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4295),
            .DIN0(D_UM_AMIGA_in_6),
            .DOUT0(N__5024),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_AMIGA_obuf_1_iopad.PULLUP=1'b1;
    IO_PAD A_AMIGA_obuf_1_iopad (
            .OE(N__12921),
            .DIN(N__12920),
            .DOUT(N__12919),
            .PACKAGEPIN(A_AMIGA[1]));
    defparam A_AMIGA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_AMIGA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO A_AMIGA_obuf_1_preio (
            .PADOEN(N__12921),
            .PADOUT(N__12920),
            .PADIN(N__12919),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4598),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_4_iopad (
            .OE(N__12912),
            .DIN(N__12911),
            .DOUT(N__12910),
            .PACKAGEPIN(D_UM_040[4]));
    defparam D_UM_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_4_preio (
            .PADOEN(N__12912),
            .PADOUT(N__12911),
            .PADIN(N__12910),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9725),
            .DIN0(D_UM_040_in_4),
            .DOUT0(N__8414),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_0_iopad (
            .OE(N__12903),
            .DIN(N__12902),
            .DOUT(N__12901),
            .PACKAGEPIN(D_UU_AMIGA[0]));
    defparam D_UU_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_0_preio (
            .PADOEN(N__12903),
            .PADOUT(N__12902),
            .PADIN(N__12901),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4976),
            .DIN0(D_UU_AMIGA_in_0),
            .DOUT0(N__5894),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_4_iopad (
            .OE(N__12894),
            .DIN(N__12893),
            .DOUT(N__12892),
            .PACKAGEPIN(D_LL_040[4]));
    defparam D_LL_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_4_preio (
            .PADOEN(N__12894),
            .PADOUT(N__12893),
            .PADIN(N__12892),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9422),
            .DIN0(D_LL_040_in_4),
            .DOUT0(N__5261),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_7_iopad (
            .OE(N__12885),
            .DIN(N__12884),
            .DOUT(N__12883),
            .PACKAGEPIN(D_LL_AMIGA[7]));
    defparam D_LL_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_7_preio (
            .PADOEN(N__12885),
            .PADOUT(N__12884),
            .PADIN(N__12883),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4256),
            .DIN0(D_LL_AMIGA_in_7),
            .DOUT0(N__8894),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_4_iopad (
            .OE(N__12876),
            .DIN(N__12875),
            .DOUT(N__12874),
            .PACKAGEPIN(D_UU_040[4]));
    defparam D_UU_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_4_preio (
            .PADOEN(N__12876),
            .PADOUT(N__12875),
            .PADIN(N__12874),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9503),
            .DIN0(D_UU_040_in_4),
            .DOUT0(N__7562),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_5_iopad (
            .OE(N__12867),
            .DIN(N__12866),
            .DOUT(N__12865),
            .PACKAGEPIN(D_UM_AMIGA[5]));
    defparam D_UM_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_5_preio (
            .PADOEN(N__12867),
            .PADOUT(N__12866),
            .PADIN(N__12865),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4961),
            .DIN0(D_UM_AMIGA_in_5),
            .DOUT0(N__5324),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__3278 (
            .O(N__12848),
            .I(N__12845));
    LocalMux I__3277 (
            .O(N__12845),
            .I(N__12828));
    ClkMux I__3276 (
            .O(N__12844),
            .I(N__12659));
    ClkMux I__3275 (
            .O(N__12843),
            .I(N__12659));
    ClkMux I__3274 (
            .O(N__12842),
            .I(N__12659));
    ClkMux I__3273 (
            .O(N__12841),
            .I(N__12659));
    ClkMux I__3272 (
            .O(N__12840),
            .I(N__12659));
    ClkMux I__3271 (
            .O(N__12839),
            .I(N__12659));
    ClkMux I__3270 (
            .O(N__12838),
            .I(N__12659));
    ClkMux I__3269 (
            .O(N__12837),
            .I(N__12659));
    ClkMux I__3268 (
            .O(N__12836),
            .I(N__12659));
    ClkMux I__3267 (
            .O(N__12835),
            .I(N__12659));
    ClkMux I__3266 (
            .O(N__12834),
            .I(N__12659));
    ClkMux I__3265 (
            .O(N__12833),
            .I(N__12659));
    ClkMux I__3264 (
            .O(N__12832),
            .I(N__12659));
    ClkMux I__3263 (
            .O(N__12831),
            .I(N__12659));
    Glb2LocalMux I__3262 (
            .O(N__12828),
            .I(N__12659));
    ClkMux I__3261 (
            .O(N__12827),
            .I(N__12659));
    ClkMux I__3260 (
            .O(N__12826),
            .I(N__12659));
    ClkMux I__3259 (
            .O(N__12825),
            .I(N__12659));
    ClkMux I__3258 (
            .O(N__12824),
            .I(N__12659));
    ClkMux I__3257 (
            .O(N__12823),
            .I(N__12659));
    ClkMux I__3256 (
            .O(N__12822),
            .I(N__12659));
    ClkMux I__3255 (
            .O(N__12821),
            .I(N__12659));
    ClkMux I__3254 (
            .O(N__12820),
            .I(N__12659));
    ClkMux I__3253 (
            .O(N__12819),
            .I(N__12659));
    ClkMux I__3252 (
            .O(N__12818),
            .I(N__12659));
    ClkMux I__3251 (
            .O(N__12817),
            .I(N__12659));
    ClkMux I__3250 (
            .O(N__12816),
            .I(N__12659));
    ClkMux I__3249 (
            .O(N__12815),
            .I(N__12659));
    ClkMux I__3248 (
            .O(N__12814),
            .I(N__12659));
    ClkMux I__3247 (
            .O(N__12813),
            .I(N__12659));
    ClkMux I__3246 (
            .O(N__12812),
            .I(N__12659));
    ClkMux I__3245 (
            .O(N__12811),
            .I(N__12659));
    ClkMux I__3244 (
            .O(N__12810),
            .I(N__12659));
    ClkMux I__3243 (
            .O(N__12809),
            .I(N__12659));
    ClkMux I__3242 (
            .O(N__12808),
            .I(N__12659));
    ClkMux I__3241 (
            .O(N__12807),
            .I(N__12659));
    ClkMux I__3240 (
            .O(N__12806),
            .I(N__12659));
    ClkMux I__3239 (
            .O(N__12805),
            .I(N__12659));
    ClkMux I__3238 (
            .O(N__12804),
            .I(N__12659));
    ClkMux I__3237 (
            .O(N__12803),
            .I(N__12659));
    ClkMux I__3236 (
            .O(N__12802),
            .I(N__12659));
    ClkMux I__3235 (
            .O(N__12801),
            .I(N__12659));
    ClkMux I__3234 (
            .O(N__12800),
            .I(N__12659));
    ClkMux I__3233 (
            .O(N__12799),
            .I(N__12659));
    ClkMux I__3232 (
            .O(N__12798),
            .I(N__12659));
    ClkMux I__3231 (
            .O(N__12797),
            .I(N__12659));
    ClkMux I__3230 (
            .O(N__12796),
            .I(N__12659));
    ClkMux I__3229 (
            .O(N__12795),
            .I(N__12659));
    ClkMux I__3228 (
            .O(N__12794),
            .I(N__12659));
    ClkMux I__3227 (
            .O(N__12793),
            .I(N__12659));
    ClkMux I__3226 (
            .O(N__12792),
            .I(N__12659));
    ClkMux I__3225 (
            .O(N__12791),
            .I(N__12659));
    ClkMux I__3224 (
            .O(N__12790),
            .I(N__12659));
    ClkMux I__3223 (
            .O(N__12789),
            .I(N__12659));
    ClkMux I__3222 (
            .O(N__12788),
            .I(N__12659));
    ClkMux I__3221 (
            .O(N__12787),
            .I(N__12659));
    ClkMux I__3220 (
            .O(N__12786),
            .I(N__12659));
    ClkMux I__3219 (
            .O(N__12785),
            .I(N__12659));
    ClkMux I__3218 (
            .O(N__12784),
            .I(N__12659));
    ClkMux I__3217 (
            .O(N__12783),
            .I(N__12659));
    ClkMux I__3216 (
            .O(N__12782),
            .I(N__12659));
    GlobalMux I__3215 (
            .O(N__12659),
            .I(CLK40));
    CEMux I__3214 (
            .O(N__12656),
            .I(N__12521));
    CEMux I__3213 (
            .O(N__12655),
            .I(N__12521));
    CEMux I__3212 (
            .O(N__12654),
            .I(N__12521));
    CEMux I__3211 (
            .O(N__12653),
            .I(N__12521));
    CEMux I__3210 (
            .O(N__12652),
            .I(N__12521));
    CEMux I__3209 (
            .O(N__12651),
            .I(N__12521));
    CEMux I__3208 (
            .O(N__12650),
            .I(N__12521));
    CEMux I__3207 (
            .O(N__12649),
            .I(N__12521));
    CEMux I__3206 (
            .O(N__12648),
            .I(N__12521));
    CEMux I__3205 (
            .O(N__12647),
            .I(N__12521));
    CEMux I__3204 (
            .O(N__12646),
            .I(N__12521));
    CEMux I__3203 (
            .O(N__12645),
            .I(N__12521));
    CEMux I__3202 (
            .O(N__12644),
            .I(N__12521));
    CEMux I__3201 (
            .O(N__12643),
            .I(N__12521));
    CEMux I__3200 (
            .O(N__12642),
            .I(N__12521));
    CEMux I__3199 (
            .O(N__12641),
            .I(N__12521));
    CEMux I__3198 (
            .O(N__12640),
            .I(N__12521));
    CEMux I__3197 (
            .O(N__12639),
            .I(N__12521));
    CEMux I__3196 (
            .O(N__12638),
            .I(N__12521));
    CEMux I__3195 (
            .O(N__12637),
            .I(N__12521));
    CEMux I__3194 (
            .O(N__12636),
            .I(N__12521));
    CEMux I__3193 (
            .O(N__12635),
            .I(N__12521));
    CEMux I__3192 (
            .O(N__12634),
            .I(N__12521));
    CEMux I__3191 (
            .O(N__12633),
            .I(N__12521));
    CEMux I__3190 (
            .O(N__12632),
            .I(N__12521));
    CEMux I__3189 (
            .O(N__12631),
            .I(N__12521));
    CEMux I__3188 (
            .O(N__12630),
            .I(N__12521));
    CEMux I__3187 (
            .O(N__12629),
            .I(N__12521));
    CEMux I__3186 (
            .O(N__12628),
            .I(N__12521));
    CEMux I__3185 (
            .O(N__12627),
            .I(N__12521));
    CEMux I__3184 (
            .O(N__12626),
            .I(N__12521));
    CEMux I__3183 (
            .O(N__12625),
            .I(N__12521));
    CEMux I__3182 (
            .O(N__12624),
            .I(N__12521));
    CEMux I__3181 (
            .O(N__12623),
            .I(N__12521));
    CEMux I__3180 (
            .O(N__12622),
            .I(N__12521));
    CEMux I__3179 (
            .O(N__12621),
            .I(N__12521));
    CEMux I__3178 (
            .O(N__12620),
            .I(N__12521));
    CEMux I__3177 (
            .O(N__12619),
            .I(N__12521));
    CEMux I__3176 (
            .O(N__12618),
            .I(N__12521));
    CEMux I__3175 (
            .O(N__12617),
            .I(N__12521));
    CEMux I__3174 (
            .O(N__12616),
            .I(N__12521));
    CEMux I__3173 (
            .O(N__12615),
            .I(N__12521));
    CEMux I__3172 (
            .O(N__12614),
            .I(N__12521));
    CEMux I__3171 (
            .O(N__12613),
            .I(N__12521));
    CEMux I__3170 (
            .O(N__12612),
            .I(N__12521));
    GlobalMux I__3169 (
            .O(N__12521),
            .I(N__12518));
    gio2CtrlBuf I__3168 (
            .O(N__12518),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_g_0 ));
    InMux I__3167 (
            .O(N__12515),
            .I(N__12512));
    LocalMux I__3166 (
            .O(N__12512),
            .I(N__12459));
    SRMux I__3165 (
            .O(N__12511),
            .I(N__12356));
    SRMux I__3164 (
            .O(N__12510),
            .I(N__12356));
    SRMux I__3163 (
            .O(N__12509),
            .I(N__12356));
    SRMux I__3162 (
            .O(N__12508),
            .I(N__12356));
    SRMux I__3161 (
            .O(N__12507),
            .I(N__12356));
    SRMux I__3160 (
            .O(N__12506),
            .I(N__12356));
    SRMux I__3159 (
            .O(N__12505),
            .I(N__12356));
    SRMux I__3158 (
            .O(N__12504),
            .I(N__12356));
    SRMux I__3157 (
            .O(N__12503),
            .I(N__12356));
    SRMux I__3156 (
            .O(N__12502),
            .I(N__12356));
    SRMux I__3155 (
            .O(N__12501),
            .I(N__12356));
    SRMux I__3154 (
            .O(N__12500),
            .I(N__12356));
    SRMux I__3153 (
            .O(N__12499),
            .I(N__12356));
    SRMux I__3152 (
            .O(N__12498),
            .I(N__12356));
    SRMux I__3151 (
            .O(N__12497),
            .I(N__12356));
    SRMux I__3150 (
            .O(N__12496),
            .I(N__12356));
    SRMux I__3149 (
            .O(N__12495),
            .I(N__12356));
    SRMux I__3148 (
            .O(N__12494),
            .I(N__12356));
    SRMux I__3147 (
            .O(N__12493),
            .I(N__12356));
    SRMux I__3146 (
            .O(N__12492),
            .I(N__12356));
    SRMux I__3145 (
            .O(N__12491),
            .I(N__12356));
    SRMux I__3144 (
            .O(N__12490),
            .I(N__12356));
    SRMux I__3143 (
            .O(N__12489),
            .I(N__12356));
    SRMux I__3142 (
            .O(N__12488),
            .I(N__12356));
    SRMux I__3141 (
            .O(N__12487),
            .I(N__12356));
    SRMux I__3140 (
            .O(N__12486),
            .I(N__12356));
    SRMux I__3139 (
            .O(N__12485),
            .I(N__12356));
    SRMux I__3138 (
            .O(N__12484),
            .I(N__12356));
    SRMux I__3137 (
            .O(N__12483),
            .I(N__12356));
    SRMux I__3136 (
            .O(N__12482),
            .I(N__12356));
    SRMux I__3135 (
            .O(N__12481),
            .I(N__12356));
    SRMux I__3134 (
            .O(N__12480),
            .I(N__12356));
    SRMux I__3133 (
            .O(N__12479),
            .I(N__12356));
    SRMux I__3132 (
            .O(N__12478),
            .I(N__12356));
    SRMux I__3131 (
            .O(N__12477),
            .I(N__12356));
    SRMux I__3130 (
            .O(N__12476),
            .I(N__12356));
    SRMux I__3129 (
            .O(N__12475),
            .I(N__12356));
    SRMux I__3128 (
            .O(N__12474),
            .I(N__12356));
    SRMux I__3127 (
            .O(N__12473),
            .I(N__12356));
    SRMux I__3126 (
            .O(N__12472),
            .I(N__12356));
    SRMux I__3125 (
            .O(N__12471),
            .I(N__12356));
    SRMux I__3124 (
            .O(N__12470),
            .I(N__12356));
    SRMux I__3123 (
            .O(N__12469),
            .I(N__12356));
    SRMux I__3122 (
            .O(N__12468),
            .I(N__12356));
    SRMux I__3121 (
            .O(N__12467),
            .I(N__12356));
    SRMux I__3120 (
            .O(N__12466),
            .I(N__12356));
    SRMux I__3119 (
            .O(N__12465),
            .I(N__12356));
    SRMux I__3118 (
            .O(N__12464),
            .I(N__12356));
    SRMux I__3117 (
            .O(N__12463),
            .I(N__12356));
    SRMux I__3116 (
            .O(N__12462),
            .I(N__12356));
    Glb2LocalMux I__3115 (
            .O(N__12459),
            .I(N__12356));
    GlobalMux I__3114 (
            .O(N__12356),
            .I(N__12353));
    gio2CtrlBuf I__3113 (
            .O(N__12353),
            .I(RESETn_c_i_g));
    InMux I__3112 (
            .O(N__12350),
            .I(N__12347));
    LocalMux I__3111 (
            .O(N__12347),
            .I(READ_CYCLE_ACTIVE_rep11_i_ess));
    IoInMux I__3110 (
            .O(N__12344),
            .I(N__12341));
    LocalMux I__3109 (
            .O(N__12341),
            .I(N__12338));
    Span4Mux_s3_h I__3108 (
            .O(N__12338),
            .I(N__12335));
    Span4Mux_v I__3107 (
            .O(N__12335),
            .I(N__12332));
    Odrv4 I__3106 (
            .O(N__12332),
            .I(N_192_i));
    InMux I__3105 (
            .O(N__12329),
            .I(N__12326));
    LocalMux I__3104 (
            .O(N__12326),
            .I(READ_CYCLE_ACTIVE_rep3_i_ess));
    IoInMux I__3103 (
            .O(N__12323),
            .I(N__12320));
    LocalMux I__3102 (
            .O(N__12320),
            .I(N__12317));
    IoSpan4Mux I__3101 (
            .O(N__12317),
            .I(N__12314));
    Span4Mux_s3_v I__3100 (
            .O(N__12314),
            .I(N__12311));
    Span4Mux_v I__3099 (
            .O(N__12311),
            .I(N__12308));
    Odrv4 I__3098 (
            .O(N__12308),
            .I(N_184_i));
    InMux I__3097 (
            .O(N__12305),
            .I(N__12302));
    LocalMux I__3096 (
            .O(N__12302),
            .I(READ_CYCLE_ACTIVE_rep15_i_ess));
    IoInMux I__3095 (
            .O(N__12299),
            .I(N__12296));
    LocalMux I__3094 (
            .O(N__12296),
            .I(N__12293));
    IoSpan4Mux I__3093 (
            .O(N__12293),
            .I(N__12290));
    Span4Mux_s3_h I__3092 (
            .O(N__12290),
            .I(N__12287));
    Odrv4 I__3091 (
            .O(N__12287),
            .I(N_196_i));
    InMux I__3090 (
            .O(N__12284),
            .I(N__12281));
    LocalMux I__3089 (
            .O(N__12281),
            .I(READ_CYCLE_ACTIVE_rep1_i_ess));
    IoInMux I__3088 (
            .O(N__12278),
            .I(N__12275));
    LocalMux I__3087 (
            .O(N__12275),
            .I(N__12272));
    Span12Mux_s4_h I__3086 (
            .O(N__12272),
            .I(N__12269));
    Odrv12 I__3085 (
            .O(N__12269),
            .I(N_182_i));
    InMux I__3084 (
            .O(N__12266),
            .I(N__12263));
    LocalMux I__3083 (
            .O(N__12263),
            .I(READ_CYCLE_ACTIVE_rep13_i_ess));
    CascadeMux I__3082 (
            .O(N__12260),
            .I(N__12253));
    InMux I__3081 (
            .O(N__12259),
            .I(N__12248));
    InMux I__3080 (
            .O(N__12258),
            .I(N__12245));
    InMux I__3079 (
            .O(N__12257),
            .I(N__12239));
    InMux I__3078 (
            .O(N__12256),
            .I(N__12236));
    InMux I__3077 (
            .O(N__12253),
            .I(N__12231));
    InMux I__3076 (
            .O(N__12252),
            .I(N__12231));
    InMux I__3075 (
            .O(N__12251),
            .I(N__12223));
    LocalMux I__3074 (
            .O(N__12248),
            .I(N__12218));
    LocalMux I__3073 (
            .O(N__12245),
            .I(N__12218));
    InMux I__3072 (
            .O(N__12244),
            .I(N__12213));
    InMux I__3071 (
            .O(N__12243),
            .I(N__12210));
    InMux I__3070 (
            .O(N__12242),
            .I(N__12207));
    LocalMux I__3069 (
            .O(N__12239),
            .I(N__12197));
    LocalMux I__3068 (
            .O(N__12236),
            .I(N__12197));
    LocalMux I__3067 (
            .O(N__12231),
            .I(N__12194));
    InMux I__3066 (
            .O(N__12230),
            .I(N__12189));
    InMux I__3065 (
            .O(N__12229),
            .I(N__12189));
    InMux I__3064 (
            .O(N__12228),
            .I(N__12186));
    InMux I__3063 (
            .O(N__12227),
            .I(N__12183));
    InMux I__3062 (
            .O(N__12226),
            .I(N__12180));
    LocalMux I__3061 (
            .O(N__12223),
            .I(N__12175));
    Span4Mux_v I__3060 (
            .O(N__12218),
            .I(N__12175));
    InMux I__3059 (
            .O(N__12217),
            .I(N__12172));
    CascadeMux I__3058 (
            .O(N__12216),
            .I(N__12168));
    LocalMux I__3057 (
            .O(N__12213),
            .I(N__12159));
    LocalMux I__3056 (
            .O(N__12210),
            .I(N__12159));
    LocalMux I__3055 (
            .O(N__12207),
            .I(N__12159));
    InMux I__3054 (
            .O(N__12206),
            .I(N__12156));
    InMux I__3053 (
            .O(N__12205),
            .I(N__12153));
    InMux I__3052 (
            .O(N__12204),
            .I(N__12150));
    InMux I__3051 (
            .O(N__12203),
            .I(N__12147));
    InMux I__3050 (
            .O(N__12202),
            .I(N__12144));
    Span4Mux_v I__3049 (
            .O(N__12197),
            .I(N__12127));
    Span4Mux_h I__3048 (
            .O(N__12194),
            .I(N__12127));
    LocalMux I__3047 (
            .O(N__12189),
            .I(N__12127));
    LocalMux I__3046 (
            .O(N__12186),
            .I(N__12127));
    LocalMux I__3045 (
            .O(N__12183),
            .I(N__12127));
    LocalMux I__3044 (
            .O(N__12180),
            .I(N__12127));
    Span4Mux_h I__3043 (
            .O(N__12175),
            .I(N__12127));
    LocalMux I__3042 (
            .O(N__12172),
            .I(N__12127));
    InMux I__3041 (
            .O(N__12171),
            .I(N__12124));
    InMux I__3040 (
            .O(N__12168),
            .I(N__12121));
    InMux I__3039 (
            .O(N__12167),
            .I(N__12118));
    InMux I__3038 (
            .O(N__12166),
            .I(N__12113));
    Span4Mux_v I__3037 (
            .O(N__12159),
            .I(N__12106));
    LocalMux I__3036 (
            .O(N__12156),
            .I(N__12106));
    LocalMux I__3035 (
            .O(N__12153),
            .I(N__12106));
    LocalMux I__3034 (
            .O(N__12150),
            .I(N__12095));
    LocalMux I__3033 (
            .O(N__12147),
            .I(N__12095));
    LocalMux I__3032 (
            .O(N__12144),
            .I(N__12095));
    Span4Mux_v I__3031 (
            .O(N__12127),
            .I(N__12095));
    LocalMux I__3030 (
            .O(N__12124),
            .I(N__12095));
    LocalMux I__3029 (
            .O(N__12121),
            .I(N__12084));
    LocalMux I__3028 (
            .O(N__12118),
            .I(N__12084));
    InMux I__3027 (
            .O(N__12117),
            .I(N__12081));
    InMux I__3026 (
            .O(N__12116),
            .I(N__12078));
    LocalMux I__3025 (
            .O(N__12113),
            .I(N__12075));
    Span4Mux_v I__3024 (
            .O(N__12106),
            .I(N__12068));
    Span4Mux_v I__3023 (
            .O(N__12095),
            .I(N__12068));
    InMux I__3022 (
            .O(N__12094),
            .I(N__12065));
    InMux I__3021 (
            .O(N__12093),
            .I(N__12062));
    InMux I__3020 (
            .O(N__12092),
            .I(N__12059));
    InMux I__3019 (
            .O(N__12091),
            .I(N__12056));
    InMux I__3018 (
            .O(N__12090),
            .I(N__12053));
    InMux I__3017 (
            .O(N__12089),
            .I(N__12039));
    Span4Mux_v I__3016 (
            .O(N__12084),
            .I(N__12032));
    LocalMux I__3015 (
            .O(N__12081),
            .I(N__12032));
    LocalMux I__3014 (
            .O(N__12078),
            .I(N__12032));
    Span4Mux_v I__3013 (
            .O(N__12075),
            .I(N__12029));
    InMux I__3012 (
            .O(N__12074),
            .I(N__12024));
    InMux I__3011 (
            .O(N__12073),
            .I(N__12024));
    Span4Mux_h I__3010 (
            .O(N__12068),
            .I(N__12017));
    LocalMux I__3009 (
            .O(N__12065),
            .I(N__12017));
    LocalMux I__3008 (
            .O(N__12062),
            .I(N__12014));
    LocalMux I__3007 (
            .O(N__12059),
            .I(N__12008));
    LocalMux I__3006 (
            .O(N__12056),
            .I(N__12008));
    LocalMux I__3005 (
            .O(N__12053),
            .I(N__12005));
    InMux I__3004 (
            .O(N__12052),
            .I(N__11998));
    InMux I__3003 (
            .O(N__12051),
            .I(N__11998));
    InMux I__3002 (
            .O(N__12050),
            .I(N__11998));
    InMux I__3001 (
            .O(N__12049),
            .I(N__11995));
    InMux I__3000 (
            .O(N__12048),
            .I(N__11986));
    InMux I__2999 (
            .O(N__12047),
            .I(N__11986));
    InMux I__2998 (
            .O(N__12046),
            .I(N__11986));
    InMux I__2997 (
            .O(N__12045),
            .I(N__11981));
    InMux I__2996 (
            .O(N__12044),
            .I(N__11981));
    InMux I__2995 (
            .O(N__12043),
            .I(N__11976));
    InMux I__2994 (
            .O(N__12042),
            .I(N__11976));
    LocalMux I__2993 (
            .O(N__12039),
            .I(N__11966));
    Sp12to4 I__2992 (
            .O(N__12032),
            .I(N__11966));
    Span4Mux_h I__2991 (
            .O(N__12029),
            .I(N__11961));
    LocalMux I__2990 (
            .O(N__12024),
            .I(N__11961));
    InMux I__2989 (
            .O(N__12023),
            .I(N__11956));
    InMux I__2988 (
            .O(N__12022),
            .I(N__11956));
    Span4Mux_h I__2987 (
            .O(N__12017),
            .I(N__11951));
    Span4Mux_v I__2986 (
            .O(N__12014),
            .I(N__11951));
    InMux I__2985 (
            .O(N__12013),
            .I(N__11948));
    Span4Mux_v I__2984 (
            .O(N__12008),
            .I(N__11945));
    Span4Mux_v I__2983 (
            .O(N__12005),
            .I(N__11942));
    LocalMux I__2982 (
            .O(N__11998),
            .I(N__11939));
    LocalMux I__2981 (
            .O(N__11995),
            .I(N__11934));
    InMux I__2980 (
            .O(N__11994),
            .I(N__11929));
    InMux I__2979 (
            .O(N__11993),
            .I(N__11929));
    LocalMux I__2978 (
            .O(N__11986),
            .I(N__11920));
    LocalMux I__2977 (
            .O(N__11981),
            .I(N__11920));
    LocalMux I__2976 (
            .O(N__11976),
            .I(N__11917));
    InMux I__2975 (
            .O(N__11975),
            .I(N__11908));
    InMux I__2974 (
            .O(N__11974),
            .I(N__11908));
    InMux I__2973 (
            .O(N__11973),
            .I(N__11908));
    InMux I__2972 (
            .O(N__11972),
            .I(N__11908));
    InMux I__2971 (
            .O(N__11971),
            .I(N__11905));
    Span12Mux_v I__2970 (
            .O(N__11966),
            .I(N__11897));
    Sp12to4 I__2969 (
            .O(N__11961),
            .I(N__11894));
    LocalMux I__2968 (
            .O(N__11956),
            .I(N__11891));
    Span4Mux_v I__2967 (
            .O(N__11951),
            .I(N__11888));
    LocalMux I__2966 (
            .O(N__11948),
            .I(N__11885));
    Span4Mux_v I__2965 (
            .O(N__11945),
            .I(N__11882));
    Span4Mux_h I__2964 (
            .O(N__11942),
            .I(N__11877));
    Span4Mux_v I__2963 (
            .O(N__11939),
            .I(N__11877));
    InMux I__2962 (
            .O(N__11938),
            .I(N__11874));
    InMux I__2961 (
            .O(N__11937),
            .I(N__11871));
    Span4Mux_v I__2960 (
            .O(N__11934),
            .I(N__11868));
    LocalMux I__2959 (
            .O(N__11929),
            .I(N__11865));
    InMux I__2958 (
            .O(N__11928),
            .I(N__11858));
    InMux I__2957 (
            .O(N__11927),
            .I(N__11858));
    InMux I__2956 (
            .O(N__11926),
            .I(N__11858));
    InMux I__2955 (
            .O(N__11925),
            .I(N__11855));
    Span4Mux_v I__2954 (
            .O(N__11920),
            .I(N__11848));
    Span4Mux_h I__2953 (
            .O(N__11917),
            .I(N__11848));
    LocalMux I__2952 (
            .O(N__11908),
            .I(N__11848));
    LocalMux I__2951 (
            .O(N__11905),
            .I(N__11845));
    InMux I__2950 (
            .O(N__11904),
            .I(N__11840));
    InMux I__2949 (
            .O(N__11903),
            .I(N__11840));
    InMux I__2948 (
            .O(N__11902),
            .I(N__11833));
    InMux I__2947 (
            .O(N__11901),
            .I(N__11833));
    InMux I__2946 (
            .O(N__11900),
            .I(N__11833));
    Span12Mux_h I__2945 (
            .O(N__11897),
            .I(N__11830));
    Span12Mux_v I__2944 (
            .O(N__11894),
            .I(N__11825));
    Span12Mux_s9_h I__2943 (
            .O(N__11891),
            .I(N__11825));
    Sp12to4 I__2942 (
            .O(N__11888),
            .I(N__11820));
    Span12Mux_v I__2941 (
            .O(N__11885),
            .I(N__11820));
    Span4Mux_v I__2940 (
            .O(N__11882),
            .I(N__11815));
    Span4Mux_v I__2939 (
            .O(N__11877),
            .I(N__11815));
    LocalMux I__2938 (
            .O(N__11874),
            .I(N__11810));
    LocalMux I__2937 (
            .O(N__11871),
            .I(N__11810));
    Span4Mux_h I__2936 (
            .O(N__11868),
            .I(N__11801));
    Span4Mux_v I__2935 (
            .O(N__11865),
            .I(N__11801));
    LocalMux I__2934 (
            .O(N__11858),
            .I(N__11801));
    LocalMux I__2933 (
            .O(N__11855),
            .I(N__11801));
    Span4Mux_v I__2932 (
            .O(N__11848),
            .I(N__11792));
    Span4Mux_h I__2931 (
            .O(N__11845),
            .I(N__11792));
    LocalMux I__2930 (
            .O(N__11840),
            .I(N__11792));
    LocalMux I__2929 (
            .O(N__11833),
            .I(N__11792));
    Span12Mux_h I__2928 (
            .O(N__11830),
            .I(N__11789));
    Span12Mux_h I__2927 (
            .O(N__11825),
            .I(N__11786));
    Span12Mux_h I__2926 (
            .O(N__11820),
            .I(N__11779));
    Sp12to4 I__2925 (
            .O(N__11815),
            .I(N__11779));
    Span12Mux_v I__2924 (
            .O(N__11810),
            .I(N__11779));
    Span4Mux_v I__2923 (
            .O(N__11801),
            .I(N__11774));
    Span4Mux_v I__2922 (
            .O(N__11792),
            .I(N__11774));
    Odrv12 I__2921 (
            .O(N__11789),
            .I(BGn_c));
    Odrv12 I__2920 (
            .O(N__11786),
            .I(BGn_c));
    Odrv12 I__2919 (
            .O(N__11779),
            .I(BGn_c));
    Odrv4 I__2918 (
            .O(N__11774),
            .I(BGn_c));
    CascadeMux I__2917 (
            .O(N__11765),
            .I(N__11761));
    InMux I__2916 (
            .O(N__11764),
            .I(N__11755));
    InMux I__2915 (
            .O(N__11761),
            .I(N__11752));
    CascadeMux I__2914 (
            .O(N__11760),
            .I(N__11749));
    CascadeMux I__2913 (
            .O(N__11759),
            .I(N__11745));
    CascadeMux I__2912 (
            .O(N__11758),
            .I(N__11741));
    LocalMux I__2911 (
            .O(N__11755),
            .I(N__11734));
    LocalMux I__2910 (
            .O(N__11752),
            .I(N__11734));
    InMux I__2909 (
            .O(N__11749),
            .I(N__11731));
    InMux I__2908 (
            .O(N__11748),
            .I(N__11726));
    InMux I__2907 (
            .O(N__11745),
            .I(N__11726));
    InMux I__2906 (
            .O(N__11744),
            .I(N__11723));
    InMux I__2905 (
            .O(N__11741),
            .I(N__11720));
    CascadeMux I__2904 (
            .O(N__11740),
            .I(N__11717));
    CascadeMux I__2903 (
            .O(N__11739),
            .I(N__11712));
    Span4Mux_v I__2902 (
            .O(N__11734),
            .I(N__11692));
    LocalMux I__2901 (
            .O(N__11731),
            .I(N__11692));
    LocalMux I__2900 (
            .O(N__11726),
            .I(N__11692));
    LocalMux I__2899 (
            .O(N__11723),
            .I(N__11692));
    LocalMux I__2898 (
            .O(N__11720),
            .I(N__11692));
    InMux I__2897 (
            .O(N__11717),
            .I(N__11689));
    CascadeMux I__2896 (
            .O(N__11716),
            .I(N__11685));
    InMux I__2895 (
            .O(N__11715),
            .I(N__11677));
    InMux I__2894 (
            .O(N__11712),
            .I(N__11677));
    InMux I__2893 (
            .O(N__11711),
            .I(N__11677));
    InMux I__2892 (
            .O(N__11710),
            .I(N__11674));
    InMux I__2891 (
            .O(N__11709),
            .I(N__11671));
    CascadeMux I__2890 (
            .O(N__11708),
            .I(N__11668));
    CascadeMux I__2889 (
            .O(N__11707),
            .I(N__11663));
    CascadeMux I__2888 (
            .O(N__11706),
            .I(N__11659));
    CascadeMux I__2887 (
            .O(N__11705),
            .I(N__11656));
    InMux I__2886 (
            .O(N__11704),
            .I(N__11651));
    CascadeMux I__2885 (
            .O(N__11703),
            .I(N__11646));
    Span4Mux_v I__2884 (
            .O(N__11692),
            .I(N__11641));
    LocalMux I__2883 (
            .O(N__11689),
            .I(N__11641));
    InMux I__2882 (
            .O(N__11688),
            .I(N__11636));
    InMux I__2881 (
            .O(N__11685),
            .I(N__11636));
    InMux I__2880 (
            .O(N__11684),
            .I(N__11633));
    LocalMux I__2879 (
            .O(N__11677),
            .I(N__11623));
    LocalMux I__2878 (
            .O(N__11674),
            .I(N__11623));
    LocalMux I__2877 (
            .O(N__11671),
            .I(N__11623));
    InMux I__2876 (
            .O(N__11668),
            .I(N__11618));
    InMux I__2875 (
            .O(N__11667),
            .I(N__11618));
    InMux I__2874 (
            .O(N__11666),
            .I(N__11609));
    InMux I__2873 (
            .O(N__11663),
            .I(N__11609));
    InMux I__2872 (
            .O(N__11662),
            .I(N__11609));
    InMux I__2871 (
            .O(N__11659),
            .I(N__11609));
    InMux I__2870 (
            .O(N__11656),
            .I(N__11602));
    CascadeMux I__2869 (
            .O(N__11655),
            .I(N__11598));
    CascadeMux I__2868 (
            .O(N__11654),
            .I(N__11590));
    LocalMux I__2867 (
            .O(N__11651),
            .I(N__11581));
    InMux I__2866 (
            .O(N__11650),
            .I(N__11576));
    InMux I__2865 (
            .O(N__11649),
            .I(N__11576));
    InMux I__2864 (
            .O(N__11646),
            .I(N__11573));
    Span4Mux_v I__2863 (
            .O(N__11641),
            .I(N__11566));
    LocalMux I__2862 (
            .O(N__11636),
            .I(N__11566));
    LocalMux I__2861 (
            .O(N__11633),
            .I(N__11566));
    InMux I__2860 (
            .O(N__11632),
            .I(N__11561));
    InMux I__2859 (
            .O(N__11631),
            .I(N__11561));
    CascadeMux I__2858 (
            .O(N__11630),
            .I(N__11555));
    Span4Mux_v I__2857 (
            .O(N__11623),
            .I(N__11547));
    LocalMux I__2856 (
            .O(N__11618),
            .I(N__11547));
    LocalMux I__2855 (
            .O(N__11609),
            .I(N__11547));
    InMux I__2854 (
            .O(N__11608),
            .I(N__11544));
    InMux I__2853 (
            .O(N__11607),
            .I(N__11539));
    InMux I__2852 (
            .O(N__11606),
            .I(N__11539));
    InMux I__2851 (
            .O(N__11605),
            .I(N__11532));
    LocalMux I__2850 (
            .O(N__11602),
            .I(N__11529));
    InMux I__2849 (
            .O(N__11601),
            .I(N__11526));
    InMux I__2848 (
            .O(N__11598),
            .I(N__11523));
    InMux I__2847 (
            .O(N__11597),
            .I(N__11515));
    InMux I__2846 (
            .O(N__11596),
            .I(N__11515));
    InMux I__2845 (
            .O(N__11595),
            .I(N__11515));
    InMux I__2844 (
            .O(N__11594),
            .I(N__11508));
    InMux I__2843 (
            .O(N__11593),
            .I(N__11508));
    InMux I__2842 (
            .O(N__11590),
            .I(N__11502));
    InMux I__2841 (
            .O(N__11589),
            .I(N__11499));
    InMux I__2840 (
            .O(N__11588),
            .I(N__11496));
    CascadeMux I__2839 (
            .O(N__11587),
            .I(N__11493));
    CascadeMux I__2838 (
            .O(N__11586),
            .I(N__11490));
    CascadeMux I__2837 (
            .O(N__11585),
            .I(N__11485));
    CascadeMux I__2836 (
            .O(N__11584),
            .I(N__11482));
    Span4Mux_v I__2835 (
            .O(N__11581),
            .I(N__11479));
    LocalMux I__2834 (
            .O(N__11576),
            .I(N__11474));
    LocalMux I__2833 (
            .O(N__11573),
            .I(N__11474));
    Span4Mux_v I__2832 (
            .O(N__11566),
            .I(N__11469));
    LocalMux I__2831 (
            .O(N__11561),
            .I(N__11469));
    InMux I__2830 (
            .O(N__11560),
            .I(N__11466));
    InMux I__2829 (
            .O(N__11559),
            .I(N__11461));
    InMux I__2828 (
            .O(N__11558),
            .I(N__11461));
    InMux I__2827 (
            .O(N__11555),
            .I(N__11458));
    CascadeMux I__2826 (
            .O(N__11554),
            .I(N__11454));
    Span4Mux_v I__2825 (
            .O(N__11547),
            .I(N__11448));
    LocalMux I__2824 (
            .O(N__11544),
            .I(N__11448));
    LocalMux I__2823 (
            .O(N__11539),
            .I(N__11445));
    InMux I__2822 (
            .O(N__11538),
            .I(N__11442));
    InMux I__2821 (
            .O(N__11537),
            .I(N__11435));
    InMux I__2820 (
            .O(N__11536),
            .I(N__11435));
    InMux I__2819 (
            .O(N__11535),
            .I(N__11435));
    LocalMux I__2818 (
            .O(N__11532),
            .I(N__11432));
    Span4Mux_h I__2817 (
            .O(N__11529),
            .I(N__11425));
    LocalMux I__2816 (
            .O(N__11526),
            .I(N__11425));
    LocalMux I__2815 (
            .O(N__11523),
            .I(N__11425));
    InMux I__2814 (
            .O(N__11522),
            .I(N__11422));
    LocalMux I__2813 (
            .O(N__11515),
            .I(N__11419));
    InMux I__2812 (
            .O(N__11514),
            .I(N__11416));
    InMux I__2811 (
            .O(N__11513),
            .I(N__11413));
    LocalMux I__2810 (
            .O(N__11508),
            .I(N__11410));
    InMux I__2809 (
            .O(N__11507),
            .I(N__11407));
    InMux I__2808 (
            .O(N__11506),
            .I(N__11404));
    InMux I__2807 (
            .O(N__11505),
            .I(N__11401));
    LocalMux I__2806 (
            .O(N__11502),
            .I(N__11396));
    LocalMux I__2805 (
            .O(N__11499),
            .I(N__11396));
    LocalMux I__2804 (
            .O(N__11496),
            .I(N__11393));
    InMux I__2803 (
            .O(N__11493),
            .I(N__11390));
    InMux I__2802 (
            .O(N__11490),
            .I(N__11383));
    InMux I__2801 (
            .O(N__11489),
            .I(N__11383));
    InMux I__2800 (
            .O(N__11488),
            .I(N__11383));
    InMux I__2799 (
            .O(N__11485),
            .I(N__11380));
    InMux I__2798 (
            .O(N__11482),
            .I(N__11377));
    Span4Mux_v I__2797 (
            .O(N__11479),
            .I(N__11374));
    Span4Mux_v I__2796 (
            .O(N__11474),
            .I(N__11371));
    Span4Mux_h I__2795 (
            .O(N__11469),
            .I(N__11364));
    LocalMux I__2794 (
            .O(N__11466),
            .I(N__11364));
    LocalMux I__2793 (
            .O(N__11461),
            .I(N__11364));
    LocalMux I__2792 (
            .O(N__11458),
            .I(N__11361));
    InMux I__2791 (
            .O(N__11457),
            .I(N__11356));
    InMux I__2790 (
            .O(N__11454),
            .I(N__11356));
    CascadeMux I__2789 (
            .O(N__11453),
            .I(N__11353));
    Span4Mux_v I__2788 (
            .O(N__11448),
            .I(N__11346));
    Span4Mux_v I__2787 (
            .O(N__11445),
            .I(N__11346));
    LocalMux I__2786 (
            .O(N__11442),
            .I(N__11346));
    LocalMux I__2785 (
            .O(N__11435),
            .I(N__11343));
    Span4Mux_v I__2784 (
            .O(N__11432),
            .I(N__11339));
    Span4Mux_h I__2783 (
            .O(N__11425),
            .I(N__11334));
    LocalMux I__2782 (
            .O(N__11422),
            .I(N__11334));
    Span4Mux_h I__2781 (
            .O(N__11419),
            .I(N__11327));
    LocalMux I__2780 (
            .O(N__11416),
            .I(N__11327));
    LocalMux I__2779 (
            .O(N__11413),
            .I(N__11327));
    Span4Mux_h I__2778 (
            .O(N__11410),
            .I(N__11324));
    LocalMux I__2777 (
            .O(N__11407),
            .I(N__11321));
    LocalMux I__2776 (
            .O(N__11404),
            .I(N__11316));
    LocalMux I__2775 (
            .O(N__11401),
            .I(N__11316));
    Span12Mux_v I__2774 (
            .O(N__11396),
            .I(N__11309));
    Span12Mux_s6_h I__2773 (
            .O(N__11393),
            .I(N__11309));
    LocalMux I__2772 (
            .O(N__11390),
            .I(N__11309));
    LocalMux I__2771 (
            .O(N__11383),
            .I(N__11306));
    LocalMux I__2770 (
            .O(N__11380),
            .I(N__11303));
    LocalMux I__2769 (
            .O(N__11377),
            .I(N__11300));
    Span4Mux_v I__2768 (
            .O(N__11374),
            .I(N__11293));
    Span4Mux_h I__2767 (
            .O(N__11371),
            .I(N__11293));
    Span4Mux_v I__2766 (
            .O(N__11364),
            .I(N__11293));
    Span12Mux_s6_h I__2765 (
            .O(N__11361),
            .I(N__11290));
    LocalMux I__2764 (
            .O(N__11356),
            .I(N__11287));
    InMux I__2763 (
            .O(N__11353),
            .I(N__11284));
    Span4Mux_v I__2762 (
            .O(N__11346),
            .I(N__11279));
    Span4Mux_v I__2761 (
            .O(N__11343),
            .I(N__11279));
    InMux I__2760 (
            .O(N__11342),
            .I(N__11276));
    Span4Mux_v I__2759 (
            .O(N__11339),
            .I(N__11271));
    Span4Mux_h I__2758 (
            .O(N__11334),
            .I(N__11271));
    Span4Mux_h I__2757 (
            .O(N__11327),
            .I(N__11268));
    Span4Mux_v I__2756 (
            .O(N__11324),
            .I(N__11265));
    Span4Mux_v I__2755 (
            .O(N__11321),
            .I(N__11262));
    Span12Mux_v I__2754 (
            .O(N__11316),
            .I(N__11259));
    Span12Mux_h I__2753 (
            .O(N__11309),
            .I(N__11254));
    Span12Mux_h I__2752 (
            .O(N__11306),
            .I(N__11254));
    Span12Mux_h I__2751 (
            .O(N__11303),
            .I(N__11251));
    Span12Mux_v I__2750 (
            .O(N__11300),
            .I(N__11246));
    Sp12to4 I__2749 (
            .O(N__11293),
            .I(N__11246));
    Span12Mux_h I__2748 (
            .O(N__11290),
            .I(N__11241));
    Span12Mux_h I__2747 (
            .O(N__11287),
            .I(N__11241));
    LocalMux I__2746 (
            .O(N__11284),
            .I(N__11238));
    Sp12to4 I__2745 (
            .O(N__11279),
            .I(N__11233));
    LocalMux I__2744 (
            .O(N__11276),
            .I(N__11233));
    Span4Mux_v I__2743 (
            .O(N__11271),
            .I(N__11230));
    Span4Mux_v I__2742 (
            .O(N__11268),
            .I(N__11227));
    IoSpan4Mux I__2741 (
            .O(N__11265),
            .I(N__11224));
    Span4Mux_v I__2740 (
            .O(N__11262),
            .I(N__11221));
    Span12Mux_h I__2739 (
            .O(N__11259),
            .I(N__11216));
    Span12Mux_v I__2738 (
            .O(N__11254),
            .I(N__11216));
    Span12Mux_v I__2737 (
            .O(N__11251),
            .I(N__11211));
    Span12Mux_h I__2736 (
            .O(N__11246),
            .I(N__11211));
    Span12Mux_v I__2735 (
            .O(N__11241),
            .I(N__11204));
    Span12Mux_h I__2734 (
            .O(N__11238),
            .I(N__11204));
    Span12Mux_h I__2733 (
            .O(N__11233),
            .I(N__11204));
    Span4Mux_h I__2732 (
            .O(N__11230),
            .I(N__11199));
    Span4Mux_h I__2731 (
            .O(N__11227),
            .I(N__11199));
    IoSpan4Mux I__2730 (
            .O(N__11224),
            .I(N__11194));
    IoSpan4Mux I__2729 (
            .O(N__11221),
            .I(N__11194));
    Odrv12 I__2728 (
            .O(N__11216),
            .I(TS_CPUn_c));
    Odrv12 I__2727 (
            .O(N__11211),
            .I(TS_CPUn_c));
    Odrv12 I__2726 (
            .O(N__11204),
            .I(TS_CPUn_c));
    Odrv4 I__2725 (
            .O(N__11199),
            .I(TS_CPUn_c));
    Odrv4 I__2724 (
            .O(N__11194),
            .I(TS_CPUn_c));
    CascadeMux I__2723 (
            .O(N__11183),
            .I(N__11178));
    CascadeMux I__2722 (
            .O(N__11182),
            .I(N__11175));
    InMux I__2721 (
            .O(N__11181),
            .I(N__11169));
    InMux I__2720 (
            .O(N__11178),
            .I(N__11169));
    InMux I__2719 (
            .O(N__11175),
            .I(N__11163));
    InMux I__2718 (
            .O(N__11174),
            .I(N__11158));
    LocalMux I__2717 (
            .O(N__11169),
            .I(N__11154));
    InMux I__2716 (
            .O(N__11168),
            .I(N__11151));
    CascadeMux I__2715 (
            .O(N__11167),
            .I(N__11145));
    CascadeMux I__2714 (
            .O(N__11166),
            .I(N__11139));
    LocalMux I__2713 (
            .O(N__11163),
            .I(N__11134));
    InMux I__2712 (
            .O(N__11162),
            .I(N__11127));
    InMux I__2711 (
            .O(N__11161),
            .I(N__11123));
    LocalMux I__2710 (
            .O(N__11158),
            .I(N__11120));
    InMux I__2709 (
            .O(N__11157),
            .I(N__11117));
    Span4Mux_v I__2708 (
            .O(N__11154),
            .I(N__11114));
    LocalMux I__2707 (
            .O(N__11151),
            .I(N__11110));
    InMux I__2706 (
            .O(N__11150),
            .I(N__11104));
    InMux I__2705 (
            .O(N__11149),
            .I(N__11104));
    InMux I__2704 (
            .O(N__11148),
            .I(N__11101));
    InMux I__2703 (
            .O(N__11145),
            .I(N__11098));
    InMux I__2702 (
            .O(N__11144),
            .I(N__11095));
    InMux I__2701 (
            .O(N__11143),
            .I(N__11092));
    InMux I__2700 (
            .O(N__11142),
            .I(N__11087));
    InMux I__2699 (
            .O(N__11139),
            .I(N__11087));
    InMux I__2698 (
            .O(N__11138),
            .I(N__11084));
    CascadeMux I__2697 (
            .O(N__11137),
            .I(N__11080));
    Span4Mux_h I__2696 (
            .O(N__11134),
            .I(N__11073));
    CascadeMux I__2695 (
            .O(N__11133),
            .I(N__11070));
    CascadeMux I__2694 (
            .O(N__11132),
            .I(N__11061));
    CascadeMux I__2693 (
            .O(N__11131),
            .I(N__11058));
    CascadeMux I__2692 (
            .O(N__11130),
            .I(N__11055));
    LocalMux I__2691 (
            .O(N__11127),
            .I(N__11050));
    InMux I__2690 (
            .O(N__11126),
            .I(N__11047));
    LocalMux I__2689 (
            .O(N__11123),
            .I(N__11044));
    Span4Mux_v I__2688 (
            .O(N__11120),
            .I(N__11039));
    LocalMux I__2687 (
            .O(N__11117),
            .I(N__11039));
    Span4Mux_v I__2686 (
            .O(N__11114),
            .I(N__11034));
    InMux I__2685 (
            .O(N__11113),
            .I(N__11031));
    Span4Mux_v I__2684 (
            .O(N__11110),
            .I(N__11028));
    InMux I__2683 (
            .O(N__11109),
            .I(N__11025));
    LocalMux I__2682 (
            .O(N__11104),
            .I(N__11016));
    LocalMux I__2681 (
            .O(N__11101),
            .I(N__11016));
    LocalMux I__2680 (
            .O(N__11098),
            .I(N__11016));
    LocalMux I__2679 (
            .O(N__11095),
            .I(N__11007));
    LocalMux I__2678 (
            .O(N__11092),
            .I(N__11007));
    LocalMux I__2677 (
            .O(N__11087),
            .I(N__11007));
    LocalMux I__2676 (
            .O(N__11084),
            .I(N__11007));
    InMux I__2675 (
            .O(N__11083),
            .I(N__11004));
    InMux I__2674 (
            .O(N__11080),
            .I(N__11001));
    InMux I__2673 (
            .O(N__11079),
            .I(N__10998));
    InMux I__2672 (
            .O(N__11078),
            .I(N__10995));
    InMux I__2671 (
            .O(N__11077),
            .I(N__10989));
    CascadeMux I__2670 (
            .O(N__11076),
            .I(N__10986));
    Span4Mux_v I__2669 (
            .O(N__11073),
            .I(N__10983));
    InMux I__2668 (
            .O(N__11070),
            .I(N__10980));
    CascadeMux I__2667 (
            .O(N__11069),
            .I(N__10977));
    CascadeMux I__2666 (
            .O(N__11068),
            .I(N__10974));
    CascadeMux I__2665 (
            .O(N__11067),
            .I(N__10970));
    InMux I__2664 (
            .O(N__11066),
            .I(N__10962));
    CascadeMux I__2663 (
            .O(N__11065),
            .I(N__10958));
    CascadeMux I__2662 (
            .O(N__11064),
            .I(N__10955));
    InMux I__2661 (
            .O(N__11061),
            .I(N__10946));
    InMux I__2660 (
            .O(N__11058),
            .I(N__10946));
    InMux I__2659 (
            .O(N__11055),
            .I(N__10946));
    InMux I__2658 (
            .O(N__11054),
            .I(N__10943));
    InMux I__2657 (
            .O(N__11053),
            .I(N__10940));
    Span4Mux_h I__2656 (
            .O(N__11050),
            .I(N__10935));
    LocalMux I__2655 (
            .O(N__11047),
            .I(N__10935));
    Span4Mux_v I__2654 (
            .O(N__11044),
            .I(N__10932));
    Span4Mux_h I__2653 (
            .O(N__11039),
            .I(N__10929));
    InMux I__2652 (
            .O(N__11038),
            .I(N__10926));
    InMux I__2651 (
            .O(N__11037),
            .I(N__10923));
    Span4Mux_h I__2650 (
            .O(N__11034),
            .I(N__10918));
    LocalMux I__2649 (
            .O(N__11031),
            .I(N__10918));
    Span4Mux_v I__2648 (
            .O(N__11028),
            .I(N__10913));
    LocalMux I__2647 (
            .O(N__11025),
            .I(N__10913));
    InMux I__2646 (
            .O(N__11024),
            .I(N__10908));
    InMux I__2645 (
            .O(N__11023),
            .I(N__10908));
    Span4Mux_v I__2644 (
            .O(N__11016),
            .I(N__10905));
    Span4Mux_v I__2643 (
            .O(N__11007),
            .I(N__10894));
    LocalMux I__2642 (
            .O(N__11004),
            .I(N__10894));
    LocalMux I__2641 (
            .O(N__11001),
            .I(N__10894));
    LocalMux I__2640 (
            .O(N__10998),
            .I(N__10894));
    LocalMux I__2639 (
            .O(N__10995),
            .I(N__10894));
    InMux I__2638 (
            .O(N__10994),
            .I(N__10891));
    InMux I__2637 (
            .O(N__10993),
            .I(N__10888));
    CascadeMux I__2636 (
            .O(N__10992),
            .I(N__10885));
    LocalMux I__2635 (
            .O(N__10989),
            .I(N__10880));
    InMux I__2634 (
            .O(N__10986),
            .I(N__10877));
    Span4Mux_v I__2633 (
            .O(N__10983),
            .I(N__10871));
    LocalMux I__2632 (
            .O(N__10980),
            .I(N__10871));
    InMux I__2631 (
            .O(N__10977),
            .I(N__10866));
    InMux I__2630 (
            .O(N__10974),
            .I(N__10866));
    InMux I__2629 (
            .O(N__10973),
            .I(N__10859));
    InMux I__2628 (
            .O(N__10970),
            .I(N__10859));
    InMux I__2627 (
            .O(N__10969),
            .I(N__10859));
    InMux I__2626 (
            .O(N__10968),
            .I(N__10856));
    CascadeMux I__2625 (
            .O(N__10967),
            .I(N__10848));
    CascadeMux I__2624 (
            .O(N__10966),
            .I(N__10844));
    CascadeMux I__2623 (
            .O(N__10965),
            .I(N__10840));
    LocalMux I__2622 (
            .O(N__10962),
            .I(N__10836));
    InMux I__2621 (
            .O(N__10961),
            .I(N__10831));
    InMux I__2620 (
            .O(N__10958),
            .I(N__10831));
    InMux I__2619 (
            .O(N__10955),
            .I(N__10828));
    CascadeMux I__2618 (
            .O(N__10954),
            .I(N__10825));
    CascadeMux I__2617 (
            .O(N__10953),
            .I(N__10821));
    LocalMux I__2616 (
            .O(N__10946),
            .I(N__10813));
    LocalMux I__2615 (
            .O(N__10943),
            .I(N__10813));
    LocalMux I__2614 (
            .O(N__10940),
            .I(N__10813));
    Span4Mux_v I__2613 (
            .O(N__10935),
            .I(N__10810));
    Span4Mux_h I__2612 (
            .O(N__10932),
            .I(N__10801));
    Span4Mux_v I__2611 (
            .O(N__10929),
            .I(N__10801));
    LocalMux I__2610 (
            .O(N__10926),
            .I(N__10801));
    LocalMux I__2609 (
            .O(N__10923),
            .I(N__10801));
    Span4Mux_v I__2608 (
            .O(N__10918),
            .I(N__10794));
    Span4Mux_v I__2607 (
            .O(N__10913),
            .I(N__10794));
    LocalMux I__2606 (
            .O(N__10908),
            .I(N__10794));
    Span4Mux_v I__2605 (
            .O(N__10905),
            .I(N__10785));
    Span4Mux_v I__2604 (
            .O(N__10894),
            .I(N__10785));
    LocalMux I__2603 (
            .O(N__10891),
            .I(N__10785));
    LocalMux I__2602 (
            .O(N__10888),
            .I(N__10785));
    InMux I__2601 (
            .O(N__10885),
            .I(N__10782));
    InMux I__2600 (
            .O(N__10884),
            .I(N__10779));
    InMux I__2599 (
            .O(N__10883),
            .I(N__10776));
    Span4Mux_h I__2598 (
            .O(N__10880),
            .I(N__10771));
    LocalMux I__2597 (
            .O(N__10877),
            .I(N__10771));
    InMux I__2596 (
            .O(N__10876),
            .I(N__10768));
    Span4Mux_h I__2595 (
            .O(N__10871),
            .I(N__10765));
    LocalMux I__2594 (
            .O(N__10866),
            .I(N__10758));
    LocalMux I__2593 (
            .O(N__10859),
            .I(N__10758));
    LocalMux I__2592 (
            .O(N__10856),
            .I(N__10758));
    InMux I__2591 (
            .O(N__10855),
            .I(N__10751));
    InMux I__2590 (
            .O(N__10854),
            .I(N__10751));
    InMux I__2589 (
            .O(N__10853),
            .I(N__10751));
    InMux I__2588 (
            .O(N__10852),
            .I(N__10746));
    InMux I__2587 (
            .O(N__10851),
            .I(N__10746));
    InMux I__2586 (
            .O(N__10848),
            .I(N__10737));
    InMux I__2585 (
            .O(N__10847),
            .I(N__10737));
    InMux I__2584 (
            .O(N__10844),
            .I(N__10737));
    InMux I__2583 (
            .O(N__10843),
            .I(N__10737));
    InMux I__2582 (
            .O(N__10840),
            .I(N__10732));
    InMux I__2581 (
            .O(N__10839),
            .I(N__10732));
    Span4Mux_v I__2580 (
            .O(N__10836),
            .I(N__10725));
    LocalMux I__2579 (
            .O(N__10831),
            .I(N__10725));
    LocalMux I__2578 (
            .O(N__10828),
            .I(N__10725));
    InMux I__2577 (
            .O(N__10825),
            .I(N__10718));
    InMux I__2576 (
            .O(N__10824),
            .I(N__10718));
    InMux I__2575 (
            .O(N__10821),
            .I(N__10718));
    CascadeMux I__2574 (
            .O(N__10820),
            .I(N__10715));
    Span4Mux_v I__2573 (
            .O(N__10813),
            .I(N__10712));
    Span4Mux_h I__2572 (
            .O(N__10810),
            .I(N__10707));
    Span4Mux_v I__2571 (
            .O(N__10801),
            .I(N__10707));
    Span4Mux_v I__2570 (
            .O(N__10794),
            .I(N__10704));
    Span4Mux_v I__2569 (
            .O(N__10785),
            .I(N__10694));
    LocalMux I__2568 (
            .O(N__10782),
            .I(N__10694));
    LocalMux I__2567 (
            .O(N__10779),
            .I(N__10694));
    LocalMux I__2566 (
            .O(N__10776),
            .I(N__10694));
    Span4Mux_v I__2565 (
            .O(N__10771),
            .I(N__10690));
    LocalMux I__2564 (
            .O(N__10768),
            .I(N__10687));
    Span4Mux_v I__2563 (
            .O(N__10765),
            .I(N__10683));
    Span12Mux_s11_v I__2562 (
            .O(N__10758),
            .I(N__10672));
    LocalMux I__2561 (
            .O(N__10751),
            .I(N__10672));
    LocalMux I__2560 (
            .O(N__10746),
            .I(N__10672));
    LocalMux I__2559 (
            .O(N__10737),
            .I(N__10672));
    LocalMux I__2558 (
            .O(N__10732),
            .I(N__10672));
    Span4Mux_v I__2557 (
            .O(N__10725),
            .I(N__10669));
    LocalMux I__2556 (
            .O(N__10718),
            .I(N__10666));
    InMux I__2555 (
            .O(N__10715),
            .I(N__10663));
    Sp12to4 I__2554 (
            .O(N__10712),
            .I(N__10658));
    Sp12to4 I__2553 (
            .O(N__10707),
            .I(N__10658));
    Span4Mux_v I__2552 (
            .O(N__10704),
            .I(N__10655));
    InMux I__2551 (
            .O(N__10703),
            .I(N__10652));
    Span4Mux_v I__2550 (
            .O(N__10694),
            .I(N__10649));
    InMux I__2549 (
            .O(N__10693),
            .I(N__10646));
    Span4Mux_h I__2548 (
            .O(N__10690),
            .I(N__10643));
    Span4Mux_v I__2547 (
            .O(N__10687),
            .I(N__10640));
    InMux I__2546 (
            .O(N__10686),
            .I(N__10637));
    Span4Mux_v I__2545 (
            .O(N__10683),
            .I(N__10634));
    Span12Mux_v I__2544 (
            .O(N__10672),
            .I(N__10625));
    Sp12to4 I__2543 (
            .O(N__10669),
            .I(N__10625));
    Span12Mux_s8_v I__2542 (
            .O(N__10666),
            .I(N__10625));
    LocalMux I__2541 (
            .O(N__10663),
            .I(N__10625));
    Span12Mux_h I__2540 (
            .O(N__10658),
            .I(N__10622));
    Sp12to4 I__2539 (
            .O(N__10655),
            .I(N__10613));
    LocalMux I__2538 (
            .O(N__10652),
            .I(N__10613));
    Sp12to4 I__2537 (
            .O(N__10649),
            .I(N__10613));
    LocalMux I__2536 (
            .O(N__10646),
            .I(N__10613));
    Span4Mux_h I__2535 (
            .O(N__10643),
            .I(N__10606));
    Span4Mux_v I__2534 (
            .O(N__10640),
            .I(N__10606));
    LocalMux I__2533 (
            .O(N__10637),
            .I(N__10606));
    Span4Mux_v I__2532 (
            .O(N__10634),
            .I(N__10603));
    Span12Mux_h I__2531 (
            .O(N__10625),
            .I(N__10596));
    Span12Mux_v I__2530 (
            .O(N__10622),
            .I(N__10596));
    Span12Mux_h I__2529 (
            .O(N__10613),
            .I(N__10596));
    Span4Mux_v I__2528 (
            .O(N__10606),
            .I(N__10593));
    Odrv4 I__2527 (
            .O(N__10603),
            .I(LBENn_c));
    Odrv12 I__2526 (
            .O(N__10596),
            .I(LBENn_c));
    Odrv4 I__2525 (
            .O(N__10593),
            .I(LBENn_c));
    InMux I__2524 (
            .O(N__10586),
            .I(N__10577));
    CascadeMux I__2523 (
            .O(N__10585),
            .I(N__10574));
    InMux I__2522 (
            .O(N__10584),
            .I(N__10564));
    InMux I__2521 (
            .O(N__10583),
            .I(N__10561));
    InMux I__2520 (
            .O(N__10582),
            .I(N__10558));
    InMux I__2519 (
            .O(N__10581),
            .I(N__10555));
    IoInMux I__2518 (
            .O(N__10580),
            .I(N__10551));
    LocalMux I__2517 (
            .O(N__10577),
            .I(N__10545));
    InMux I__2516 (
            .O(N__10574),
            .I(N__10542));
    InMux I__2515 (
            .O(N__10573),
            .I(N__10539));
    CascadeMux I__2514 (
            .O(N__10572),
            .I(N__10536));
    InMux I__2513 (
            .O(N__10571),
            .I(N__10532));
    CascadeMux I__2512 (
            .O(N__10570),
            .I(N__10529));
    InMux I__2511 (
            .O(N__10569),
            .I(N__10524));
    CascadeMux I__2510 (
            .O(N__10568),
            .I(N__10521));
    InMux I__2509 (
            .O(N__10567),
            .I(N__10518));
    LocalMux I__2508 (
            .O(N__10564),
            .I(N__10511));
    LocalMux I__2507 (
            .O(N__10561),
            .I(N__10511));
    LocalMux I__2506 (
            .O(N__10558),
            .I(N__10511));
    LocalMux I__2505 (
            .O(N__10555),
            .I(N__10508));
    InMux I__2504 (
            .O(N__10554),
            .I(N__10505));
    LocalMux I__2503 (
            .O(N__10551),
            .I(N__10499));
    CascadeMux I__2502 (
            .O(N__10550),
            .I(N__10495));
    CascadeMux I__2501 (
            .O(N__10549),
            .I(N__10490));
    CascadeMux I__2500 (
            .O(N__10548),
            .I(N__10487));
    Span4Mux_v I__2499 (
            .O(N__10545),
            .I(N__10478));
    LocalMux I__2498 (
            .O(N__10542),
            .I(N__10478));
    LocalMux I__2497 (
            .O(N__10539),
            .I(N__10478));
    InMux I__2496 (
            .O(N__10536),
            .I(N__10473));
    InMux I__2495 (
            .O(N__10535),
            .I(N__10473));
    LocalMux I__2494 (
            .O(N__10532),
            .I(N__10470));
    InMux I__2493 (
            .O(N__10529),
            .I(N__10465));
    InMux I__2492 (
            .O(N__10528),
            .I(N__10465));
    InMux I__2491 (
            .O(N__10527),
            .I(N__10462));
    LocalMux I__2490 (
            .O(N__10524),
            .I(N__10458));
    InMux I__2489 (
            .O(N__10521),
            .I(N__10455));
    LocalMux I__2488 (
            .O(N__10518),
            .I(N__10451));
    Span4Mux_v I__2487 (
            .O(N__10511),
            .I(N__10434));
    Span4Mux_h I__2486 (
            .O(N__10508),
            .I(N__10434));
    LocalMux I__2485 (
            .O(N__10505),
            .I(N__10434));
    InMux I__2484 (
            .O(N__10504),
            .I(N__10431));
    InMux I__2483 (
            .O(N__10503),
            .I(N__10428));
    InMux I__2482 (
            .O(N__10502),
            .I(N__10425));
    Span4Mux_s3_v I__2481 (
            .O(N__10499),
            .I(N__10422));
    InMux I__2480 (
            .O(N__10498),
            .I(N__10419));
    InMux I__2479 (
            .O(N__10495),
            .I(N__10416));
    InMux I__2478 (
            .O(N__10494),
            .I(N__10411));
    InMux I__2477 (
            .O(N__10493),
            .I(N__10411));
    InMux I__2476 (
            .O(N__10490),
            .I(N__10406));
    InMux I__2475 (
            .O(N__10487),
            .I(N__10406));
    InMux I__2474 (
            .O(N__10486),
            .I(N__10403));
    InMux I__2473 (
            .O(N__10485),
            .I(N__10400));
    Span4Mux_v I__2472 (
            .O(N__10478),
            .I(N__10395));
    LocalMux I__2471 (
            .O(N__10473),
            .I(N__10395));
    Span4Mux_v I__2470 (
            .O(N__10470),
            .I(N__10392));
    LocalMux I__2469 (
            .O(N__10465),
            .I(N__10389));
    LocalMux I__2468 (
            .O(N__10462),
            .I(N__10386));
    InMux I__2467 (
            .O(N__10461),
            .I(N__10383));
    Span4Mux_v I__2466 (
            .O(N__10458),
            .I(N__10376));
    LocalMux I__2465 (
            .O(N__10455),
            .I(N__10376));
    CascadeMux I__2464 (
            .O(N__10454),
            .I(N__10373));
    Span4Mux_v I__2463 (
            .O(N__10451),
            .I(N__10369));
    InMux I__2462 (
            .O(N__10450),
            .I(N__10366));
    InMux I__2461 (
            .O(N__10449),
            .I(N__10361));
    InMux I__2460 (
            .O(N__10448),
            .I(N__10361));
    CascadeMux I__2459 (
            .O(N__10447),
            .I(N__10358));
    CascadeMux I__2458 (
            .O(N__10446),
            .I(N__10355));
    CascadeMux I__2457 (
            .O(N__10445),
            .I(N__10352));
    InMux I__2456 (
            .O(N__10444),
            .I(N__10347));
    InMux I__2455 (
            .O(N__10443),
            .I(N__10340));
    InMux I__2454 (
            .O(N__10442),
            .I(N__10340));
    InMux I__2453 (
            .O(N__10441),
            .I(N__10340));
    Span4Mux_v I__2452 (
            .O(N__10434),
            .I(N__10327));
    LocalMux I__2451 (
            .O(N__10431),
            .I(N__10327));
    LocalMux I__2450 (
            .O(N__10428),
            .I(N__10327));
    LocalMux I__2449 (
            .O(N__10425),
            .I(N__10327));
    Span4Mux_v I__2448 (
            .O(N__10422),
            .I(N__10312));
    LocalMux I__2447 (
            .O(N__10419),
            .I(N__10312));
    LocalMux I__2446 (
            .O(N__10416),
            .I(N__10312));
    LocalMux I__2445 (
            .O(N__10411),
            .I(N__10312));
    LocalMux I__2444 (
            .O(N__10406),
            .I(N__10312));
    LocalMux I__2443 (
            .O(N__10403),
            .I(N__10312));
    LocalMux I__2442 (
            .O(N__10400),
            .I(N__10312));
    Span4Mux_v I__2441 (
            .O(N__10395),
            .I(N__10309));
    Span4Mux_h I__2440 (
            .O(N__10392),
            .I(N__10300));
    Span4Mux_v I__2439 (
            .O(N__10389),
            .I(N__10300));
    Span4Mux_h I__2438 (
            .O(N__10386),
            .I(N__10300));
    LocalMux I__2437 (
            .O(N__10383),
            .I(N__10300));
    InMux I__2436 (
            .O(N__10382),
            .I(N__10297));
    InMux I__2435 (
            .O(N__10381),
            .I(N__10294));
    Span4Mux_v I__2434 (
            .O(N__10376),
            .I(N__10291));
    InMux I__2433 (
            .O(N__10373),
            .I(N__10288));
    CascadeMux I__2432 (
            .O(N__10372),
            .I(N__10285));
    Span4Mux_h I__2431 (
            .O(N__10369),
            .I(N__10282));
    LocalMux I__2430 (
            .O(N__10366),
            .I(N__10277));
    LocalMux I__2429 (
            .O(N__10361),
            .I(N__10277));
    InMux I__2428 (
            .O(N__10358),
            .I(N__10274));
    InMux I__2427 (
            .O(N__10355),
            .I(N__10271));
    InMux I__2426 (
            .O(N__10352),
            .I(N__10268));
    CascadeMux I__2425 (
            .O(N__10351),
            .I(N__10265));
    CascadeMux I__2424 (
            .O(N__10350),
            .I(N__10262));
    LocalMux I__2423 (
            .O(N__10347),
            .I(N__10257));
    LocalMux I__2422 (
            .O(N__10340),
            .I(N__10257));
    InMux I__2421 (
            .O(N__10339),
            .I(N__10252));
    InMux I__2420 (
            .O(N__10338),
            .I(N__10252));
    CascadeMux I__2419 (
            .O(N__10337),
            .I(N__10245));
    CascadeMux I__2418 (
            .O(N__10336),
            .I(N__10242));
    Span4Mux_v I__2417 (
            .O(N__10327),
            .I(N__10227));
    Span4Mux_v I__2416 (
            .O(N__10312),
            .I(N__10227));
    Span4Mux_h I__2415 (
            .O(N__10309),
            .I(N__10222));
    Span4Mux_v I__2414 (
            .O(N__10300),
            .I(N__10222));
    LocalMux I__2413 (
            .O(N__10297),
            .I(N__10217));
    LocalMux I__2412 (
            .O(N__10294),
            .I(N__10217));
    Span4Mux_h I__2411 (
            .O(N__10291),
            .I(N__10212));
    LocalMux I__2410 (
            .O(N__10288),
            .I(N__10212));
    InMux I__2409 (
            .O(N__10285),
            .I(N__10209));
    Span4Mux_h I__2408 (
            .O(N__10282),
            .I(N__10206));
    Span4Mux_v I__2407 (
            .O(N__10277),
            .I(N__10201));
    LocalMux I__2406 (
            .O(N__10274),
            .I(N__10201));
    LocalMux I__2405 (
            .O(N__10271),
            .I(N__10196));
    LocalMux I__2404 (
            .O(N__10268),
            .I(N__10196));
    InMux I__2403 (
            .O(N__10265),
            .I(N__10193));
    InMux I__2402 (
            .O(N__10262),
            .I(N__10190));
    Span4Mux_h I__2401 (
            .O(N__10257),
            .I(N__10185));
    LocalMux I__2400 (
            .O(N__10252),
            .I(N__10185));
    InMux I__2399 (
            .O(N__10251),
            .I(N__10176));
    InMux I__2398 (
            .O(N__10250),
            .I(N__10176));
    InMux I__2397 (
            .O(N__10249),
            .I(N__10176));
    InMux I__2396 (
            .O(N__10248),
            .I(N__10176));
    InMux I__2395 (
            .O(N__10245),
            .I(N__10171));
    InMux I__2394 (
            .O(N__10242),
            .I(N__10171));
    CascadeMux I__2393 (
            .O(N__10241),
            .I(N__10167));
    CascadeMux I__2392 (
            .O(N__10240),
            .I(N__10164));
    InMux I__2391 (
            .O(N__10239),
            .I(N__10157));
    InMux I__2390 (
            .O(N__10238),
            .I(N__10157));
    InMux I__2389 (
            .O(N__10237),
            .I(N__10157));
    InMux I__2388 (
            .O(N__10236),
            .I(N__10152));
    InMux I__2387 (
            .O(N__10235),
            .I(N__10152));
    CascadeMux I__2386 (
            .O(N__10234),
            .I(N__10149));
    CascadeMux I__2385 (
            .O(N__10233),
            .I(N__10145));
    CascadeMux I__2384 (
            .O(N__10232),
            .I(N__10142));
    Sp12to4 I__2383 (
            .O(N__10227),
            .I(N__10137));
    Sp12to4 I__2382 (
            .O(N__10222),
            .I(N__10137));
    Span12Mux_s11_h I__2381 (
            .O(N__10217),
            .I(N__10134));
    Sp12to4 I__2380 (
            .O(N__10212),
            .I(N__10131));
    LocalMux I__2379 (
            .O(N__10209),
            .I(N__10128));
    Span4Mux_h I__2378 (
            .O(N__10206),
            .I(N__10123));
    Span4Mux_v I__2377 (
            .O(N__10201),
            .I(N__10123));
    Span4Mux_h I__2376 (
            .O(N__10196),
            .I(N__10116));
    LocalMux I__2375 (
            .O(N__10193),
            .I(N__10116));
    LocalMux I__2374 (
            .O(N__10190),
            .I(N__10116));
    Span4Mux_v I__2373 (
            .O(N__10185),
            .I(N__10111));
    LocalMux I__2372 (
            .O(N__10176),
            .I(N__10111));
    LocalMux I__2371 (
            .O(N__10171),
            .I(N__10108));
    InMux I__2370 (
            .O(N__10170),
            .I(N__10101));
    InMux I__2369 (
            .O(N__10167),
            .I(N__10101));
    InMux I__2368 (
            .O(N__10164),
            .I(N__10101));
    LocalMux I__2367 (
            .O(N__10157),
            .I(N__10098));
    LocalMux I__2366 (
            .O(N__10152),
            .I(N__10095));
    InMux I__2365 (
            .O(N__10149),
            .I(N__10088));
    InMux I__2364 (
            .O(N__10148),
            .I(N__10088));
    InMux I__2363 (
            .O(N__10145),
            .I(N__10088));
    InMux I__2362 (
            .O(N__10142),
            .I(N__10085));
    Span12Mux_h I__2361 (
            .O(N__10137),
            .I(N__10082));
    Span12Mux_h I__2360 (
            .O(N__10134),
            .I(N__10079));
    Span12Mux_s11_v I__2359 (
            .O(N__10131),
            .I(N__10074));
    Span12Mux_s11_h I__2358 (
            .O(N__10128),
            .I(N__10074));
    Span4Mux_v I__2357 (
            .O(N__10123),
            .I(N__10069));
    Span4Mux_v I__2356 (
            .O(N__10116),
            .I(N__10069));
    Span4Mux_v I__2355 (
            .O(N__10111),
            .I(N__10062));
    Span4Mux_h I__2354 (
            .O(N__10108),
            .I(N__10062));
    LocalMux I__2353 (
            .O(N__10101),
            .I(N__10062));
    Span4Mux_h I__2352 (
            .O(N__10098),
            .I(N__10053));
    Span4Mux_v I__2351 (
            .O(N__10095),
            .I(N__10053));
    LocalMux I__2350 (
            .O(N__10088),
            .I(N__10053));
    LocalMux I__2349 (
            .O(N__10085),
            .I(N__10053));
    Span12Mux_h I__2348 (
            .O(N__10082),
            .I(N__10050));
    Span12Mux_v I__2347 (
            .O(N__10079),
            .I(N__10045));
    Span12Mux_h I__2346 (
            .O(N__10074),
            .I(N__10045));
    Span4Mux_h I__2345 (
            .O(N__10069),
            .I(N__10042));
    Span4Mux_v I__2344 (
            .O(N__10062),
            .I(N__10037));
    Span4Mux_v I__2343 (
            .O(N__10053),
            .I(N__10037));
    Odrv12 I__2342 (
            .O(N__10050),
            .I(RnW_c));
    Odrv12 I__2341 (
            .O(N__10045),
            .I(RnW_c));
    Odrv4 I__2340 (
            .O(N__10042),
            .I(RnW_c));
    Odrv4 I__2339 (
            .O(N__10037),
            .I(RnW_c));
    InMux I__2338 (
            .O(N__10028),
            .I(N__10025));
    LocalMux I__2337 (
            .O(N__10025),
            .I(READ_CYCLE_ACTIVE_rep12_i_ess));
    InMux I__2336 (
            .O(N__10022),
            .I(N__10019));
    LocalMux I__2335 (
            .O(N__10019),
            .I(READ_CYCLE_ACTIVE_rep29_i_ess));
    IoInMux I__2334 (
            .O(N__10016),
            .I(N__10013));
    LocalMux I__2333 (
            .O(N__10013),
            .I(N__10010));
    Span4Mux_s3_h I__2332 (
            .O(N__10010),
            .I(N__10007));
    Odrv4 I__2331 (
            .O(N__10007),
            .I(N_195_i));
    InMux I__2330 (
            .O(N__10004),
            .I(N__10001));
    LocalMux I__2329 (
            .O(N__10001),
            .I(READ_CYCLE_ACTIVE_rep14_i_ess));
    InMux I__2328 (
            .O(N__9998),
            .I(N__9995));
    LocalMux I__2327 (
            .O(N__9995),
            .I(READ_CYCLE_ACTIVE_rep22_i_ess));
    IoInMux I__2326 (
            .O(N__9992),
            .I(N__9989));
    LocalMux I__2325 (
            .O(N__9989),
            .I(N__9986));
    Span4Mux_s3_h I__2324 (
            .O(N__9986),
            .I(N__9983));
    Odrv4 I__2323 (
            .O(N__9983),
            .I(N_203_i));
    InMux I__2322 (
            .O(N__9980),
            .I(N__9977));
    LocalMux I__2321 (
            .O(N__9977),
            .I(N__9974));
    Odrv4 I__2320 (
            .O(N__9974),
            .I(READ_CYCLE_ACTIVE_rep23_i_ess));
    IoInMux I__2319 (
            .O(N__9971),
            .I(N__9968));
    LocalMux I__2318 (
            .O(N__9968),
            .I(N__9965));
    IoSpan4Mux I__2317 (
            .O(N__9965),
            .I(N__9962));
    Span4Mux_s3_h I__2316 (
            .O(N__9962),
            .I(N__9959));
    Odrv4 I__2315 (
            .O(N__9959),
            .I(N_204_i));
    InMux I__2314 (
            .O(N__9956),
            .I(N__9953));
    LocalMux I__2313 (
            .O(N__9953),
            .I(READ_CYCLE_ACTIVE_rep9_i_ess));
    IoInMux I__2312 (
            .O(N__9950),
            .I(N__9947));
    LocalMux I__2311 (
            .O(N__9947),
            .I(N__9944));
    Span4Mux_s3_h I__2310 (
            .O(N__9944),
            .I(N__9941));
    Span4Mux_v I__2309 (
            .O(N__9941),
            .I(N__9938));
    Odrv4 I__2308 (
            .O(N__9938),
            .I(N_190_i));
    InMux I__2307 (
            .O(N__9935),
            .I(N__9932));
    LocalMux I__2306 (
            .O(N__9932),
            .I(READ_CYCLE_ACTIVE_rep16_i_ess));
    InMux I__2305 (
            .O(N__9929),
            .I(N__9926));
    LocalMux I__2304 (
            .O(N__9926),
            .I(READ_CYCLE_ACTIVE_rep20_i_ess));
    IoInMux I__2303 (
            .O(N__9923),
            .I(N__9920));
    LocalMux I__2302 (
            .O(N__9920),
            .I(N__9917));
    Span4Mux_s3_h I__2301 (
            .O(N__9917),
            .I(N__9914));
    Odrv4 I__2300 (
            .O(N__9914),
            .I(N_201_i));
    InMux I__2299 (
            .O(N__9911),
            .I(N__9908));
    LocalMux I__2298 (
            .O(N__9908),
            .I(READ_CYCLE_ACTIVE_rep8_i_ess));
    IoInMux I__2297 (
            .O(N__9905),
            .I(N__9902));
    LocalMux I__2296 (
            .O(N__9902),
            .I(N__9899));
    Odrv12 I__2295 (
            .O(N__9899),
            .I(N_189_i));
    InMux I__2294 (
            .O(N__9896),
            .I(N__9893));
    LocalMux I__2293 (
            .O(N__9893),
            .I(READ_CYCLE_ACTIVE_rep21_i_ess));
    IoInMux I__2292 (
            .O(N__9890),
            .I(N__9887));
    LocalMux I__2291 (
            .O(N__9887),
            .I(N__9884));
    IoSpan4Mux I__2290 (
            .O(N__9884),
            .I(N__9881));
    Span4Mux_s3_h I__2289 (
            .O(N__9881),
            .I(N__9878));
    Odrv4 I__2288 (
            .O(N__9878),
            .I(N_202_i));
    IoInMux I__2287 (
            .O(N__9875),
            .I(N__9872));
    LocalMux I__2286 (
            .O(N__9872),
            .I(N__9869));
    Span12Mux_s11_h I__2285 (
            .O(N__9869),
            .I(N__9866));
    Span12Mux_v I__2284 (
            .O(N__9866),
            .I(N__9863));
    Odrv12 I__2283 (
            .O(N__9863),
            .I(N_210_i));
    IoInMux I__2282 (
            .O(N__9860),
            .I(N__9857));
    LocalMux I__2281 (
            .O(N__9857),
            .I(N__9854));
    Odrv12 I__2280 (
            .O(N__9854),
            .I(N_191_i));
    InMux I__2279 (
            .O(N__9851),
            .I(N__9848));
    LocalMux I__2278 (
            .O(N__9848),
            .I(READ_CYCLE_ACTIVE_rep10_i_ess));
    InMux I__2277 (
            .O(N__9845),
            .I(N__9842));
    LocalMux I__2276 (
            .O(N__9842),
            .I(READ_CYCLE_ACTIVE_rep26_i_ess));
    IoInMux I__2275 (
            .O(N__9839),
            .I(N__9836));
    LocalMux I__2274 (
            .O(N__9836),
            .I(N__9833));
    Span4Mux_s3_h I__2273 (
            .O(N__9833),
            .I(N__9830));
    Span4Mux_v I__2272 (
            .O(N__9830),
            .I(N__9827));
    Odrv4 I__2271 (
            .O(N__9827),
            .I(N_207_i));
    InMux I__2270 (
            .O(N__9824),
            .I(N__9821));
    LocalMux I__2269 (
            .O(N__9821),
            .I(READ_CYCLE_ACTIVE_rep30_i_ess));
    InMux I__2268 (
            .O(N__9818),
            .I(N__9815));
    LocalMux I__2267 (
            .O(N__9815),
            .I(READ_CYCLE_ACTIVE_rep17_i_ess));
    IoInMux I__2266 (
            .O(N__9812),
            .I(N__9809));
    LocalMux I__2265 (
            .O(N__9809),
            .I(N__9806));
    Span4Mux_s3_h I__2264 (
            .O(N__9806),
            .I(N__9803));
    Span4Mux_v I__2263 (
            .O(N__9803),
            .I(N__9800));
    Odrv4 I__2262 (
            .O(N__9800),
            .I(N_198_i));
    InMux I__2261 (
            .O(N__9797),
            .I(N__9794));
    LocalMux I__2260 (
            .O(N__9794),
            .I(READ_CYCLE_ACTIVE_rep18_i_ess));
    IoInMux I__2259 (
            .O(N__9791),
            .I(N__9788));
    LocalMux I__2258 (
            .O(N__9788),
            .I(N__9785));
    Span12Mux_s4_h I__2257 (
            .O(N__9785),
            .I(N__9782));
    Odrv12 I__2256 (
            .O(N__9782),
            .I(N_199_i));
    InMux I__2255 (
            .O(N__9779),
            .I(N__9776));
    LocalMux I__2254 (
            .O(N__9776),
            .I(READ_CYCLE_ACTIVE_rep31_i_ess));
    IoInMux I__2253 (
            .O(N__9773),
            .I(N__9770));
    LocalMux I__2252 (
            .O(N__9770),
            .I(N__9767));
    Span4Mux_s3_h I__2251 (
            .O(N__9767),
            .I(N__9764));
    Span4Mux_v I__2250 (
            .O(N__9764),
            .I(N__9761));
    Odrv4 I__2249 (
            .O(N__9761),
            .I(N_212_i));
    IoInMux I__2248 (
            .O(N__9758),
            .I(N__9755));
    LocalMux I__2247 (
            .O(N__9755),
            .I(N__9752));
    Span4Mux_s3_h I__2246 (
            .O(N__9752),
            .I(N__9749));
    Span4Mux_v I__2245 (
            .O(N__9749),
            .I(N__9746));
    Odrv4 I__2244 (
            .O(N__9746),
            .I(N_197_i));
    IoInMux I__2243 (
            .O(N__9743),
            .I(N__9740));
    LocalMux I__2242 (
            .O(N__9740),
            .I(N__9737));
    Span4Mux_s3_h I__2241 (
            .O(N__9737),
            .I(N__9734));
    Odrv4 I__2240 (
            .O(N__9734),
            .I(N_200_i));
    InMux I__2239 (
            .O(N__9731),
            .I(N__9728));
    LocalMux I__2238 (
            .O(N__9728),
            .I(READ_CYCLE_ACTIVE_rep19_i_ess));
    IoInMux I__2237 (
            .O(N__9725),
            .I(N__9722));
    LocalMux I__2236 (
            .O(N__9722),
            .I(N__9719));
    Span4Mux_s3_v I__2235 (
            .O(N__9719),
            .I(N__9716));
    Span4Mux_h I__2234 (
            .O(N__9716),
            .I(N__9713));
    Odrv4 I__2233 (
            .O(N__9713),
            .I(N_193_i));
    IoInMux I__2232 (
            .O(N__9710),
            .I(N__9707));
    LocalMux I__2231 (
            .O(N__9707),
            .I(N__9704));
    Span4Mux_s2_v I__2230 (
            .O(N__9704),
            .I(N__9701));
    Span4Mux_v I__2229 (
            .O(N__9701),
            .I(N__9698));
    Odrv4 I__2228 (
            .O(N__9698),
            .I(N_194_i));
    IoInMux I__2227 (
            .O(N__9695),
            .I(N__9692));
    LocalMux I__2226 (
            .O(N__9692),
            .I(N__9689));
    Span4Mux_s3_h I__2225 (
            .O(N__9689),
            .I(N__9686));
    Span4Mux_v I__2224 (
            .O(N__9686),
            .I(N__9683));
    Odrv4 I__2223 (
            .O(N__9683),
            .I(N_205_i));
    IoInMux I__2222 (
            .O(N__9680),
            .I(N__9677));
    LocalMux I__2221 (
            .O(N__9677),
            .I(N__9674));
    IoSpan4Mux I__2220 (
            .O(N__9674),
            .I(N__9671));
    Span4Mux_s3_h I__2219 (
            .O(N__9671),
            .I(N__9668));
    Odrv4 I__2218 (
            .O(N__9668),
            .I(N_206_i));
    IoInMux I__2217 (
            .O(N__9665),
            .I(N__9662));
    LocalMux I__2216 (
            .O(N__9662),
            .I(N__9659));
    Span4Mux_s3_h I__2215 (
            .O(N__9659),
            .I(N__9656));
    Span4Mux_v I__2214 (
            .O(N__9656),
            .I(N__9653));
    Odrv4 I__2213 (
            .O(N__9653),
            .I(N_208_i));
    InMux I__2212 (
            .O(N__9650),
            .I(N__9647));
    LocalMux I__2211 (
            .O(N__9647),
            .I(READ_CYCLE_ACTIVE_rep25_i_ess));
    InMux I__2210 (
            .O(N__9644),
            .I(N__9641));
    LocalMux I__2209 (
            .O(N__9641),
            .I(READ_CYCLE_ACTIVE_rep24_i_ess));
    InMux I__2208 (
            .O(N__9638),
            .I(N__9635));
    LocalMux I__2207 (
            .O(N__9635),
            .I(READ_CYCLE_ACTIVE_rep27_i_ess));
    IoInMux I__2206 (
            .O(N__9632),
            .I(N__9629));
    LocalMux I__2205 (
            .O(N__9629),
            .I(N__9626));
    Span4Mux_s3_h I__2204 (
            .O(N__9626),
            .I(N__9623));
    Span4Mux_v I__2203 (
            .O(N__9623),
            .I(N__9620));
    Odrv4 I__2202 (
            .O(N__9620),
            .I(N_211_i));
    IoInMux I__2201 (
            .O(N__9617),
            .I(N__9613));
    IoInMux I__2200 (
            .O(N__9616),
            .I(N__9610));
    LocalMux I__2199 (
            .O(N__9613),
            .I(N__9607));
    LocalMux I__2198 (
            .O(N__9610),
            .I(N__9603));
    IoSpan4Mux I__2197 (
            .O(N__9607),
            .I(N__9600));
    IoInMux I__2196 (
            .O(N__9606),
            .I(N__9597));
    IoSpan4Mux I__2195 (
            .O(N__9603),
            .I(N__9593));
    IoSpan4Mux I__2194 (
            .O(N__9600),
            .I(N__9588));
    LocalMux I__2193 (
            .O(N__9597),
            .I(N__9588));
    IoInMux I__2192 (
            .O(N__9596),
            .I(N__9585));
    Sp12to4 I__2191 (
            .O(N__9593),
            .I(N__9582));
    IoSpan4Mux I__2190 (
            .O(N__9588),
            .I(N__9579));
    LocalMux I__2189 (
            .O(N__9585),
            .I(N__9576));
    Span12Mux_s6_h I__2188 (
            .O(N__9582),
            .I(N__9573));
    Span4Mux_s3_v I__2187 (
            .O(N__9579),
            .I(N__9570));
    IoSpan4Mux I__2186 (
            .O(N__9576),
            .I(N__9567));
    Span12Mux_h I__2185 (
            .O(N__9573),
            .I(N__9564));
    Sp12to4 I__2184 (
            .O(N__9570),
            .I(N__9561));
    Span4Mux_s3_h I__2183 (
            .O(N__9567),
            .I(N__9558));
    Odrv12 I__2182 (
            .O(N__9564),
            .I(GB_BUFFER_CLK40_THRU_CO));
    Odrv12 I__2181 (
            .O(N__9561),
            .I(GB_BUFFER_CLK40_THRU_CO));
    Odrv4 I__2180 (
            .O(N__9558),
            .I(GB_BUFFER_CLK40_THRU_CO));
    InMux I__2179 (
            .O(N__9551),
            .I(N__9548));
    LocalMux I__2178 (
            .O(N__9548),
            .I(READ_CYCLE_ACTIVE_rep5_i_ess));
    IoInMux I__2177 (
            .O(N__9545),
            .I(N__9542));
    LocalMux I__2176 (
            .O(N__9542),
            .I(N__9539));
    Span4Mux_s2_v I__2175 (
            .O(N__9539),
            .I(N__9536));
    Span4Mux_v I__2174 (
            .O(N__9536),
            .I(N__9533));
    Odrv4 I__2173 (
            .O(N__9533),
            .I(N_186_i));
    InMux I__2172 (
            .O(N__9530),
            .I(N__9527));
    LocalMux I__2171 (
            .O(N__9527),
            .I(READ_CYCLE_ACTIVE_rep6_i_ess));
    IoInMux I__2170 (
            .O(N__9524),
            .I(N__9521));
    LocalMux I__2169 (
            .O(N__9521),
            .I(N__9518));
    Span4Mux_s2_v I__2168 (
            .O(N__9518),
            .I(N__9515));
    Span4Mux_v I__2167 (
            .O(N__9515),
            .I(N__9512));
    Odrv4 I__2166 (
            .O(N__9512),
            .I(N_187_i));
    InMux I__2165 (
            .O(N__9509),
            .I(N__9506));
    LocalMux I__2164 (
            .O(N__9506),
            .I(READ_CYCLE_ACTIVE_rep4_i_ess));
    IoInMux I__2163 (
            .O(N__9503),
            .I(N__9500));
    LocalMux I__2162 (
            .O(N__9500),
            .I(N__9497));
    Span4Mux_s2_v I__2161 (
            .O(N__9497),
            .I(N__9494));
    Span4Mux_v I__2160 (
            .O(N__9494),
            .I(N__9491));
    Odrv4 I__2159 (
            .O(N__9491),
            .I(N_185_i));
    InMux I__2158 (
            .O(N__9488),
            .I(N__9485));
    LocalMux I__2157 (
            .O(N__9485),
            .I(READ_CYCLE_ACTIVE_rep2_i_ess));
    IoInMux I__2156 (
            .O(N__9482),
            .I(N__9479));
    LocalMux I__2155 (
            .O(N__9479),
            .I(N__9476));
    Span4Mux_s2_v I__2154 (
            .O(N__9476),
            .I(N__9473));
    Span4Mux_v I__2153 (
            .O(N__9473),
            .I(N__9470));
    Odrv4 I__2152 (
            .O(N__9470),
            .I(N_183_i));
    InMux I__2151 (
            .O(N__9467),
            .I(N__9464));
    LocalMux I__2150 (
            .O(N__9464),
            .I(READ_CYCLE_ACTIVE_rep0_i_ess));
    IoInMux I__2149 (
            .O(N__9461),
            .I(N__9458));
    LocalMux I__2148 (
            .O(N__9458),
            .I(N__9455));
    Span4Mux_s0_v I__2147 (
            .O(N__9455),
            .I(N__9452));
    Span4Mux_v I__2146 (
            .O(N__9452),
            .I(N__9449));
    Span4Mux_v I__2145 (
            .O(N__9449),
            .I(N__9446));
    Odrv4 I__2144 (
            .O(N__9446),
            .I(N_181_i));
    InMux I__2143 (
            .O(N__9443),
            .I(N__9440));
    LocalMux I__2142 (
            .O(N__9440),
            .I(READ_CYCLE_ACTIVE_rep7_i_ess));
    IoInMux I__2141 (
            .O(N__9437),
            .I(N__9434));
    LocalMux I__2140 (
            .O(N__9434),
            .I(N__9431));
    Span4Mux_s2_v I__2139 (
            .O(N__9431),
            .I(N__9428));
    Span4Mux_v I__2138 (
            .O(N__9428),
            .I(N__9425));
    Odrv4 I__2137 (
            .O(N__9425),
            .I(N_188_i));
    IoInMux I__2136 (
            .O(N__9422),
            .I(N__9419));
    LocalMux I__2135 (
            .O(N__9419),
            .I(N__9416));
    IoSpan4Mux I__2134 (
            .O(N__9416),
            .I(N__9413));
    IoSpan4Mux I__2133 (
            .O(N__9413),
            .I(N__9410));
    Span4Mux_s2_h I__2132 (
            .O(N__9410),
            .I(N__9407));
    Odrv4 I__2131 (
            .O(N__9407),
            .I(N_209_i));
    InMux I__2130 (
            .O(N__9404),
            .I(N__9401));
    LocalMux I__2129 (
            .O(N__9401),
            .I(READ_CYCLE_ACTIVE_rep28_i_ess));
    InMux I__2128 (
            .O(N__9398),
            .I(N__9395));
    LocalMux I__2127 (
            .O(N__9395),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ));
    InMux I__2126 (
            .O(N__9392),
            .I(N__9388));
    InMux I__2125 (
            .O(N__9391),
            .I(N__9385));
    LocalMux I__2124 (
            .O(N__9388),
            .I(N__9381));
    LocalMux I__2123 (
            .O(N__9385),
            .I(N__9378));
    InMux I__2122 (
            .O(N__9384),
            .I(N__9375));
    Span4Mux_v I__2121 (
            .O(N__9381),
            .I(N__9372));
    Span4Mux_h I__2120 (
            .O(N__9378),
            .I(N__9367));
    LocalMux I__2119 (
            .O(N__9375),
            .I(N__9367));
    Span4Mux_v I__2118 (
            .O(N__9372),
            .I(N__9362));
    Span4Mux_h I__2117 (
            .O(N__9367),
            .I(N__9362));
    Span4Mux_v I__2116 (
            .O(N__9362),
            .I(N__9359));
    Sp12to4 I__2115 (
            .O(N__9359),
            .I(N__9356));
    Span12Mux_h I__2114 (
            .O(N__9356),
            .I(N__9353));
    Odrv12 I__2113 (
            .O(N__9353),
            .I(D_UM_AMIGA_in_2));
    IoInMux I__2112 (
            .O(N__9350),
            .I(N__9347));
    LocalMux I__2111 (
            .O(N__9347),
            .I(N__9344));
    Span12Mux_s6_h I__2110 (
            .O(N__9344),
            .I(N__9341));
    Odrv12 I__2109 (
            .O(N__9341),
            .I(un1_D_UM_AMIGA_2));
    InMux I__2108 (
            .O(N__9338),
            .I(N__9335));
    LocalMux I__2107 (
            .O(N__9335),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ));
    InMux I__2106 (
            .O(N__9332),
            .I(N__9329));
    LocalMux I__2105 (
            .O(N__9329),
            .I(N__9325));
    InMux I__2104 (
            .O(N__9328),
            .I(N__9322));
    Span4Mux_v I__2103 (
            .O(N__9325),
            .I(N__9318));
    LocalMux I__2102 (
            .O(N__9322),
            .I(N__9315));
    InMux I__2101 (
            .O(N__9321),
            .I(N__9312));
    Span4Mux_v I__2100 (
            .O(N__9318),
            .I(N__9309));
    Span4Mux_v I__2099 (
            .O(N__9315),
            .I(N__9306));
    LocalMux I__2098 (
            .O(N__9312),
            .I(N__9303));
    Sp12to4 I__2097 (
            .O(N__9309),
            .I(N__9296));
    Sp12to4 I__2096 (
            .O(N__9306),
            .I(N__9296));
    Span12Mux_v I__2095 (
            .O(N__9303),
            .I(N__9296));
    Span12Mux_h I__2094 (
            .O(N__9296),
            .I(N__9293));
    Span12Mux_v I__2093 (
            .O(N__9293),
            .I(N__9290));
    Odrv12 I__2092 (
            .O(N__9290),
            .I(D_UM_AMIGA_in_6));
    IoInMux I__2091 (
            .O(N__9287),
            .I(N__9284));
    LocalMux I__2090 (
            .O(N__9284),
            .I(N__9281));
    IoSpan4Mux I__2089 (
            .O(N__9281),
            .I(N__9278));
    Span4Mux_s2_h I__2088 (
            .O(N__9278),
            .I(N__9275));
    Sp12to4 I__2087 (
            .O(N__9275),
            .I(N__9272));
    Odrv12 I__2086 (
            .O(N__9272),
            .I(un1_D_UM_AMIGA_6));
    IoInMux I__2085 (
            .O(N__9269),
            .I(N__9265));
    InMux I__2084 (
            .O(N__9268),
            .I(N__9262));
    LocalMux I__2083 (
            .O(N__9265),
            .I(N__9259));
    LocalMux I__2082 (
            .O(N__9262),
            .I(N__9256));
    Span4Mux_s2_h I__2081 (
            .O(N__9259),
            .I(N__9253));
    Sp12to4 I__2080 (
            .O(N__9256),
            .I(N__9250));
    Span4Mux_v I__2079 (
            .O(N__9253),
            .I(N__9247));
    Span12Mux_v I__2078 (
            .O(N__9250),
            .I(N__9244));
    Sp12to4 I__2077 (
            .O(N__9247),
            .I(N__9241));
    Span12Mux_v I__2076 (
            .O(N__9244),
            .I(N__9238));
    Span12Mux_h I__2075 (
            .O(N__9241),
            .I(N__9235));
    Span12Mux_h I__2074 (
            .O(N__9238),
            .I(N__9232));
    Span12Mux_h I__2073 (
            .O(N__9235),
            .I(N__9229));
    Odrv12 I__2072 (
            .O(N__9232),
            .I(D_LL_040_in_4));
    Odrv12 I__2071 (
            .O(N__9229),
            .I(D_LL_040_in_4));
    InMux I__2070 (
            .O(N__9224),
            .I(N__9221));
    LocalMux I__2069 (
            .O(N__9221),
            .I(N__9218));
    Span4Mux_v I__2068 (
            .O(N__9218),
            .I(N__9215));
    Sp12to4 I__2067 (
            .O(N__9215),
            .I(N__9212));
    Span12Mux_h I__2066 (
            .O(N__9212),
            .I(N__9209));
    Odrv12 I__2065 (
            .O(N__9209),
            .I(D_UM_040_in_4));
    IoInMux I__2064 (
            .O(N__9206),
            .I(N__9203));
    LocalMux I__2063 (
            .O(N__9203),
            .I(N__9200));
    IoSpan4Mux I__2062 (
            .O(N__9200),
            .I(N__9197));
    Span4Mux_s3_h I__2061 (
            .O(N__9197),
            .I(N__9194));
    Span4Mux_h I__2060 (
            .O(N__9194),
            .I(N__9191));
    Span4Mux_h I__2059 (
            .O(N__9191),
            .I(N__9188));
    Span4Mux_h I__2058 (
            .O(N__9188),
            .I(N__9185));
    Odrv4 I__2057 (
            .O(N__9185),
            .I(un1_D_UM_040_4));
    InMux I__2056 (
            .O(N__9182),
            .I(N__9179));
    LocalMux I__2055 (
            .O(N__9179),
            .I(N__9176));
    Span4Mux_v I__2054 (
            .O(N__9176),
            .I(N__9173));
    Span4Mux_h I__2053 (
            .O(N__9173),
            .I(N__9170));
    Span4Mux_h I__2052 (
            .O(N__9170),
            .I(N__9167));
    Odrv4 I__2051 (
            .O(N__9167),
            .I(D_UU_040_in_4));
    IoInMux I__2050 (
            .O(N__9164),
            .I(N__9161));
    LocalMux I__2049 (
            .O(N__9161),
            .I(N__9158));
    Span4Mux_s1_h I__2048 (
            .O(N__9158),
            .I(N__9155));
    Sp12to4 I__2047 (
            .O(N__9155),
            .I(N__9151));
    InMux I__2046 (
            .O(N__9154),
            .I(N__9148));
    Span12Mux_v I__2045 (
            .O(N__9151),
            .I(N__9145));
    LocalMux I__2044 (
            .O(N__9148),
            .I(N__9142));
    Span12Mux_h I__2043 (
            .O(N__9145),
            .I(N__9139));
    Span12Mux_h I__2042 (
            .O(N__9142),
            .I(N__9136));
    Span12Mux_h I__2041 (
            .O(N__9139),
            .I(N__9131));
    Span12Mux_v I__2040 (
            .O(N__9136),
            .I(N__9131));
    Odrv12 I__2039 (
            .O(N__9131),
            .I(D_LM_040_in_4));
    IoInMux I__2038 (
            .O(N__9128),
            .I(N__9125));
    LocalMux I__2037 (
            .O(N__9125),
            .I(N__9122));
    IoSpan4Mux I__2036 (
            .O(N__9122),
            .I(N__9119));
    Sp12to4 I__2035 (
            .O(N__9119),
            .I(N__9116));
    Span12Mux_s6_v I__2034 (
            .O(N__9116),
            .I(N__9113));
    Odrv12 I__2033 (
            .O(N__9113),
            .I(un1_D_UU_040_4));
    InMux I__2032 (
            .O(N__9110),
            .I(N__9097));
    InMux I__2031 (
            .O(N__9109),
            .I(N__9097));
    InMux I__2030 (
            .O(N__9108),
            .I(N__9097));
    InMux I__2029 (
            .O(N__9107),
            .I(N__9092));
    CascadeMux I__2028 (
            .O(N__9106),
            .I(N__9086));
    InMux I__2027 (
            .O(N__9105),
            .I(N__9080));
    InMux I__2026 (
            .O(N__9104),
            .I(N__9080));
    LocalMux I__2025 (
            .O(N__9097),
            .I(N__9077));
    InMux I__2024 (
            .O(N__9096),
            .I(N__9074));
    InMux I__2023 (
            .O(N__9095),
            .I(N__9071));
    LocalMux I__2022 (
            .O(N__9092),
            .I(N__9068));
    InMux I__2021 (
            .O(N__9091),
            .I(N__9063));
    InMux I__2020 (
            .O(N__9090),
            .I(N__9063));
    InMux I__2019 (
            .O(N__9089),
            .I(N__9056));
    InMux I__2018 (
            .O(N__9086),
            .I(N__9056));
    InMux I__2017 (
            .O(N__9085),
            .I(N__9056));
    LocalMux I__2016 (
            .O(N__9080),
            .I(N__9053));
    Span4Mux_h I__2015 (
            .O(N__9077),
            .I(N__9046));
    LocalMux I__2014 (
            .O(N__9074),
            .I(N__9046));
    LocalMux I__2013 (
            .O(N__9071),
            .I(N__9043));
    Span4Mux_h I__2012 (
            .O(N__9068),
            .I(N__9038));
    LocalMux I__2011 (
            .O(N__9063),
            .I(N__9038));
    LocalMux I__2010 (
            .O(N__9056),
            .I(N__9033));
    Span4Mux_h I__2009 (
            .O(N__9053),
            .I(N__9033));
    InMux I__2008 (
            .O(N__9052),
            .I(N__9030));
    InMux I__2007 (
            .O(N__9051),
            .I(N__9027));
    Span4Mux_v I__2006 (
            .O(N__9046),
            .I(N__9022));
    Sp12to4 I__2005 (
            .O(N__9043),
            .I(N__9011));
    Sp12to4 I__2004 (
            .O(N__9038),
            .I(N__9011));
    Sp12to4 I__2003 (
            .O(N__9033),
            .I(N__9011));
    LocalMux I__2002 (
            .O(N__9030),
            .I(N__9011));
    LocalMux I__2001 (
            .O(N__9027),
            .I(N__9011));
    InMux I__2000 (
            .O(N__9026),
            .I(N__9008));
    CascadeMux I__1999 (
            .O(N__9025),
            .I(N__9005));
    Span4Mux_v I__1998 (
            .O(N__9022),
            .I(N__9002));
    Span12Mux_v I__1997 (
            .O(N__9011),
            .I(N__8999));
    LocalMux I__1996 (
            .O(N__9008),
            .I(N__8996));
    InMux I__1995 (
            .O(N__9005),
            .I(N__8993));
    Odrv4 I__1994 (
            .O(N__9002),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    Odrv12 I__1993 (
            .O(N__8999),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    Odrv12 I__1992 (
            .O(N__8996),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    LocalMux I__1991 (
            .O(N__8993),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    InMux I__1990 (
            .O(N__8984),
            .I(N__8981));
    LocalMux I__1989 (
            .O(N__8981),
            .I(N__8978));
    Odrv4 I__1988 (
            .O(N__8978),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ));
    InMux I__1987 (
            .O(N__8975),
            .I(N__8972));
    LocalMux I__1986 (
            .O(N__8972),
            .I(N__8968));
    InMux I__1985 (
            .O(N__8971),
            .I(N__8964));
    Span4Mux_v I__1984 (
            .O(N__8968),
            .I(N__8961));
    InMux I__1983 (
            .O(N__8967),
            .I(N__8958));
    LocalMux I__1982 (
            .O(N__8964),
            .I(N__8955));
    Span4Mux_v I__1981 (
            .O(N__8961),
            .I(N__8952));
    LocalMux I__1980 (
            .O(N__8958),
            .I(N__8949));
    Span4Mux_v I__1979 (
            .O(N__8955),
            .I(N__8946));
    Span4Mux_v I__1978 (
            .O(N__8952),
            .I(N__8943));
    Span4Mux_v I__1977 (
            .O(N__8949),
            .I(N__8940));
    Sp12to4 I__1976 (
            .O(N__8946),
            .I(N__8933));
    Sp12to4 I__1975 (
            .O(N__8943),
            .I(N__8933));
    Sp12to4 I__1974 (
            .O(N__8940),
            .I(N__8933));
    Span12Mux_h I__1973 (
            .O(N__8933),
            .I(N__8930));
    Odrv12 I__1972 (
            .O(N__8930),
            .I(D_UM_AMIGA_in_0));
    IoInMux I__1971 (
            .O(N__8927),
            .I(N__8924));
    LocalMux I__1970 (
            .O(N__8924),
            .I(N__8921));
    Span12Mux_s8_h I__1969 (
            .O(N__8921),
            .I(N__8918));
    Odrv12 I__1968 (
            .O(N__8918),
            .I(un1_D_UM_AMIGA_0));
    InMux I__1967 (
            .O(N__8915),
            .I(N__8912));
    LocalMux I__1966 (
            .O(N__8912),
            .I(N__8909));
    Span4Mux_v I__1965 (
            .O(N__8909),
            .I(N__8906));
    Span4Mux_v I__1964 (
            .O(N__8906),
            .I(N__8903));
    Sp12to4 I__1963 (
            .O(N__8903),
            .I(N__8900));
    Span12Mux_h I__1962 (
            .O(N__8900),
            .I(N__8897));
    Odrv12 I__1961 (
            .O(N__8897),
            .I(D_UM_040_in_7));
    IoInMux I__1960 (
            .O(N__8894),
            .I(N__8891));
    LocalMux I__1959 (
            .O(N__8891),
            .I(N__8887));
    InMux I__1958 (
            .O(N__8890),
            .I(N__8884));
    IoSpan4Mux I__1957 (
            .O(N__8887),
            .I(N__8881));
    LocalMux I__1956 (
            .O(N__8884),
            .I(N__8878));
    Span4Mux_s3_h I__1955 (
            .O(N__8881),
            .I(N__8875));
    Span4Mux_h I__1954 (
            .O(N__8878),
            .I(N__8872));
    Sp12to4 I__1953 (
            .O(N__8875),
            .I(N__8869));
    Sp12to4 I__1952 (
            .O(N__8872),
            .I(N__8866));
    Span12Mux_v I__1951 (
            .O(N__8869),
            .I(N__8863));
    Span12Mux_v I__1950 (
            .O(N__8866),
            .I(N__8860));
    Span12Mux_h I__1949 (
            .O(N__8863),
            .I(N__8857));
    Span12Mux_v I__1948 (
            .O(N__8860),
            .I(N__8854));
    Span12Mux_h I__1947 (
            .O(N__8857),
            .I(N__8851));
    Span12Mux_h I__1946 (
            .O(N__8854),
            .I(N__8848));
    Odrv12 I__1945 (
            .O(N__8851),
            .I(D_LL_040_in_7));
    Odrv12 I__1944 (
            .O(N__8848),
            .I(D_LL_040_in_7));
    IoInMux I__1943 (
            .O(N__8843),
            .I(N__8840));
    LocalMux I__1942 (
            .O(N__8840),
            .I(N__8837));
    Span12Mux_s5_h I__1941 (
            .O(N__8837),
            .I(N__8834));
    Span12Mux_h I__1940 (
            .O(N__8834),
            .I(N__8831));
    Odrv12 I__1939 (
            .O(N__8831),
            .I(un1_D_UM_040_7));
    InMux I__1938 (
            .O(N__8828),
            .I(N__8824));
    InMux I__1937 (
            .O(N__8827),
            .I(N__8818));
    LocalMux I__1936 (
            .O(N__8824),
            .I(N__8812));
    InMux I__1935 (
            .O(N__8823),
            .I(N__8809));
    InMux I__1934 (
            .O(N__8822),
            .I(N__8804));
    InMux I__1933 (
            .O(N__8821),
            .I(N__8801));
    LocalMux I__1932 (
            .O(N__8818),
            .I(N__8793));
    InMux I__1931 (
            .O(N__8817),
            .I(N__8788));
    InMux I__1930 (
            .O(N__8816),
            .I(N__8785));
    InMux I__1929 (
            .O(N__8815),
            .I(N__8782));
    Span4Mux_h I__1928 (
            .O(N__8812),
            .I(N__8776));
    LocalMux I__1927 (
            .O(N__8809),
            .I(N__8776));
    InMux I__1926 (
            .O(N__8808),
            .I(N__8773));
    InMux I__1925 (
            .O(N__8807),
            .I(N__8770));
    LocalMux I__1924 (
            .O(N__8804),
            .I(N__8763));
    LocalMux I__1923 (
            .O(N__8801),
            .I(N__8763));
    InMux I__1922 (
            .O(N__8800),
            .I(N__8758));
    InMux I__1921 (
            .O(N__8799),
            .I(N__8758));
    InMux I__1920 (
            .O(N__8798),
            .I(N__8751));
    InMux I__1919 (
            .O(N__8797),
            .I(N__8751));
    InMux I__1918 (
            .O(N__8796),
            .I(N__8748));
    Span4Mux_v I__1917 (
            .O(N__8793),
            .I(N__8742));
    InMux I__1916 (
            .O(N__8792),
            .I(N__8736));
    InMux I__1915 (
            .O(N__8791),
            .I(N__8736));
    LocalMux I__1914 (
            .O(N__8788),
            .I(N__8731));
    LocalMux I__1913 (
            .O(N__8785),
            .I(N__8728));
    LocalMux I__1912 (
            .O(N__8782),
            .I(N__8725));
    InMux I__1911 (
            .O(N__8781),
            .I(N__8722));
    Span4Mux_h I__1910 (
            .O(N__8776),
            .I(N__8714));
    LocalMux I__1909 (
            .O(N__8773),
            .I(N__8714));
    LocalMux I__1908 (
            .O(N__8770),
            .I(N__8714));
    InMux I__1907 (
            .O(N__8769),
            .I(N__8711));
    InMux I__1906 (
            .O(N__8768),
            .I(N__8707));
    Span4Mux_h I__1905 (
            .O(N__8763),
            .I(N__8702));
    LocalMux I__1904 (
            .O(N__8758),
            .I(N__8702));
    InMux I__1903 (
            .O(N__8757),
            .I(N__8699));
    InMux I__1902 (
            .O(N__8756),
            .I(N__8696));
    LocalMux I__1901 (
            .O(N__8751),
            .I(N__8691));
    LocalMux I__1900 (
            .O(N__8748),
            .I(N__8691));
    InMux I__1899 (
            .O(N__8747),
            .I(N__8688));
    InMux I__1898 (
            .O(N__8746),
            .I(N__8685));
    InMux I__1897 (
            .O(N__8745),
            .I(N__8682));
    Span4Mux_v I__1896 (
            .O(N__8742),
            .I(N__8679));
    InMux I__1895 (
            .O(N__8741),
            .I(N__8676));
    LocalMux I__1894 (
            .O(N__8736),
            .I(N__8673));
    InMux I__1893 (
            .O(N__8735),
            .I(N__8670));
    InMux I__1892 (
            .O(N__8734),
            .I(N__8667));
    Span4Mux_h I__1891 (
            .O(N__8731),
            .I(N__8657));
    Span4Mux_h I__1890 (
            .O(N__8728),
            .I(N__8657));
    Span4Mux_v I__1889 (
            .O(N__8725),
            .I(N__8657));
    LocalMux I__1888 (
            .O(N__8722),
            .I(N__8657));
    InMux I__1887 (
            .O(N__8721),
            .I(N__8654));
    Span4Mux_v I__1886 (
            .O(N__8714),
            .I(N__8649));
    LocalMux I__1885 (
            .O(N__8711),
            .I(N__8649));
    InMux I__1884 (
            .O(N__8710),
            .I(N__8646));
    LocalMux I__1883 (
            .O(N__8707),
            .I(N__8642));
    Sp12to4 I__1882 (
            .O(N__8702),
            .I(N__8637));
    LocalMux I__1881 (
            .O(N__8699),
            .I(N__8637));
    LocalMux I__1880 (
            .O(N__8696),
            .I(N__8634));
    Span4Mux_v I__1879 (
            .O(N__8691),
            .I(N__8625));
    LocalMux I__1878 (
            .O(N__8688),
            .I(N__8625));
    LocalMux I__1877 (
            .O(N__8685),
            .I(N__8625));
    LocalMux I__1876 (
            .O(N__8682),
            .I(N__8625));
    Span4Mux_v I__1875 (
            .O(N__8679),
            .I(N__8616));
    LocalMux I__1874 (
            .O(N__8676),
            .I(N__8616));
    Span4Mux_v I__1873 (
            .O(N__8673),
            .I(N__8616));
    LocalMux I__1872 (
            .O(N__8670),
            .I(N__8616));
    LocalMux I__1871 (
            .O(N__8667),
            .I(N__8613));
    InMux I__1870 (
            .O(N__8666),
            .I(N__8610));
    Span4Mux_v I__1869 (
            .O(N__8657),
            .I(N__8605));
    LocalMux I__1868 (
            .O(N__8654),
            .I(N__8605));
    Span4Mux_h I__1867 (
            .O(N__8649),
            .I(N__8600));
    LocalMux I__1866 (
            .O(N__8646),
            .I(N__8600));
    InMux I__1865 (
            .O(N__8645),
            .I(N__8597));
    Span12Mux_v I__1864 (
            .O(N__8642),
            .I(N__8593));
    Span12Mux_v I__1863 (
            .O(N__8637),
            .I(N__8588));
    Span12Mux_v I__1862 (
            .O(N__8634),
            .I(N__8588));
    Span4Mux_v I__1861 (
            .O(N__8625),
            .I(N__8583));
    Span4Mux_h I__1860 (
            .O(N__8616),
            .I(N__8583));
    Span12Mux_s9_v I__1859 (
            .O(N__8613),
            .I(N__8578));
    LocalMux I__1858 (
            .O(N__8610),
            .I(N__8578));
    Span4Mux_v I__1857 (
            .O(N__8605),
            .I(N__8571));
    Span4Mux_v I__1856 (
            .O(N__8600),
            .I(N__8571));
    LocalMux I__1855 (
            .O(N__8597),
            .I(N__8571));
    InMux I__1854 (
            .O(N__8596),
            .I(N__8568));
    Odrv12 I__1853 (
            .O(N__8593),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv12 I__1852 (
            .O(N__8588),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv4 I__1851 (
            .O(N__8583),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv12 I__1850 (
            .O(N__8578),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv4 I__1849 (
            .O(N__8571),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    LocalMux I__1848 (
            .O(N__8568),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    InMux I__1847 (
            .O(N__8555),
            .I(N__8552));
    LocalMux I__1846 (
            .O(N__8552),
            .I(N__8549));
    Span4Mux_v I__1845 (
            .O(N__8549),
            .I(N__8546));
    Sp12to4 I__1844 (
            .O(N__8546),
            .I(N__8543));
    Span12Mux_h I__1843 (
            .O(N__8543),
            .I(N__8540));
    Odrv12 I__1842 (
            .O(N__8540),
            .I(D_UU_040_in_7));
    IoInMux I__1841 (
            .O(N__8537),
            .I(N__8534));
    LocalMux I__1840 (
            .O(N__8534),
            .I(N__8531));
    IoSpan4Mux I__1839 (
            .O(N__8531),
            .I(N__8528));
    Span4Mux_s2_h I__1838 (
            .O(N__8528),
            .I(N__8524));
    InMux I__1837 (
            .O(N__8527),
            .I(N__8521));
    Sp12to4 I__1836 (
            .O(N__8524),
            .I(N__8518));
    LocalMux I__1835 (
            .O(N__8521),
            .I(N__8515));
    Span12Mux_h I__1834 (
            .O(N__8518),
            .I(N__8512));
    Span12Mux_s9_v I__1833 (
            .O(N__8515),
            .I(N__8509));
    Span12Mux_h I__1832 (
            .O(N__8512),
            .I(N__8506));
    Span12Mux_h I__1831 (
            .O(N__8509),
            .I(N__8503));
    Odrv12 I__1830 (
            .O(N__8506),
            .I(D_LM_040_in_7));
    Odrv12 I__1829 (
            .O(N__8503),
            .I(D_LM_040_in_7));
    IoInMux I__1828 (
            .O(N__8498),
            .I(N__8495));
    LocalMux I__1827 (
            .O(N__8495),
            .I(N__8492));
    IoSpan4Mux I__1826 (
            .O(N__8492),
            .I(N__8489));
    Span4Mux_s3_v I__1825 (
            .O(N__8489),
            .I(N__8486));
    Span4Mux_h I__1824 (
            .O(N__8486),
            .I(N__8483));
    Span4Mux_h I__1823 (
            .O(N__8483),
            .I(N__8480));
    Span4Mux_h I__1822 (
            .O(N__8480),
            .I(N__8477));
    Odrv4 I__1821 (
            .O(N__8477),
            .I(un1_D_UU_040_7));
    InMux I__1820 (
            .O(N__8474),
            .I(N__8471));
    LocalMux I__1819 (
            .O(N__8471),
            .I(N__8468));
    Odrv12 I__1818 (
            .O(N__8468),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ));
    InMux I__1817 (
            .O(N__8465),
            .I(N__8461));
    InMux I__1816 (
            .O(N__8464),
            .I(N__8458));
    LocalMux I__1815 (
            .O(N__8461),
            .I(N__8454));
    LocalMux I__1814 (
            .O(N__8458),
            .I(N__8451));
    InMux I__1813 (
            .O(N__8457),
            .I(N__8448));
    Span4Mux_v I__1812 (
            .O(N__8454),
            .I(N__8445));
    Span4Mux_v I__1811 (
            .O(N__8451),
            .I(N__8440));
    LocalMux I__1810 (
            .O(N__8448),
            .I(N__8440));
    Span4Mux_v I__1809 (
            .O(N__8445),
            .I(N__8437));
    Span4Mux_v I__1808 (
            .O(N__8440),
            .I(N__8434));
    Sp12to4 I__1807 (
            .O(N__8437),
            .I(N__8431));
    Span4Mux_v I__1806 (
            .O(N__8434),
            .I(N__8428));
    Span12Mux_h I__1805 (
            .O(N__8431),
            .I(N__8425));
    Sp12to4 I__1804 (
            .O(N__8428),
            .I(N__8422));
    Span12Mux_v I__1803 (
            .O(N__8425),
            .I(N__8417));
    Span12Mux_h I__1802 (
            .O(N__8422),
            .I(N__8417));
    Odrv12 I__1801 (
            .O(N__8417),
            .I(D_UM_AMIGA_in_4));
    IoInMux I__1800 (
            .O(N__8414),
            .I(N__8411));
    LocalMux I__1799 (
            .O(N__8411),
            .I(N__8408));
    IoSpan4Mux I__1798 (
            .O(N__8408),
            .I(N__8405));
    Span4Mux_s2_v I__1797 (
            .O(N__8405),
            .I(N__8402));
    Sp12to4 I__1796 (
            .O(N__8402),
            .I(N__8399));
    Span12Mux_s10_v I__1795 (
            .O(N__8399),
            .I(N__8396));
    Odrv12 I__1794 (
            .O(N__8396),
            .I(un1_D_UM_AMIGA_4));
    InMux I__1793 (
            .O(N__8393),
            .I(N__8390));
    LocalMux I__1792 (
            .O(N__8390),
            .I(N__8387));
    Span4Mux_v I__1791 (
            .O(N__8387),
            .I(N__8384));
    Sp12to4 I__1790 (
            .O(N__8384),
            .I(N__8381));
    Span12Mux_h I__1789 (
            .O(N__8381),
            .I(N__8378));
    Odrv12 I__1788 (
            .O(N__8378),
            .I(D_LM_AMIGA_in_7));
    InMux I__1787 (
            .O(N__8375),
            .I(N__8372));
    LocalMux I__1786 (
            .O(N__8372),
            .I(N__8367));
    InMux I__1785 (
            .O(N__8371),
            .I(N__8364));
    InMux I__1784 (
            .O(N__8370),
            .I(N__8361));
    Sp12to4 I__1783 (
            .O(N__8367),
            .I(N__8358));
    LocalMux I__1782 (
            .O(N__8364),
            .I(N__8353));
    LocalMux I__1781 (
            .O(N__8361),
            .I(N__8353));
    Span12Mux_h I__1780 (
            .O(N__8358),
            .I(N__8350));
    Span12Mux_v I__1779 (
            .O(N__8353),
            .I(N__8347));
    Span12Mux_v I__1778 (
            .O(N__8350),
            .I(N__8342));
    Span12Mux_h I__1777 (
            .O(N__8347),
            .I(N__8342));
    Odrv12 I__1776 (
            .O(N__8342),
            .I(D_UU_AMIGA_in_7));
    IoInMux I__1775 (
            .O(N__8339),
            .I(N__8336));
    LocalMux I__1774 (
            .O(N__8336),
            .I(N__8333));
    Span12Mux_s7_h I__1773 (
            .O(N__8333),
            .I(N__8330));
    Odrv12 I__1772 (
            .O(N__8330),
            .I(un2_D_LM_AMIGA_7));
    InMux I__1771 (
            .O(N__8327),
            .I(N__8324));
    LocalMux I__1770 (
            .O(N__8324),
            .I(N__8321));
    Odrv12 I__1769 (
            .O(N__8321),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ));
    InMux I__1768 (
            .O(N__8318),
            .I(N__8315));
    LocalMux I__1767 (
            .O(N__8315),
            .I(N__8312));
    Span4Mux_v I__1766 (
            .O(N__8312),
            .I(N__8307));
    InMux I__1765 (
            .O(N__8311),
            .I(N__8304));
    InMux I__1764 (
            .O(N__8310),
            .I(N__8301));
    Sp12to4 I__1763 (
            .O(N__8307),
            .I(N__8296));
    LocalMux I__1762 (
            .O(N__8304),
            .I(N__8296));
    LocalMux I__1761 (
            .O(N__8301),
            .I(N__8293));
    Span12Mux_h I__1760 (
            .O(N__8296),
            .I(N__8290));
    Span12Mux_v I__1759 (
            .O(N__8293),
            .I(N__8287));
    Span12Mux_v I__1758 (
            .O(N__8290),
            .I(N__8284));
    Span12Mux_h I__1757 (
            .O(N__8287),
            .I(N__8281));
    Odrv12 I__1756 (
            .O(N__8284),
            .I(D_UM_AMIGA_in_7));
    Odrv12 I__1755 (
            .O(N__8281),
            .I(D_UM_AMIGA_in_7));
    IoInMux I__1754 (
            .O(N__8276),
            .I(N__8273));
    LocalMux I__1753 (
            .O(N__8273),
            .I(N__8270));
    Span12Mux_s4_h I__1752 (
            .O(N__8270),
            .I(N__8267));
    Span12Mux_h I__1751 (
            .O(N__8267),
            .I(N__8264));
    Odrv12 I__1750 (
            .O(N__8264),
            .I(un1_D_UM_AMIGA_7));
    InMux I__1749 (
            .O(N__8261),
            .I(N__8257));
    InMux I__1748 (
            .O(N__8260),
            .I(N__8253));
    LocalMux I__1747 (
            .O(N__8257),
            .I(N__8250));
    InMux I__1746 (
            .O(N__8256),
            .I(N__8247));
    LocalMux I__1745 (
            .O(N__8253),
            .I(N__8244));
    Sp12to4 I__1744 (
            .O(N__8250),
            .I(N__8241));
    LocalMux I__1743 (
            .O(N__8247),
            .I(N__8238));
    Span4Mux_v I__1742 (
            .O(N__8244),
            .I(N__8235));
    Span12Mux_v I__1741 (
            .O(N__8241),
            .I(N__8232));
    Span12Mux_h I__1740 (
            .O(N__8238),
            .I(N__8229));
    Sp12to4 I__1739 (
            .O(N__8235),
            .I(N__8226));
    Span12Mux_h I__1738 (
            .O(N__8232),
            .I(N__8223));
    Span12Mux_v I__1737 (
            .O(N__8229),
            .I(N__8218));
    Span12Mux_h I__1736 (
            .O(N__8226),
            .I(N__8218));
    Odrv12 I__1735 (
            .O(N__8223),
            .I(D_UM_AMIGA_in_5));
    Odrv12 I__1734 (
            .O(N__8218),
            .I(D_UM_AMIGA_in_5));
    InMux I__1733 (
            .O(N__8213),
            .I(N__8210));
    LocalMux I__1732 (
            .O(N__8210),
            .I(N__8207));
    Span12Mux_s8_v I__1731 (
            .O(N__8207),
            .I(N__8204));
    Odrv12 I__1730 (
            .O(N__8204),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ));
    IoInMux I__1729 (
            .O(N__8201),
            .I(N__8198));
    LocalMux I__1728 (
            .O(N__8198),
            .I(N__8195));
    IoSpan4Mux I__1727 (
            .O(N__8195),
            .I(N__8192));
    IoSpan4Mux I__1726 (
            .O(N__8192),
            .I(N__8189));
    IoSpan4Mux I__1725 (
            .O(N__8189),
            .I(N__8186));
    Span4Mux_s2_v I__1724 (
            .O(N__8186),
            .I(N__8183));
    Span4Mux_v I__1723 (
            .O(N__8183),
            .I(N__8180));
    Odrv4 I__1722 (
            .O(N__8180),
            .I(un1_D_UM_AMIGA_5));
    InMux I__1721 (
            .O(N__8177),
            .I(N__8174));
    LocalMux I__1720 (
            .O(N__8174),
            .I(N__8171));
    Span4Mux_v I__1719 (
            .O(N__8171),
            .I(N__8168));
    Sp12to4 I__1718 (
            .O(N__8168),
            .I(N__8165));
    Span12Mux_h I__1717 (
            .O(N__8165),
            .I(N__8162));
    Odrv12 I__1716 (
            .O(N__8162),
            .I(D_UU_040_in_2));
    InMux I__1715 (
            .O(N__8159),
            .I(N__8156));
    LocalMux I__1714 (
            .O(N__8156),
            .I(N__8152));
    IoInMux I__1713 (
            .O(N__8155),
            .I(N__8149));
    Span4Mux_h I__1712 (
            .O(N__8152),
            .I(N__8146));
    LocalMux I__1711 (
            .O(N__8149),
            .I(N__8143));
    Sp12to4 I__1710 (
            .O(N__8146),
            .I(N__8140));
    Span12Mux_s9_h I__1709 (
            .O(N__8143),
            .I(N__8137));
    Span12Mux_v I__1708 (
            .O(N__8140),
            .I(N__8134));
    Span12Mux_h I__1707 (
            .O(N__8137),
            .I(N__8131));
    Span12Mux_v I__1706 (
            .O(N__8134),
            .I(N__8128));
    Span12Mux_v I__1705 (
            .O(N__8131),
            .I(N__8125));
    Span12Mux_h I__1704 (
            .O(N__8128),
            .I(N__8122));
    Odrv12 I__1703 (
            .O(N__8125),
            .I(D_LM_040_in_2));
    Odrv12 I__1702 (
            .O(N__8122),
            .I(D_LM_040_in_2));
    IoInMux I__1701 (
            .O(N__8117),
            .I(N__8114));
    LocalMux I__1700 (
            .O(N__8114),
            .I(N__8111));
    IoSpan4Mux I__1699 (
            .O(N__8111),
            .I(N__8108));
    IoSpan4Mux I__1698 (
            .O(N__8108),
            .I(N__8105));
    Span4Mux_s3_v I__1697 (
            .O(N__8105),
            .I(N__8102));
    Span4Mux_h I__1696 (
            .O(N__8102),
            .I(N__8099));
    Odrv4 I__1695 (
            .O(N__8099),
            .I(un1_D_UU_040_2));
    InMux I__1694 (
            .O(N__8096),
            .I(N__8093));
    LocalMux I__1693 (
            .O(N__8093),
            .I(N__8090));
    Span4Mux_v I__1692 (
            .O(N__8090),
            .I(N__8087));
    Span4Mux_v I__1691 (
            .O(N__8087),
            .I(N__8084));
    Sp12to4 I__1690 (
            .O(N__8084),
            .I(N__8081));
    Span12Mux_h I__1689 (
            .O(N__8081),
            .I(N__8078));
    Odrv12 I__1688 (
            .O(N__8078),
            .I(D_UU_040_in_5));
    IoInMux I__1687 (
            .O(N__8075),
            .I(N__8072));
    LocalMux I__1686 (
            .O(N__8072),
            .I(N__8069));
    IoSpan4Mux I__1685 (
            .O(N__8069),
            .I(N__8065));
    InMux I__1684 (
            .O(N__8068),
            .I(N__8062));
    IoSpan4Mux I__1683 (
            .O(N__8065),
            .I(N__8059));
    LocalMux I__1682 (
            .O(N__8062),
            .I(N__8056));
    Span4Mux_s2_h I__1681 (
            .O(N__8059),
            .I(N__8053));
    Span4Mux_v I__1680 (
            .O(N__8056),
            .I(N__8050));
    Sp12to4 I__1679 (
            .O(N__8053),
            .I(N__8047));
    Sp12to4 I__1678 (
            .O(N__8050),
            .I(N__8044));
    Span12Mux_h I__1677 (
            .O(N__8047),
            .I(N__8041));
    Span12Mux_h I__1676 (
            .O(N__8044),
            .I(N__8038));
    Span12Mux_h I__1675 (
            .O(N__8041),
            .I(N__8035));
    Span12Mux_v I__1674 (
            .O(N__8038),
            .I(N__8032));
    Odrv12 I__1673 (
            .O(N__8035),
            .I(D_LM_040_in_5));
    Odrv12 I__1672 (
            .O(N__8032),
            .I(D_LM_040_in_5));
    IoInMux I__1671 (
            .O(N__8027),
            .I(N__8024));
    LocalMux I__1670 (
            .O(N__8024),
            .I(N__8021));
    Span4Mux_s3_h I__1669 (
            .O(N__8021),
            .I(N__8018));
    Sp12to4 I__1668 (
            .O(N__8018),
            .I(N__8015));
    Span12Mux_s7_v I__1667 (
            .O(N__8015),
            .I(N__8012));
    Span12Mux_h I__1666 (
            .O(N__8012),
            .I(N__8009));
    Odrv12 I__1665 (
            .O(N__8009),
            .I(un1_D_UU_040_5));
    InMux I__1664 (
            .O(N__8006),
            .I(N__8002));
    InMux I__1663 (
            .O(N__8005),
            .I(N__7999));
    LocalMux I__1662 (
            .O(N__8002),
            .I(N__7996));
    LocalMux I__1661 (
            .O(N__7999),
            .I(N__7993));
    Span4Mux_v I__1660 (
            .O(N__7996),
            .I(N__7989));
    Span4Mux_v I__1659 (
            .O(N__7993),
            .I(N__7986));
    InMux I__1658 (
            .O(N__7992),
            .I(N__7983));
    Span4Mux_v I__1657 (
            .O(N__7989),
            .I(N__7980));
    Span4Mux_v I__1656 (
            .O(N__7986),
            .I(N__7975));
    LocalMux I__1655 (
            .O(N__7983),
            .I(N__7975));
    Span4Mux_v I__1654 (
            .O(N__7980),
            .I(N__7970));
    Span4Mux_v I__1653 (
            .O(N__7975),
            .I(N__7970));
    Sp12to4 I__1652 (
            .O(N__7970),
            .I(N__7967));
    Span12Mux_h I__1651 (
            .O(N__7967),
            .I(N__7964));
    Odrv12 I__1650 (
            .O(N__7964),
            .I(D_UU_AMIGA_in_3));
    InMux I__1649 (
            .O(N__7961),
            .I(N__7958));
    LocalMux I__1648 (
            .O(N__7958),
            .I(N__7955));
    Span12Mux_s7_v I__1647 (
            .O(N__7955),
            .I(N__7952));
    Odrv12 I__1646 (
            .O(N__7952),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ));
    IoInMux I__1645 (
            .O(N__7949),
            .I(N__7946));
    LocalMux I__1644 (
            .O(N__7946),
            .I(N__7943));
    Span4Mux_s2_v I__1643 (
            .O(N__7943),
            .I(N__7940));
    Span4Mux_h I__1642 (
            .O(N__7940),
            .I(N__7937));
    Span4Mux_v I__1641 (
            .O(N__7937),
            .I(N__7934));
    Sp12to4 I__1640 (
            .O(N__7934),
            .I(N__7931));
    Odrv12 I__1639 (
            .O(N__7931),
            .I(un1_D_UU_AMIGA_3));
    InMux I__1638 (
            .O(N__7928),
            .I(N__7924));
    InMux I__1637 (
            .O(N__7927),
            .I(N__7921));
    LocalMux I__1636 (
            .O(N__7924),
            .I(N__7917));
    LocalMux I__1635 (
            .O(N__7921),
            .I(N__7914));
    InMux I__1634 (
            .O(N__7920),
            .I(N__7911));
    Span12Mux_v I__1633 (
            .O(N__7917),
            .I(N__7904));
    Span12Mux_s9_v I__1632 (
            .O(N__7914),
            .I(N__7904));
    LocalMux I__1631 (
            .O(N__7911),
            .I(N__7904));
    Span12Mux_h I__1630 (
            .O(N__7904),
            .I(N__7901));
    Odrv12 I__1629 (
            .O(N__7901),
            .I(D_UU_AMIGA_in_6));
    InMux I__1628 (
            .O(N__7898),
            .I(N__7895));
    LocalMux I__1627 (
            .O(N__7895),
            .I(N__7892));
    Span12Mux_s11_v I__1626 (
            .O(N__7892),
            .I(N__7889));
    Odrv12 I__1625 (
            .O(N__7889),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ));
    IoInMux I__1624 (
            .O(N__7886),
            .I(N__7883));
    LocalMux I__1623 (
            .O(N__7883),
            .I(N__7880));
    Span4Mux_s0_v I__1622 (
            .O(N__7880),
            .I(N__7877));
    Sp12to4 I__1621 (
            .O(N__7877),
            .I(N__7874));
    Span12Mux_h I__1620 (
            .O(N__7874),
            .I(N__7871));
    Odrv12 I__1619 (
            .O(N__7871),
            .I(un1_D_UU_AMIGA_6));
    CEMux I__1618 (
            .O(N__7868),
            .I(N__7862));
    CEMux I__1617 (
            .O(N__7867),
            .I(N__7859));
    CEMux I__1616 (
            .O(N__7866),
            .I(N__7854));
    CEMux I__1615 (
            .O(N__7865),
            .I(N__7851));
    LocalMux I__1614 (
            .O(N__7862),
            .I(N__7848));
    LocalMux I__1613 (
            .O(N__7859),
            .I(N__7845));
    CEMux I__1612 (
            .O(N__7858),
            .I(N__7842));
    CEMux I__1611 (
            .O(N__7857),
            .I(N__7839));
    LocalMux I__1610 (
            .O(N__7854),
            .I(N__7836));
    LocalMux I__1609 (
            .O(N__7851),
            .I(N__7833));
    Span4Mux_v I__1608 (
            .O(N__7848),
            .I(N__7826));
    Span4Mux_h I__1607 (
            .O(N__7845),
            .I(N__7826));
    LocalMux I__1606 (
            .O(N__7842),
            .I(N__7826));
    LocalMux I__1605 (
            .O(N__7839),
            .I(N__7823));
    Span4Mux_v I__1604 (
            .O(N__7836),
            .I(N__7820));
    Span4Mux_h I__1603 (
            .O(N__7833),
            .I(N__7817));
    Span4Mux_v I__1602 (
            .O(N__7826),
            .I(N__7814));
    Odrv4 I__1601 (
            .O(N__7823),
            .I(\U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0 ));
    Odrv4 I__1600 (
            .O(N__7820),
            .I(\U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0 ));
    Odrv4 I__1599 (
            .O(N__7817),
            .I(\U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0 ));
    Odrv4 I__1598 (
            .O(N__7814),
            .I(\U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0 ));
    SRMux I__1597 (
            .O(N__7805),
            .I(N__7802));
    LocalMux I__1596 (
            .O(N__7802),
            .I(N__7799));
    Span4Mux_h I__1595 (
            .O(N__7799),
            .I(N__7791));
    SRMux I__1594 (
            .O(N__7798),
            .I(N__7788));
    SRMux I__1593 (
            .O(N__7797),
            .I(N__7785));
    SRMux I__1592 (
            .O(N__7796),
            .I(N__7782));
    SRMux I__1591 (
            .O(N__7795),
            .I(N__7779));
    SRMux I__1590 (
            .O(N__7794),
            .I(N__7776));
    Odrv4 I__1589 (
            .O(N__7791),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1 ));
    LocalMux I__1588 (
            .O(N__7788),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1 ));
    LocalMux I__1587 (
            .O(N__7785),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1 ));
    LocalMux I__1586 (
            .O(N__7782),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1 ));
    LocalMux I__1585 (
            .O(N__7779),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1 ));
    LocalMux I__1584 (
            .O(N__7776),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1 ));
    InMux I__1583 (
            .O(N__7763),
            .I(N__7760));
    LocalMux I__1582 (
            .O(N__7760),
            .I(N__7757));
    Glb2LocalMux I__1581 (
            .O(N__7757),
            .I(N__7754));
    GlobalMux I__1580 (
            .O(N__7754),
            .I(CLK80));
    IoInMux I__1579 (
            .O(N__7751),
            .I(N__7747));
    IoInMux I__1578 (
            .O(N__7750),
            .I(N__7744));
    LocalMux I__1577 (
            .O(N__7747),
            .I(N__7741));
    LocalMux I__1576 (
            .O(N__7744),
            .I(N__7738));
    Span4Mux_s3_v I__1575 (
            .O(N__7741),
            .I(N__7735));
    IoSpan4Mux I__1574 (
            .O(N__7738),
            .I(N__7732));
    Span4Mux_v I__1573 (
            .O(N__7735),
            .I(N__7729));
    Span4Mux_s3_h I__1572 (
            .O(N__7732),
            .I(N__7726));
    Span4Mux_v I__1571 (
            .O(N__7729),
            .I(N__7723));
    Span4Mux_h I__1570 (
            .O(N__7726),
            .I(N__7720));
    Span4Mux_v I__1569 (
            .O(N__7723),
            .I(N__7717));
    Sp12to4 I__1568 (
            .O(N__7720),
            .I(N__7714));
    Odrv4 I__1567 (
            .O(N__7717),
            .I(GB_BUFFER_CLK80_THRU_CO));
    Odrv12 I__1566 (
            .O(N__7714),
            .I(GB_BUFFER_CLK80_THRU_CO));
    InMux I__1565 (
            .O(N__7709),
            .I(N__7706));
    LocalMux I__1564 (
            .O(N__7706),
            .I(N__7703));
    Odrv4 I__1563 (
            .O(N__7703),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ));
    InMux I__1562 (
            .O(N__7700),
            .I(N__7695));
    InMux I__1561 (
            .O(N__7699),
            .I(N__7692));
    InMux I__1560 (
            .O(N__7698),
            .I(N__7689));
    LocalMux I__1559 (
            .O(N__7695),
            .I(N__7684));
    LocalMux I__1558 (
            .O(N__7692),
            .I(N__7684));
    LocalMux I__1557 (
            .O(N__7689),
            .I(N__7681));
    Span4Mux_v I__1556 (
            .O(N__7684),
            .I(N__7678));
    Span4Mux_v I__1555 (
            .O(N__7681),
            .I(N__7675));
    Sp12to4 I__1554 (
            .O(N__7678),
            .I(N__7672));
    Span4Mux_h I__1553 (
            .O(N__7675),
            .I(N__7669));
    Span12Mux_h I__1552 (
            .O(N__7672),
            .I(N__7664));
    Sp12to4 I__1551 (
            .O(N__7669),
            .I(N__7664));
    Odrv12 I__1550 (
            .O(N__7664),
            .I(D_UU_AMIGA_in_2));
    IoInMux I__1549 (
            .O(N__7661),
            .I(N__7658));
    LocalMux I__1548 (
            .O(N__7658),
            .I(N__7655));
    IoSpan4Mux I__1547 (
            .O(N__7655),
            .I(N__7652));
    Span4Mux_s0_v I__1546 (
            .O(N__7652),
            .I(N__7649));
    Sp12to4 I__1545 (
            .O(N__7649),
            .I(N__7646));
    Span12Mux_v I__1544 (
            .O(N__7646),
            .I(N__7643));
    Odrv12 I__1543 (
            .O(N__7643),
            .I(un1_D_UU_AMIGA_2));
    InMux I__1542 (
            .O(N__7640),
            .I(N__7637));
    LocalMux I__1541 (
            .O(N__7637),
            .I(N__7634));
    Odrv12 I__1540 (
            .O(N__7634),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ));
    IoInMux I__1539 (
            .O(N__7631),
            .I(N__7628));
    LocalMux I__1538 (
            .O(N__7628),
            .I(N__7625));
    Span4Mux_s0_v I__1537 (
            .O(N__7625),
            .I(N__7622));
    Sp12to4 I__1536 (
            .O(N__7622),
            .I(N__7619));
    Span12Mux_s9_h I__1535 (
            .O(N__7619),
            .I(N__7616));
    Span12Mux_v I__1534 (
            .O(N__7616),
            .I(N__7613));
    Odrv12 I__1533 (
            .O(N__7613),
            .I(un1_D_UU_AMIGA_7));
    InMux I__1532 (
            .O(N__7610),
            .I(N__7607));
    LocalMux I__1531 (
            .O(N__7607),
            .I(N__7604));
    Odrv4 I__1530 (
            .O(N__7604),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ));
    InMux I__1529 (
            .O(N__7601),
            .I(N__7596));
    InMux I__1528 (
            .O(N__7600),
            .I(N__7593));
    InMux I__1527 (
            .O(N__7599),
            .I(N__7590));
    LocalMux I__1526 (
            .O(N__7596),
            .I(N__7585));
    LocalMux I__1525 (
            .O(N__7593),
            .I(N__7585));
    LocalMux I__1524 (
            .O(N__7590),
            .I(N__7582));
    Span4Mux_v I__1523 (
            .O(N__7585),
            .I(N__7579));
    Span12Mux_h I__1522 (
            .O(N__7582),
            .I(N__7576));
    Sp12to4 I__1521 (
            .O(N__7579),
            .I(N__7573));
    Span12Mux_v I__1520 (
            .O(N__7576),
            .I(N__7570));
    Span12Mux_h I__1519 (
            .O(N__7573),
            .I(N__7567));
    Odrv12 I__1518 (
            .O(N__7570),
            .I(D_UU_AMIGA_in_4));
    Odrv12 I__1517 (
            .O(N__7567),
            .I(D_UU_AMIGA_in_4));
    IoInMux I__1516 (
            .O(N__7562),
            .I(N__7559));
    LocalMux I__1515 (
            .O(N__7559),
            .I(N__7556));
    IoSpan4Mux I__1514 (
            .O(N__7556),
            .I(N__7553));
    Span4Mux_s2_v I__1513 (
            .O(N__7553),
            .I(N__7550));
    Sp12to4 I__1512 (
            .O(N__7550),
            .I(N__7547));
    Span12Mux_h I__1511 (
            .O(N__7547),
            .I(N__7544));
    Odrv12 I__1510 (
            .O(N__7544),
            .I(un1_D_UU_AMIGA_4));
    InMux I__1509 (
            .O(N__7541),
            .I(N__7537));
    InMux I__1508 (
            .O(N__7540),
            .I(N__7533));
    LocalMux I__1507 (
            .O(N__7537),
            .I(N__7530));
    InMux I__1506 (
            .O(N__7536),
            .I(N__7527));
    LocalMux I__1505 (
            .O(N__7533),
            .I(N__7524));
    Span4Mux_v I__1504 (
            .O(N__7530),
            .I(N__7519));
    LocalMux I__1503 (
            .O(N__7527),
            .I(N__7519));
    Sp12to4 I__1502 (
            .O(N__7524),
            .I(N__7516));
    Span4Mux_v I__1501 (
            .O(N__7519),
            .I(N__7513));
    Span12Mux_v I__1500 (
            .O(N__7516),
            .I(N__7510));
    Span4Mux_v I__1499 (
            .O(N__7513),
            .I(N__7507));
    Span12Mux_v I__1498 (
            .O(N__7510),
            .I(N__7504));
    Sp12to4 I__1497 (
            .O(N__7507),
            .I(N__7501));
    Span12Mux_h I__1496 (
            .O(N__7504),
            .I(N__7498));
    Span12Mux_h I__1495 (
            .O(N__7501),
            .I(N__7495));
    Odrv12 I__1494 (
            .O(N__7498),
            .I(D_UM_AMIGA_in_3));
    Odrv12 I__1493 (
            .O(N__7495),
            .I(D_UM_AMIGA_in_3));
    InMux I__1492 (
            .O(N__7490),
            .I(N__7487));
    LocalMux I__1491 (
            .O(N__7487),
            .I(N__7484));
    Span4Mux_v I__1490 (
            .O(N__7484),
            .I(N__7481));
    Odrv4 I__1489 (
            .O(N__7481),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ));
    IoInMux I__1488 (
            .O(N__7478),
            .I(N__7475));
    LocalMux I__1487 (
            .O(N__7475),
            .I(N__7472));
    IoSpan4Mux I__1486 (
            .O(N__7472),
            .I(N__7469));
    Span4Mux_s2_h I__1485 (
            .O(N__7469),
            .I(N__7466));
    Sp12to4 I__1484 (
            .O(N__7466),
            .I(N__7463));
    Span12Mux_h I__1483 (
            .O(N__7463),
            .I(N__7460));
    Odrv12 I__1482 (
            .O(N__7460),
            .I(un1_D_UM_AMIGA_3));
    InMux I__1481 (
            .O(N__7457),
            .I(N__7454));
    LocalMux I__1480 (
            .O(N__7454),
            .I(N__7451));
    Span4Mux_v I__1479 (
            .O(N__7451),
            .I(N__7448));
    Sp12to4 I__1478 (
            .O(N__7448),
            .I(N__7445));
    Span12Mux_h I__1477 (
            .O(N__7445),
            .I(N__7442));
    Odrv12 I__1476 (
            .O(N__7442),
            .I(D_LL_AMIGA_in_5));
    IoInMux I__1475 (
            .O(N__7439),
            .I(N__7436));
    LocalMux I__1474 (
            .O(N__7436),
            .I(N__7433));
    IoSpan4Mux I__1473 (
            .O(N__7433),
            .I(N__7430));
    Span4Mux_s2_h I__1472 (
            .O(N__7430),
            .I(N__7427));
    Sp12to4 I__1471 (
            .O(N__7427),
            .I(N__7424));
    Span12Mux_h I__1470 (
            .O(N__7424),
            .I(N__7421));
    Odrv12 I__1469 (
            .O(N__7421),
            .I(un2_D_LL_AMIGA_5));
    IoInMux I__1468 (
            .O(N__7418),
            .I(N__7415));
    LocalMux I__1467 (
            .O(N__7415),
            .I(N__7411));
    CascadeMux I__1466 (
            .O(N__7414),
            .I(N__7406));
    Span4Mux_s1_v I__1465 (
            .O(N__7411),
            .I(N__7402));
    InMux I__1464 (
            .O(N__7410),
            .I(N__7399));
    InMux I__1463 (
            .O(N__7409),
            .I(N__7396));
    InMux I__1462 (
            .O(N__7406),
            .I(N__7391));
    InMux I__1461 (
            .O(N__7405),
            .I(N__7391));
    Span4Mux_v I__1460 (
            .O(N__7402),
            .I(N__7388));
    LocalMux I__1459 (
            .O(N__7399),
            .I(N__7383));
    LocalMux I__1458 (
            .O(N__7396),
            .I(N__7378));
    LocalMux I__1457 (
            .O(N__7391),
            .I(N__7378));
    Sp12to4 I__1456 (
            .O(N__7388),
            .I(N__7375));
    InMux I__1455 (
            .O(N__7387),
            .I(N__7372));
    InMux I__1454 (
            .O(N__7386),
            .I(N__7369));
    Span4Mux_v I__1453 (
            .O(N__7383),
            .I(N__7363));
    Span4Mux_v I__1452 (
            .O(N__7378),
            .I(N__7363));
    Span12Mux_h I__1451 (
            .O(N__7375),
            .I(N__7356));
    LocalMux I__1450 (
            .O(N__7372),
            .I(N__7356));
    LocalMux I__1449 (
            .O(N__7369),
            .I(N__7356));
    InMux I__1448 (
            .O(N__7368),
            .I(N__7353));
    Sp12to4 I__1447 (
            .O(N__7363),
            .I(N__7346));
    Span12Mux_v I__1446 (
            .O(N__7356),
            .I(N__7346));
    LocalMux I__1445 (
            .O(N__7353),
            .I(N__7346));
    Span12Mux_v I__1444 (
            .O(N__7346),
            .I(N__7343));
    Odrv12 I__1443 (
            .O(N__7343),
            .I(TACKn_in));
    IoInMux I__1442 (
            .O(N__7340),
            .I(N__7337));
    LocalMux I__1441 (
            .O(N__7337),
            .I(N__7334));
    Span4Mux_s1_v I__1440 (
            .O(N__7334),
            .I(N__7326));
    InMux I__1439 (
            .O(N__7333),
            .I(N__7323));
    InMux I__1438 (
            .O(N__7332),
            .I(N__7320));
    InMux I__1437 (
            .O(N__7331),
            .I(N__7317));
    InMux I__1436 (
            .O(N__7330),
            .I(N__7312));
    InMux I__1435 (
            .O(N__7329),
            .I(N__7312));
    Span4Mux_v I__1434 (
            .O(N__7326),
            .I(N__7308));
    LocalMux I__1433 (
            .O(N__7323),
            .I(N__7299));
    LocalMux I__1432 (
            .O(N__7320),
            .I(N__7299));
    LocalMux I__1431 (
            .O(N__7317),
            .I(N__7299));
    LocalMux I__1430 (
            .O(N__7312),
            .I(N__7299));
    InMux I__1429 (
            .O(N__7311),
            .I(N__7296));
    Span4Mux_v I__1428 (
            .O(N__7308),
            .I(N__7293));
    Span4Mux_v I__1427 (
            .O(N__7299),
            .I(N__7288));
    LocalMux I__1426 (
            .O(N__7296),
            .I(N__7288));
    Sp12to4 I__1425 (
            .O(N__7293),
            .I(N__7285));
    Span4Mux_v I__1424 (
            .O(N__7288),
            .I(N__7282));
    Span12Mux_h I__1423 (
            .O(N__7285),
            .I(N__7279));
    Span4Mux_h I__1422 (
            .O(N__7282),
            .I(N__7276));
    Span12Mux_v I__1421 (
            .O(N__7279),
            .I(N__7271));
    Sp12to4 I__1420 (
            .O(N__7276),
            .I(N__7271));
    Odrv12 I__1419 (
            .O(N__7271),
            .I(TEAn_c));
    InMux I__1418 (
            .O(N__7268),
            .I(N__7264));
    InMux I__1417 (
            .O(N__7267),
            .I(N__7261));
    LocalMux I__1416 (
            .O(N__7264),
            .I(N__7256));
    LocalMux I__1415 (
            .O(N__7261),
            .I(N__7256));
    Span4Mux_v I__1414 (
            .O(N__7256),
            .I(N__7250));
    InMux I__1413 (
            .O(N__7255),
            .I(N__7247));
    CascadeMux I__1412 (
            .O(N__7254),
            .I(N__7243));
    InMux I__1411 (
            .O(N__7253),
            .I(N__7237));
    Span4Mux_v I__1410 (
            .O(N__7250),
            .I(N__7232));
    LocalMux I__1409 (
            .O(N__7247),
            .I(N__7232));
    InMux I__1408 (
            .O(N__7246),
            .I(N__7227));
    InMux I__1407 (
            .O(N__7243),
            .I(N__7227));
    InMux I__1406 (
            .O(N__7242),
            .I(N__7224));
    InMux I__1405 (
            .O(N__7241),
            .I(N__7221));
    InMux I__1404 (
            .O(N__7240),
            .I(N__7218));
    LocalMux I__1403 (
            .O(N__7237),
            .I(N__7207));
    Sp12to4 I__1402 (
            .O(N__7232),
            .I(N__7207));
    LocalMux I__1401 (
            .O(N__7227),
            .I(N__7207));
    LocalMux I__1400 (
            .O(N__7224),
            .I(N__7207));
    LocalMux I__1399 (
            .O(N__7221),
            .I(N__7207));
    LocalMux I__1398 (
            .O(N__7218),
            .I(N__7204));
    Span12Mux_h I__1397 (
            .O(N__7207),
            .I(N__7201));
    Span12Mux_v I__1396 (
            .O(N__7204),
            .I(N__7198));
    Span12Mux_v I__1395 (
            .O(N__7201),
            .I(N__7195));
    Odrv12 I__1394 (
            .O(N__7198),
            .I(RESETn_c));
    Odrv12 I__1393 (
            .O(N__7195),
            .I(RESETn_c));
    InMux I__1392 (
            .O(N__7190),
            .I(N__7187));
    LocalMux I__1391 (
            .O(N__7187),
            .I(N__7183));
    CascadeMux I__1390 (
            .O(N__7186),
            .I(N__7180));
    Span4Mux_v I__1389 (
            .O(N__7183),
            .I(N__7177));
    InMux I__1388 (
            .O(N__7180),
            .I(N__7174));
    Odrv4 I__1387 (
            .O(N__7177),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ));
    LocalMux I__1386 (
            .O(N__7174),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ));
    CascadeMux I__1385 (
            .O(N__7169),
            .I(\U111_CYCLE_SM.CYCLE_STATE_srsts_i_o2_0_5_cascade_ ));
    InMux I__1384 (
            .O(N__7166),
            .I(N__7162));
    InMux I__1383 (
            .O(N__7165),
            .I(N__7158));
    LocalMux I__1382 (
            .O(N__7162),
            .I(N__7155));
    InMux I__1381 (
            .O(N__7161),
            .I(N__7151));
    LocalMux I__1380 (
            .O(N__7158),
            .I(N__7145));
    Span4Mux_v I__1379 (
            .O(N__7155),
            .I(N__7145));
    InMux I__1378 (
            .O(N__7154),
            .I(N__7142));
    LocalMux I__1377 (
            .O(N__7151),
            .I(N__7139));
    InMux I__1376 (
            .O(N__7150),
            .I(N__7136));
    Odrv4 I__1375 (
            .O(N__7145),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    LocalMux I__1374 (
            .O(N__7142),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    Odrv4 I__1373 (
            .O(N__7139),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    LocalMux I__1372 (
            .O(N__7136),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    InMux I__1371 (
            .O(N__7127),
            .I(N__7124));
    LocalMux I__1370 (
            .O(N__7124),
            .I(N__7120));
    CascadeMux I__1369 (
            .O(N__7123),
            .I(N__7117));
    Span4Mux_v I__1368 (
            .O(N__7120),
            .I(N__7114));
    InMux I__1367 (
            .O(N__7117),
            .I(N__7111));
    Odrv4 I__1366 (
            .O(N__7114),
            .I(\U111_CYCLE_SM.TA_DISZ0 ));
    LocalMux I__1365 (
            .O(N__7111),
            .I(\U111_CYCLE_SM.TA_DISZ0 ));
    IoInMux I__1364 (
            .O(N__7106),
            .I(N__7103));
    LocalMux I__1363 (
            .O(N__7103),
            .I(N__7100));
    Span4Mux_s3_v I__1362 (
            .O(N__7100),
            .I(N__7097));
    Span4Mux_h I__1361 (
            .O(N__7097),
            .I(N__7094));
    Span4Mux_v I__1360 (
            .O(N__7094),
            .I(N__7091));
    Span4Mux_v I__1359 (
            .O(N__7091),
            .I(N__7088));
    Odrv4 I__1358 (
            .O(N__7088),
            .I(TAn_1_i));
    InMux I__1357 (
            .O(N__7085),
            .I(N__7082));
    LocalMux I__1356 (
            .O(N__7082),
            .I(N__7079));
    Span4Mux_v I__1355 (
            .O(N__7079),
            .I(N__7076));
    Sp12to4 I__1354 (
            .O(N__7076),
            .I(N__7073));
    Span12Mux_h I__1353 (
            .O(N__7073),
            .I(N__7070));
    Odrv12 I__1352 (
            .O(N__7070),
            .I(D_LM_AMIGA_in_4));
    IoInMux I__1351 (
            .O(N__7067),
            .I(N__7064));
    LocalMux I__1350 (
            .O(N__7064),
            .I(N__7061));
    IoSpan4Mux I__1349 (
            .O(N__7061),
            .I(N__7058));
    Span4Mux_s2_h I__1348 (
            .O(N__7058),
            .I(N__7055));
    Span4Mux_h I__1347 (
            .O(N__7055),
            .I(N__7052));
    Sp12to4 I__1346 (
            .O(N__7052),
            .I(N__7049));
    Span12Mux_h I__1345 (
            .O(N__7049),
            .I(N__7046));
    Odrv12 I__1344 (
            .O(N__7046),
            .I(un2_D_LM_AMIGA_4));
    InMux I__1343 (
            .O(N__7043),
            .I(N__7040));
    LocalMux I__1342 (
            .O(N__7040),
            .I(N__7037));
    Span4Mux_v I__1341 (
            .O(N__7037),
            .I(N__7034));
    Odrv4 I__1340 (
            .O(N__7034),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ));
    InMux I__1339 (
            .O(N__7031),
            .I(N__7026));
    InMux I__1338 (
            .O(N__7030),
            .I(N__7023));
    InMux I__1337 (
            .O(N__7029),
            .I(N__7020));
    LocalMux I__1336 (
            .O(N__7026),
            .I(N__7017));
    LocalMux I__1335 (
            .O(N__7023),
            .I(N__7014));
    LocalMux I__1334 (
            .O(N__7020),
            .I(N__7011));
    Span4Mux_v I__1333 (
            .O(N__7017),
            .I(N__7006));
    Span4Mux_v I__1332 (
            .O(N__7014),
            .I(N__7006));
    Span4Mux_v I__1331 (
            .O(N__7011),
            .I(N__7003));
    Sp12to4 I__1330 (
            .O(N__7006),
            .I(N__6998));
    Sp12to4 I__1329 (
            .O(N__7003),
            .I(N__6998));
    Span12Mux_h I__1328 (
            .O(N__6998),
            .I(N__6995));
    Span12Mux_v I__1327 (
            .O(N__6995),
            .I(N__6992));
    Odrv12 I__1326 (
            .O(N__6992),
            .I(D_UU_AMIGA_in_5));
    IoInMux I__1325 (
            .O(N__6989),
            .I(N__6986));
    LocalMux I__1324 (
            .O(N__6986),
            .I(N__6983));
    IoSpan4Mux I__1323 (
            .O(N__6983),
            .I(N__6980));
    Sp12to4 I__1322 (
            .O(N__6980),
            .I(N__6977));
    Span12Mux_v I__1321 (
            .O(N__6977),
            .I(N__6974));
    Span12Mux_h I__1320 (
            .O(N__6974),
            .I(N__6971));
    Odrv12 I__1319 (
            .O(N__6971),
            .I(un1_D_UU_AMIGA_5));
    InMux I__1318 (
            .O(N__6968),
            .I(N__6965));
    LocalMux I__1317 (
            .O(N__6965),
            .I(N__6960));
    InMux I__1316 (
            .O(N__6964),
            .I(N__6957));
    InMux I__1315 (
            .O(N__6963),
            .I(N__6954));
    Span4Mux_v I__1314 (
            .O(N__6960),
            .I(N__6949));
    LocalMux I__1313 (
            .O(N__6957),
            .I(N__6949));
    LocalMux I__1312 (
            .O(N__6954),
            .I(N__6946));
    Span4Mux_v I__1311 (
            .O(N__6949),
            .I(N__6943));
    Sp12to4 I__1310 (
            .O(N__6946),
            .I(N__6940));
    Sp12to4 I__1309 (
            .O(N__6943),
            .I(N__6937));
    Span12Mux_v I__1308 (
            .O(N__6940),
            .I(N__6934));
    Span12Mux_h I__1307 (
            .O(N__6937),
            .I(N__6931));
    Odrv12 I__1306 (
            .O(N__6934),
            .I(D_UM_AMIGA_in_1));
    Odrv12 I__1305 (
            .O(N__6931),
            .I(D_UM_AMIGA_in_1));
    InMux I__1304 (
            .O(N__6926),
            .I(N__6923));
    LocalMux I__1303 (
            .O(N__6923),
            .I(N__6920));
    Odrv12 I__1302 (
            .O(N__6920),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ));
    IoInMux I__1301 (
            .O(N__6917),
            .I(N__6914));
    LocalMux I__1300 (
            .O(N__6914),
            .I(N__6911));
    Span4Mux_s3_h I__1299 (
            .O(N__6911),
            .I(N__6908));
    Span4Mux_h I__1298 (
            .O(N__6908),
            .I(N__6905));
    Sp12to4 I__1297 (
            .O(N__6905),
            .I(N__6902));
    Span12Mux_s11_v I__1296 (
            .O(N__6902),
            .I(N__6899));
    Odrv12 I__1295 (
            .O(N__6899),
            .I(un1_D_UM_AMIGA_1));
    InMux I__1294 (
            .O(N__6896),
            .I(N__6893));
    LocalMux I__1293 (
            .O(N__6893),
            .I(N__6890));
    Odrv12 I__1292 (
            .O(N__6890),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ));
    InMux I__1291 (
            .O(N__6887),
            .I(N__6883));
    InMux I__1290 (
            .O(N__6886),
            .I(N__6880));
    LocalMux I__1289 (
            .O(N__6883),
            .I(N__6877));
    LocalMux I__1288 (
            .O(N__6880),
            .I(N__6874));
    Span4Mux_v I__1287 (
            .O(N__6877),
            .I(N__6871));
    Span4Mux_v I__1286 (
            .O(N__6874),
            .I(N__6868));
    Sp12to4 I__1285 (
            .O(N__6871),
            .I(N__6864));
    Span4Mux_v I__1284 (
            .O(N__6868),
            .I(N__6861));
    InMux I__1283 (
            .O(N__6867),
            .I(N__6858));
    Span12Mux_h I__1282 (
            .O(N__6864),
            .I(N__6855));
    Sp12to4 I__1281 (
            .O(N__6861),
            .I(N__6850));
    LocalMux I__1280 (
            .O(N__6858),
            .I(N__6850));
    Span12Mux_v I__1279 (
            .O(N__6855),
            .I(N__6847));
    Span12Mux_h I__1278 (
            .O(N__6850),
            .I(N__6844));
    Odrv12 I__1277 (
            .O(N__6847),
            .I(D_UU_AMIGA_in_0));
    Odrv12 I__1276 (
            .O(N__6844),
            .I(D_UU_AMIGA_in_0));
    IoInMux I__1275 (
            .O(N__6839),
            .I(N__6836));
    LocalMux I__1274 (
            .O(N__6836),
            .I(N__6833));
    Span4Mux_s3_v I__1273 (
            .O(N__6833),
            .I(N__6830));
    Span4Mux_v I__1272 (
            .O(N__6830),
            .I(N__6827));
    Sp12to4 I__1271 (
            .O(N__6827),
            .I(N__6824));
    Span12Mux_h I__1270 (
            .O(N__6824),
            .I(N__6821));
    Odrv12 I__1269 (
            .O(N__6821),
            .I(un1_D_UU_AMIGA_0));
    IoInMux I__1268 (
            .O(N__6818),
            .I(N__6815));
    LocalMux I__1267 (
            .O(N__6815),
            .I(N__6812));
    Odrv12 I__1266 (
            .O(N__6812),
            .I(LBENn_c_i_0));
    InMux I__1265 (
            .O(N__6809),
            .I(N__6806));
    LocalMux I__1264 (
            .O(N__6806),
            .I(N__6803));
    Span4Mux_v I__1263 (
            .O(N__6803),
            .I(N__6800));
    Sp12to4 I__1262 (
            .O(N__6800),
            .I(N__6797));
    Span12Mux_h I__1261 (
            .O(N__6797),
            .I(N__6794));
    Odrv12 I__1260 (
            .O(N__6794),
            .I(D_LL_AMIGA_in_7));
    IoInMux I__1259 (
            .O(N__6791),
            .I(N__6788));
    LocalMux I__1258 (
            .O(N__6788),
            .I(N__6785));
    IoSpan4Mux I__1257 (
            .O(N__6785),
            .I(N__6782));
    Span4Mux_s3_h I__1256 (
            .O(N__6782),
            .I(N__6779));
    Sp12to4 I__1255 (
            .O(N__6779),
            .I(N__6776));
    Span12Mux_h I__1254 (
            .O(N__6776),
            .I(N__6773));
    Odrv12 I__1253 (
            .O(N__6773),
            .I(un2_D_LL_AMIGA_7));
    InMux I__1252 (
            .O(N__6770),
            .I(N__6767));
    LocalMux I__1251 (
            .O(N__6767),
            .I(N__6761));
    InMux I__1250 (
            .O(N__6766),
            .I(N__6757));
    InMux I__1249 (
            .O(N__6765),
            .I(N__6754));
    InMux I__1248 (
            .O(N__6764),
            .I(N__6751));
    Span12Mux_s6_h I__1247 (
            .O(N__6761),
            .I(N__6748));
    InMux I__1246 (
            .O(N__6760),
            .I(N__6745));
    LocalMux I__1245 (
            .O(N__6757),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1244 (
            .O(N__6754),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1243 (
            .O(N__6751),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    Odrv12 I__1242 (
            .O(N__6748),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1241 (
            .O(N__6745),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    CascadeMux I__1240 (
            .O(N__6734),
            .I(N__6731));
    InMux I__1239 (
            .O(N__6731),
            .I(N__6728));
    LocalMux I__1238 (
            .O(N__6728),
            .I(N__6725));
    Odrv4 I__1237 (
            .O(N__6725),
            .I(\U111_CYCLE_SM.N_119_0 ));
    InMux I__1236 (
            .O(N__6722),
            .I(N__6719));
    LocalMux I__1235 (
            .O(N__6719),
            .I(N__6716));
    Odrv4 I__1234 (
            .O(N__6716),
            .I(\U111_CYCLE_SM.N_117_0 ));
    InMux I__1233 (
            .O(N__6713),
            .I(N__6702));
    InMux I__1232 (
            .O(N__6712),
            .I(N__6702));
    InMux I__1231 (
            .O(N__6711),
            .I(N__6702));
    InMux I__1230 (
            .O(N__6710),
            .I(N__6697));
    InMux I__1229 (
            .O(N__6709),
            .I(N__6697));
    LocalMux I__1228 (
            .O(N__6702),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ));
    LocalMux I__1227 (
            .O(N__6697),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ));
    CascadeMux I__1226 (
            .O(N__6692),
            .I(\U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_cascade_ ));
    InMux I__1225 (
            .O(N__6689),
            .I(N__6686));
    LocalMux I__1224 (
            .O(N__6686),
            .I(N__6682));
    InMux I__1223 (
            .O(N__6685),
            .I(N__6679));
    Odrv4 I__1222 (
            .O(N__6682),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    LocalMux I__1221 (
            .O(N__6679),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    CascadeMux I__1220 (
            .O(N__6674),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1_cascade_ ));
    InMux I__1219 (
            .O(N__6671),
            .I(N__6668));
    LocalMux I__1218 (
            .O(N__6668),
            .I(N__6665));
    Span4Mux_h I__1217 (
            .O(N__6665),
            .I(N__6659));
    InMux I__1216 (
            .O(N__6664),
            .I(N__6656));
    InMux I__1215 (
            .O(N__6663),
            .I(N__6653));
    InMux I__1214 (
            .O(N__6662),
            .I(N__6650));
    Odrv4 I__1213 (
            .O(N__6659),
            .I(\U111_CYCLE_SM.BURST_COUNT_0_sqmuxa ));
    LocalMux I__1212 (
            .O(N__6656),
            .I(\U111_CYCLE_SM.BURST_COUNT_0_sqmuxa ));
    LocalMux I__1211 (
            .O(N__6653),
            .I(\U111_CYCLE_SM.BURST_COUNT_0_sqmuxa ));
    LocalMux I__1210 (
            .O(N__6650),
            .I(\U111_CYCLE_SM.BURST_COUNT_0_sqmuxa ));
    InMux I__1209 (
            .O(N__6641),
            .I(N__6634));
    InMux I__1208 (
            .O(N__6640),
            .I(N__6627));
    InMux I__1207 (
            .O(N__6639),
            .I(N__6627));
    InMux I__1206 (
            .O(N__6638),
            .I(N__6627));
    InMux I__1205 (
            .O(N__6637),
            .I(N__6624));
    LocalMux I__1204 (
            .O(N__6634),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ));
    LocalMux I__1203 (
            .O(N__6627),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ));
    LocalMux I__1202 (
            .O(N__6624),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ));
    InMux I__1201 (
            .O(N__6617),
            .I(N__6612));
    InMux I__1200 (
            .O(N__6616),
            .I(N__6609));
    InMux I__1199 (
            .O(N__6615),
            .I(N__6606));
    LocalMux I__1198 (
            .O(N__6612),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_0 ));
    LocalMux I__1197 (
            .O(N__6609),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_0 ));
    LocalMux I__1196 (
            .O(N__6606),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_0 ));
    InMux I__1195 (
            .O(N__6599),
            .I(N__6592));
    InMux I__1194 (
            .O(N__6598),
            .I(N__6589));
    InMux I__1193 (
            .O(N__6597),
            .I(N__6584));
    InMux I__1192 (
            .O(N__6596),
            .I(N__6584));
    InMux I__1191 (
            .O(N__6595),
            .I(N__6581));
    LocalMux I__1190 (
            .O(N__6592),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    LocalMux I__1189 (
            .O(N__6589),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    LocalMux I__1188 (
            .O(N__6584),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    LocalMux I__1187 (
            .O(N__6581),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    CascadeMux I__1186 (
            .O(N__6572),
            .I(\U111_CYCLE_SM.N_131_cascade_ ));
    InMux I__1185 (
            .O(N__6569),
            .I(N__6566));
    LocalMux I__1184 (
            .O(N__6566),
            .I(\U111_CYCLE_SM.CYCLE_STATE_srsts_0_1_0 ));
    InMux I__1183 (
            .O(N__6563),
            .I(N__6560));
    LocalMux I__1182 (
            .O(N__6560),
            .I(\U111_CYCLE_SM.TS_EN6 ));
    InMux I__1181 (
            .O(N__6557),
            .I(N__6554));
    LocalMux I__1180 (
            .O(N__6554),
            .I(N__6550));
    InMux I__1179 (
            .O(N__6553),
            .I(N__6547));
    Odrv4 I__1178 (
            .O(N__6550),
            .I(\U111_CYCLE_SM.N_144 ));
    LocalMux I__1177 (
            .O(N__6547),
            .I(\U111_CYCLE_SM.N_144 ));
    InMux I__1176 (
            .O(N__6542),
            .I(N__6539));
    LocalMux I__1175 (
            .O(N__6539),
            .I(N__6536));
    Span12Mux_s9_v I__1174 (
            .O(N__6536),
            .I(N__6533));
    Odrv12 I__1173 (
            .O(N__6533),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ));
    InMux I__1172 (
            .O(N__6530),
            .I(N__6527));
    LocalMux I__1171 (
            .O(N__6527),
            .I(N__6524));
    Span4Mux_v I__1170 (
            .O(N__6524),
            .I(N__6519));
    InMux I__1169 (
            .O(N__6523),
            .I(N__6516));
    InMux I__1168 (
            .O(N__6522),
            .I(N__6513));
    Span4Mux_v I__1167 (
            .O(N__6519),
            .I(N__6510));
    LocalMux I__1166 (
            .O(N__6516),
            .I(N__6507));
    LocalMux I__1165 (
            .O(N__6513),
            .I(N__6504));
    Span4Mux_v I__1164 (
            .O(N__6510),
            .I(N__6501));
    Span4Mux_v I__1163 (
            .O(N__6507),
            .I(N__6498));
    Span12Mux_h I__1162 (
            .O(N__6504),
            .I(N__6495));
    Sp12to4 I__1161 (
            .O(N__6501),
            .I(N__6490));
    Sp12to4 I__1160 (
            .O(N__6498),
            .I(N__6490));
    Span12Mux_v I__1159 (
            .O(N__6495),
            .I(N__6485));
    Span12Mux_h I__1158 (
            .O(N__6490),
            .I(N__6485));
    Odrv12 I__1157 (
            .O(N__6485),
            .I(D_UU_AMIGA_in_1));
    IoInMux I__1156 (
            .O(N__6482),
            .I(N__6479));
    LocalMux I__1155 (
            .O(N__6479),
            .I(N__6476));
    Span4Mux_s3_h I__1154 (
            .O(N__6476),
            .I(N__6473));
    Span4Mux_h I__1153 (
            .O(N__6473),
            .I(N__6470));
    Sp12to4 I__1152 (
            .O(N__6470),
            .I(N__6467));
    Span12Mux_s8_v I__1151 (
            .O(N__6467),
            .I(N__6464));
    Odrv12 I__1150 (
            .O(N__6464),
            .I(un1_D_UU_AMIGA_1));
    InMux I__1149 (
            .O(N__6461),
            .I(N__6458));
    LocalMux I__1148 (
            .O(N__6458),
            .I(N__6455));
    Span12Mux_v I__1147 (
            .O(N__6455),
            .I(N__6452));
    Span12Mux_h I__1146 (
            .O(N__6452),
            .I(N__6449));
    Odrv12 I__1145 (
            .O(N__6449),
            .I(D_UM_040_in_3));
    InMux I__1144 (
            .O(N__6446),
            .I(N__6442));
    IoInMux I__1143 (
            .O(N__6445),
            .I(N__6439));
    LocalMux I__1142 (
            .O(N__6442),
            .I(N__6436));
    LocalMux I__1141 (
            .O(N__6439),
            .I(N__6433));
    Span4Mux_v I__1140 (
            .O(N__6436),
            .I(N__6430));
    Span4Mux_s3_h I__1139 (
            .O(N__6433),
            .I(N__6427));
    Sp12to4 I__1138 (
            .O(N__6430),
            .I(N__6424));
    Sp12to4 I__1137 (
            .O(N__6427),
            .I(N__6421));
    Span12Mux_h I__1136 (
            .O(N__6424),
            .I(N__6418));
    Span12Mux_v I__1135 (
            .O(N__6421),
            .I(N__6415));
    Span12Mux_v I__1134 (
            .O(N__6418),
            .I(N__6412));
    Span12Mux_h I__1133 (
            .O(N__6415),
            .I(N__6409));
    Span12Mux_v I__1132 (
            .O(N__6412),
            .I(N__6404));
    Span12Mux_h I__1131 (
            .O(N__6409),
            .I(N__6404));
    Odrv12 I__1130 (
            .O(N__6404),
            .I(D_LL_040_in_3));
    IoInMux I__1129 (
            .O(N__6401),
            .I(N__6398));
    LocalMux I__1128 (
            .O(N__6398),
            .I(N__6395));
    IoSpan4Mux I__1127 (
            .O(N__6395),
            .I(N__6392));
    Span4Mux_s2_h I__1126 (
            .O(N__6392),
            .I(N__6389));
    Sp12to4 I__1125 (
            .O(N__6389),
            .I(N__6386));
    Odrv12 I__1124 (
            .O(N__6386),
            .I(un1_D_UM_040_3));
    IoInMux I__1123 (
            .O(N__6383),
            .I(N__6380));
    LocalMux I__1122 (
            .O(N__6380),
            .I(N__6377));
    IoSpan4Mux I__1121 (
            .O(N__6377),
            .I(N__6374));
    IoSpan4Mux I__1120 (
            .O(N__6374),
            .I(N__6370));
    InMux I__1119 (
            .O(N__6373),
            .I(N__6367));
    Span4Mux_s2_h I__1118 (
            .O(N__6370),
            .I(N__6364));
    LocalMux I__1117 (
            .O(N__6367),
            .I(N__6361));
    Sp12to4 I__1116 (
            .O(N__6364),
            .I(N__6358));
    Span12Mux_s10_v I__1115 (
            .O(N__6361),
            .I(N__6355));
    Span12Mux_h I__1114 (
            .O(N__6358),
            .I(N__6350));
    Span12Mux_v I__1113 (
            .O(N__6355),
            .I(N__6350));
    Span12Mux_h I__1112 (
            .O(N__6350),
            .I(N__6347));
    Odrv12 I__1111 (
            .O(N__6347),
            .I(D_LM_040_in_3));
    InMux I__1110 (
            .O(N__6344),
            .I(N__6341));
    LocalMux I__1109 (
            .O(N__6341),
            .I(N__6338));
    Span4Mux_v I__1108 (
            .O(N__6338),
            .I(N__6335));
    Span4Mux_h I__1107 (
            .O(N__6335),
            .I(N__6332));
    Sp12to4 I__1106 (
            .O(N__6332),
            .I(N__6329));
    Span12Mux_h I__1105 (
            .O(N__6329),
            .I(N__6326));
    Odrv12 I__1104 (
            .O(N__6326),
            .I(D_UU_040_in_3));
    IoInMux I__1103 (
            .O(N__6323),
            .I(N__6320));
    LocalMux I__1102 (
            .O(N__6320),
            .I(N__6317));
    Span12Mux_s6_v I__1101 (
            .O(N__6317),
            .I(N__6314));
    Odrv12 I__1100 (
            .O(N__6314),
            .I(un1_D_UU_040_3));
    InMux I__1099 (
            .O(N__6311),
            .I(N__6308));
    LocalMux I__1098 (
            .O(N__6308),
            .I(\U111_CYCLE_SM.N_124_0 ));
    CascadeMux I__1097 (
            .O(N__6305),
            .I(\U111_CYCLE_SM.N_132_cascade_ ));
    CascadeMux I__1096 (
            .O(N__6302),
            .I(N__6299));
    InMux I__1095 (
            .O(N__6299),
            .I(N__6295));
    InMux I__1094 (
            .O(N__6298),
            .I(N__6292));
    LocalMux I__1093 (
            .O(N__6295),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_1 ));
    LocalMux I__1092 (
            .O(N__6292),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_1 ));
    CascadeMux I__1091 (
            .O(N__6287),
            .I(N__6284));
    InMux I__1090 (
            .O(N__6284),
            .I(N__6281));
    LocalMux I__1089 (
            .O(N__6281),
            .I(N__6278));
    Span4Mux_v I__1088 (
            .O(N__6278),
            .I(N__6275));
    Span4Mux_v I__1087 (
            .O(N__6275),
            .I(N__6271));
    IoInMux I__1086 (
            .O(N__6274),
            .I(N__6268));
    Sp12to4 I__1085 (
            .O(N__6271),
            .I(N__6265));
    LocalMux I__1084 (
            .O(N__6268),
            .I(N__6262));
    Span12Mux_h I__1083 (
            .O(N__6265),
            .I(N__6259));
    IoSpan4Mux I__1082 (
            .O(N__6262),
            .I(N__6256));
    Odrv12 I__1081 (
            .O(N__6259),
            .I(TBIn_c));
    Odrv4 I__1080 (
            .O(N__6256),
            .I(TBIn_c));
    InMux I__1079 (
            .O(N__6251),
            .I(N__6248));
    LocalMux I__1078 (
            .O(N__6248),
            .I(\U111_CYCLE_SM.un7_CYCLE_STATE_0 ));
    CascadeMux I__1077 (
            .O(N__6245),
            .I(\U111_CYCLE_SM.un7_CYCLE_STATE_0_cascade_ ));
    CascadeMux I__1076 (
            .O(N__6242),
            .I(\U111_CYCLE_SM.CYCLE_STATE_srsts_i_1_2_cascade_ ));
    InMux I__1075 (
            .O(N__6239),
            .I(N__6229));
    InMux I__1074 (
            .O(N__6238),
            .I(N__6229));
    InMux I__1073 (
            .O(N__6237),
            .I(N__6229));
    InMux I__1072 (
            .O(N__6236),
            .I(N__6225));
    LocalMux I__1071 (
            .O(N__6229),
            .I(N__6222));
    InMux I__1070 (
            .O(N__6228),
            .I(N__6219));
    LocalMux I__1069 (
            .O(N__6225),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    Odrv4 I__1068 (
            .O(N__6222),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1067 (
            .O(N__6219),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    CascadeMux I__1066 (
            .O(N__6212),
            .I(N__6209));
    InMux I__1065 (
            .O(N__6209),
            .I(N__6203));
    InMux I__1064 (
            .O(N__6208),
            .I(N__6198));
    InMux I__1063 (
            .O(N__6207),
            .I(N__6198));
    InMux I__1062 (
            .O(N__6206),
            .I(N__6195));
    LocalMux I__1061 (
            .O(N__6203),
            .I(\U111_CYCLE_SM.PORT_MISMATCHZ0 ));
    LocalMux I__1060 (
            .O(N__6198),
            .I(\U111_CYCLE_SM.PORT_MISMATCHZ0 ));
    LocalMux I__1059 (
            .O(N__6195),
            .I(\U111_CYCLE_SM.PORT_MISMATCHZ0 ));
    InMux I__1058 (
            .O(N__6188),
            .I(N__6185));
    LocalMux I__1057 (
            .O(N__6185),
            .I(N__6177));
    InMux I__1056 (
            .O(N__6184),
            .I(N__6174));
    InMux I__1055 (
            .O(N__6183),
            .I(N__6171));
    InMux I__1054 (
            .O(N__6182),
            .I(N__6164));
    InMux I__1053 (
            .O(N__6181),
            .I(N__6164));
    InMux I__1052 (
            .O(N__6180),
            .I(N__6164));
    Odrv4 I__1051 (
            .O(N__6177),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    LocalMux I__1050 (
            .O(N__6174),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    LocalMux I__1049 (
            .O(N__6171),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    LocalMux I__1048 (
            .O(N__6164),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    InMux I__1047 (
            .O(N__6155),
            .I(N__6149));
    InMux I__1046 (
            .O(N__6154),
            .I(N__6149));
    LocalMux I__1045 (
            .O(N__6149),
            .I(N__6146));
    Sp12to4 I__1044 (
            .O(N__6146),
            .I(N__6143));
    Span12Mux_v I__1043 (
            .O(N__6143),
            .I(N__6140));
    Span12Mux_h I__1042 (
            .O(N__6140),
            .I(N__6137));
    Odrv12 I__1041 (
            .O(N__6137),
            .I(SIZ_c_1));
    CascadeMux I__1040 (
            .O(N__6134),
            .I(N__6130));
    CascadeMux I__1039 (
            .O(N__6133),
            .I(N__6127));
    InMux I__1038 (
            .O(N__6130),
            .I(N__6122));
    InMux I__1037 (
            .O(N__6127),
            .I(N__6122));
    LocalMux I__1036 (
            .O(N__6122),
            .I(N__6119));
    Span12Mux_v I__1035 (
            .O(N__6119),
            .I(N__6116));
    Span12Mux_h I__1034 (
            .O(N__6116),
            .I(N__6113));
    Odrv12 I__1033 (
            .O(N__6113),
            .I(SIZ_c_0));
    CascadeMux I__1032 (
            .O(N__6110),
            .I(N__6107));
    InMux I__1031 (
            .O(N__6107),
            .I(N__6104));
    LocalMux I__1030 (
            .O(N__6104),
            .I(N__6101));
    Span4Mux_v I__1029 (
            .O(N__6101),
            .I(N__6098));
    Span4Mux_h I__1028 (
            .O(N__6098),
            .I(N__6095));
    Odrv4 I__1027 (
            .O(N__6095),
            .I(\U111_CYCLE_SM.FLIP_WORD_2 ));
    InMux I__1026 (
            .O(N__6092),
            .I(N__6089));
    LocalMux I__1025 (
            .O(N__6089),
            .I(N__6085));
    InMux I__1024 (
            .O(N__6088),
            .I(N__6081));
    Span4Mux_v I__1023 (
            .O(N__6085),
            .I(N__6078));
    InMux I__1022 (
            .O(N__6084),
            .I(N__6075));
    LocalMux I__1021 (
            .O(N__6081),
            .I(N__6072));
    Sp12to4 I__1020 (
            .O(N__6078),
            .I(N__6067));
    LocalMux I__1019 (
            .O(N__6075),
            .I(N__6067));
    Span4Mux_h I__1018 (
            .O(N__6072),
            .I(N__6064));
    Span12Mux_h I__1017 (
            .O(N__6067),
            .I(N__6061));
    Span4Mux_v I__1016 (
            .O(N__6064),
            .I(N__6058));
    Span12Mux_v I__1015 (
            .O(N__6061),
            .I(N__6055));
    Span4Mux_v I__1014 (
            .O(N__6058),
            .I(N__6052));
    Odrv12 I__1013 (
            .O(N__6055),
            .I(PORTSIZE_c));
    Odrv4 I__1012 (
            .O(N__6052),
            .I(PORTSIZE_c));
    InMux I__1011 (
            .O(N__6047),
            .I(N__6040));
    InMux I__1010 (
            .O(N__6046),
            .I(N__6040));
    InMux I__1009 (
            .O(N__6045),
            .I(N__6037));
    LocalMux I__1008 (
            .O(N__6040),
            .I(\U111_CYCLE_SM.LW_TRANSZ0 ));
    LocalMux I__1007 (
            .O(N__6037),
            .I(\U111_CYCLE_SM.LW_TRANSZ0 ));
    InMux I__1006 (
            .O(N__6032),
            .I(N__6029));
    LocalMux I__1005 (
            .O(N__6029),
            .I(\U111_CYCLE_SM.PORT_MISMATCH_2 ));
    InMux I__1004 (
            .O(N__6026),
            .I(N__6020));
    InMux I__1003 (
            .O(N__6025),
            .I(N__6020));
    LocalMux I__1002 (
            .O(N__6020),
            .I(N__6017));
    Span4Mux_h I__1001 (
            .O(N__6017),
            .I(N__6014));
    Sp12to4 I__1000 (
            .O(N__6014),
            .I(N__6011));
    Span12Mux_v I__999 (
            .O(N__6011),
            .I(N__6007));
    InMux I__998 (
            .O(N__6010),
            .I(N__6004));
    Odrv12 I__997 (
            .O(N__6007),
            .I(\U111_CYCLE_SM.A2_ENZ0 ));
    LocalMux I__996 (
            .O(N__6004),
            .I(\U111_CYCLE_SM.A2_ENZ0 ));
    InMux I__995 (
            .O(N__5999),
            .I(N__5996));
    LocalMux I__994 (
            .O(N__5996),
            .I(N__5993));
    Span4Mux_v I__993 (
            .O(N__5993),
            .I(N__5990));
    Sp12to4 I__992 (
            .O(N__5990),
            .I(N__5987));
    Odrv12 I__991 (
            .O(N__5987),
            .I(D_LM_AMIGA_in_5));
    IoInMux I__990 (
            .O(N__5984),
            .I(N__5981));
    LocalMux I__989 (
            .O(N__5981),
            .I(N__5978));
    IoSpan4Mux I__988 (
            .O(N__5978),
            .I(N__5975));
    Sp12to4 I__987 (
            .O(N__5975),
            .I(N__5972));
    Span12Mux_s7_h I__986 (
            .O(N__5972),
            .I(N__5969));
    Span12Mux_h I__985 (
            .O(N__5969),
            .I(N__5966));
    Odrv12 I__984 (
            .O(N__5966),
            .I(un2_D_LM_AMIGA_5));
    IoInMux I__983 (
            .O(N__5963),
            .I(N__5960));
    LocalMux I__982 (
            .O(N__5960),
            .I(N__5956));
    InMux I__981 (
            .O(N__5959),
            .I(N__5953));
    IoSpan4Mux I__980 (
            .O(N__5956),
            .I(N__5950));
    LocalMux I__979 (
            .O(N__5953),
            .I(N__5947));
    Span4Mux_s2_h I__978 (
            .O(N__5950),
            .I(N__5944));
    Sp12to4 I__977 (
            .O(N__5947),
            .I(N__5941));
    Span4Mux_v I__976 (
            .O(N__5944),
            .I(N__5938));
    Span12Mux_v I__975 (
            .O(N__5941),
            .I(N__5935));
    Sp12to4 I__974 (
            .O(N__5938),
            .I(N__5932));
    Span12Mux_v I__973 (
            .O(N__5935),
            .I(N__5929));
    Span12Mux_s9_h I__972 (
            .O(N__5932),
            .I(N__5926));
    Span12Mux_h I__971 (
            .O(N__5929),
            .I(N__5923));
    Span12Mux_h I__970 (
            .O(N__5926),
            .I(N__5920));
    Odrv12 I__969 (
            .O(N__5923),
            .I(D_LM_040_in_0));
    Odrv12 I__968 (
            .O(N__5920),
            .I(D_LM_040_in_0));
    InMux I__967 (
            .O(N__5915),
            .I(N__5912));
    LocalMux I__966 (
            .O(N__5912),
            .I(N__5909));
    Span4Mux_v I__965 (
            .O(N__5909),
            .I(N__5906));
    Span4Mux_h I__964 (
            .O(N__5906),
            .I(N__5903));
    Sp12to4 I__963 (
            .O(N__5903),
            .I(N__5900));
    Span12Mux_h I__962 (
            .O(N__5900),
            .I(N__5897));
    Odrv12 I__961 (
            .O(N__5897),
            .I(D_UU_040_in_0));
    IoInMux I__960 (
            .O(N__5894),
            .I(N__5891));
    LocalMux I__959 (
            .O(N__5891),
            .I(N__5888));
    Span12Mux_s6_v I__958 (
            .O(N__5888),
            .I(N__5885));
    Odrv12 I__957 (
            .O(N__5885),
            .I(un1_D_UU_040_0));
    InMux I__956 (
            .O(N__5882),
            .I(N__5879));
    LocalMux I__955 (
            .O(N__5879),
            .I(N__5876));
    Span4Mux_v I__954 (
            .O(N__5876),
            .I(N__5873));
    Span4Mux_h I__953 (
            .O(N__5873),
            .I(N__5870));
    Sp12to4 I__952 (
            .O(N__5870),
            .I(N__5867));
    Odrv12 I__951 (
            .O(N__5867),
            .I(D_LL_AMIGA_in_6));
    IoInMux I__950 (
            .O(N__5864),
            .I(N__5861));
    LocalMux I__949 (
            .O(N__5861),
            .I(N__5858));
    Span4Mux_s3_h I__948 (
            .O(N__5858),
            .I(N__5855));
    Span4Mux_v I__947 (
            .O(N__5855),
            .I(N__5852));
    Span4Mux_v I__946 (
            .O(N__5852),
            .I(N__5849));
    Sp12to4 I__945 (
            .O(N__5849),
            .I(N__5846));
    Span12Mux_s10_h I__944 (
            .O(N__5846),
            .I(N__5843));
    Odrv12 I__943 (
            .O(N__5843),
            .I(un2_D_LL_AMIGA_6));
    InMux I__942 (
            .O(N__5840),
            .I(N__5837));
    LocalMux I__941 (
            .O(N__5837),
            .I(N__5834));
    Span4Mux_v I__940 (
            .O(N__5834),
            .I(N__5831));
    Span4Mux_h I__939 (
            .O(N__5831),
            .I(N__5828));
    Sp12to4 I__938 (
            .O(N__5828),
            .I(N__5825));
    Span12Mux_h I__937 (
            .O(N__5825),
            .I(N__5822));
    Odrv12 I__936 (
            .O(N__5822),
            .I(D_UU_040_in_6));
    IoInMux I__935 (
            .O(N__5819),
            .I(N__5816));
    LocalMux I__934 (
            .O(N__5816),
            .I(N__5812));
    InMux I__933 (
            .O(N__5815),
            .I(N__5809));
    Span4Mux_s2_h I__932 (
            .O(N__5812),
            .I(N__5806));
    LocalMux I__931 (
            .O(N__5809),
            .I(N__5803));
    Span4Mux_v I__930 (
            .O(N__5806),
            .I(N__5800));
    Span4Mux_v I__929 (
            .O(N__5803),
            .I(N__5797));
    Sp12to4 I__928 (
            .O(N__5800),
            .I(N__5794));
    Span4Mux_v I__927 (
            .O(N__5797),
            .I(N__5791));
    Span12Mux_h I__926 (
            .O(N__5794),
            .I(N__5786));
    Sp12to4 I__925 (
            .O(N__5791),
            .I(N__5786));
    Span12Mux_h I__924 (
            .O(N__5786),
            .I(N__5783));
    Odrv12 I__923 (
            .O(N__5783),
            .I(D_LM_040_in_6));
    IoInMux I__922 (
            .O(N__5780),
            .I(N__5777));
    LocalMux I__921 (
            .O(N__5777),
            .I(N__5774));
    Span4Mux_s3_v I__920 (
            .O(N__5774),
            .I(N__5771));
    Span4Mux_h I__919 (
            .O(N__5771),
            .I(N__5768));
    Span4Mux_h I__918 (
            .O(N__5768),
            .I(N__5765));
    Odrv4 I__917 (
            .O(N__5765),
            .I(un1_D_UU_040_6));
    InMux I__916 (
            .O(N__5762),
            .I(N__5759));
    LocalMux I__915 (
            .O(N__5759),
            .I(N__5756));
    Span4Mux_v I__914 (
            .O(N__5756),
            .I(N__5753));
    Sp12to4 I__913 (
            .O(N__5753),
            .I(N__5750));
    Odrv12 I__912 (
            .O(N__5750),
            .I(D_LL_AMIGA_in_3));
    IoInMux I__911 (
            .O(N__5747),
            .I(N__5744));
    LocalMux I__910 (
            .O(N__5744),
            .I(N__5741));
    Span12Mux_s7_h I__909 (
            .O(N__5741),
            .I(N__5738));
    Span12Mux_h I__908 (
            .O(N__5738),
            .I(N__5735));
    Odrv12 I__907 (
            .O(N__5735),
            .I(un2_D_LL_AMIGA_3));
    CascadeMux I__906 (
            .O(N__5732),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa_cascade_ ));
    InMux I__905 (
            .O(N__5729),
            .I(N__5725));
    InMux I__904 (
            .O(N__5728),
            .I(N__5722));
    LocalMux I__903 (
            .O(N__5725),
            .I(\U111_CYCLE_SM.un1_CYCLE_STATE_0 ));
    LocalMux I__902 (
            .O(N__5722),
            .I(\U111_CYCLE_SM.un1_CYCLE_STATE_0 ));
    CascadeMux I__901 (
            .O(N__5717),
            .I(N__5714));
    InMux I__900 (
            .O(N__5714),
            .I(N__5711));
    LocalMux I__899 (
            .O(N__5711),
            .I(\U111_CYCLE_SM.TS_EN_6 ));
    IoInMux I__898 (
            .O(N__5708),
            .I(N__5704));
    IoInMux I__897 (
            .O(N__5707),
            .I(N__5701));
    LocalMux I__896 (
            .O(N__5704),
            .I(N__5698));
    LocalMux I__895 (
            .O(N__5701),
            .I(N__5695));
    Span12Mux_s6_v I__894 (
            .O(N__5698),
            .I(N__5690));
    Span12Mux_s6_v I__893 (
            .O(N__5695),
            .I(N__5690));
    Odrv12 I__892 (
            .O(N__5690),
            .I(CONSTANT_ONE_NET));
    InMux I__891 (
            .O(N__5687),
            .I(N__5684));
    LocalMux I__890 (
            .O(N__5684),
            .I(N__5681));
    Span4Mux_v I__889 (
            .O(N__5681),
            .I(N__5678));
    Sp12to4 I__888 (
            .O(N__5678),
            .I(N__5675));
    Span12Mux_h I__887 (
            .O(N__5675),
            .I(N__5672));
    Odrv12 I__886 (
            .O(N__5672),
            .I(D_LL_AMIGA_in_2));
    IoInMux I__885 (
            .O(N__5669),
            .I(N__5666));
    LocalMux I__884 (
            .O(N__5666),
            .I(N__5663));
    Span4Mux_s2_h I__883 (
            .O(N__5663),
            .I(N__5660));
    Sp12to4 I__882 (
            .O(N__5660),
            .I(N__5657));
    Span12Mux_s8_v I__881 (
            .O(N__5657),
            .I(N__5654));
    Span12Mux_h I__880 (
            .O(N__5654),
            .I(N__5651));
    Odrv12 I__879 (
            .O(N__5651),
            .I(un2_D_LL_AMIGA_2));
    InMux I__878 (
            .O(N__5648),
            .I(N__5645));
    LocalMux I__877 (
            .O(N__5645),
            .I(N__5642));
    Span4Mux_v I__876 (
            .O(N__5642),
            .I(N__5639));
    Sp12to4 I__875 (
            .O(N__5639),
            .I(N__5636));
    Span12Mux_h I__874 (
            .O(N__5636),
            .I(N__5633));
    Odrv12 I__873 (
            .O(N__5633),
            .I(D_LM_AMIGA_in_0));
    IoInMux I__872 (
            .O(N__5630),
            .I(N__5627));
    LocalMux I__871 (
            .O(N__5627),
            .I(N__5624));
    IoSpan4Mux I__870 (
            .O(N__5624),
            .I(N__5621));
    Span4Mux_s3_h I__869 (
            .O(N__5621),
            .I(N__5618));
    Sp12to4 I__868 (
            .O(N__5618),
            .I(N__5615));
    Span12Mux_s8_h I__867 (
            .O(N__5615),
            .I(N__5612));
    Span12Mux_h I__866 (
            .O(N__5612),
            .I(N__5609));
    Odrv12 I__865 (
            .O(N__5609),
            .I(un2_D_LM_AMIGA_0));
    IoInMux I__864 (
            .O(N__5606),
            .I(N__5603));
    LocalMux I__863 (
            .O(N__5603),
            .I(N__5600));
    Span12Mux_s5_v I__862 (
            .O(N__5600),
            .I(N__5597));
    Odrv12 I__861 (
            .O(N__5597),
            .I(TSn_c));
    InMux I__860 (
            .O(N__5594),
            .I(N__5590));
    InMux I__859 (
            .O(N__5593),
            .I(N__5587));
    LocalMux I__858 (
            .O(N__5590),
            .I(\U111_CYCLE_SM.TS_ENZ0 ));
    LocalMux I__857 (
            .O(N__5587),
            .I(\U111_CYCLE_SM.TS_ENZ0 ));
    InMux I__856 (
            .O(N__5582),
            .I(N__5579));
    LocalMux I__855 (
            .O(N__5579),
            .I(N__5576));
    Span4Mux_v I__854 (
            .O(N__5576),
            .I(N__5573));
    Sp12to4 I__853 (
            .O(N__5573),
            .I(N__5570));
    Span12Mux_h I__852 (
            .O(N__5570),
            .I(N__5567));
    Span12Mux_v I__851 (
            .O(N__5567),
            .I(N__5564));
    Odrv12 I__850 (
            .O(N__5564),
            .I(D_UM_040_in_1));
    IoInMux I__849 (
            .O(N__5561),
            .I(N__5558));
    LocalMux I__848 (
            .O(N__5558),
            .I(N__5554));
    InMux I__847 (
            .O(N__5557),
            .I(N__5551));
    Span4Mux_s3_h I__846 (
            .O(N__5554),
            .I(N__5548));
    LocalMux I__845 (
            .O(N__5551),
            .I(N__5545));
    Sp12to4 I__844 (
            .O(N__5548),
            .I(N__5542));
    Span12Mux_v I__843 (
            .O(N__5545),
            .I(N__5539));
    Span12Mux_v I__842 (
            .O(N__5542),
            .I(N__5536));
    Span12Mux_v I__841 (
            .O(N__5539),
            .I(N__5533));
    Span12Mux_h I__840 (
            .O(N__5536),
            .I(N__5530));
    Span12Mux_h I__839 (
            .O(N__5533),
            .I(N__5527));
    Span12Mux_h I__838 (
            .O(N__5530),
            .I(N__5524));
    Odrv12 I__837 (
            .O(N__5527),
            .I(D_LL_040_in_1));
    Odrv12 I__836 (
            .O(N__5524),
            .I(D_LL_040_in_1));
    IoInMux I__835 (
            .O(N__5519),
            .I(N__5516));
    LocalMux I__834 (
            .O(N__5516),
            .I(N__5513));
    Span4Mux_s3_h I__833 (
            .O(N__5513),
            .I(N__5510));
    Span4Mux_h I__832 (
            .O(N__5510),
            .I(N__5507));
    Span4Mux_h I__831 (
            .O(N__5507),
            .I(N__5504));
    Odrv4 I__830 (
            .O(N__5504),
            .I(un1_D_UM_040_1));
    InMux I__829 (
            .O(N__5501),
            .I(N__5498));
    LocalMux I__828 (
            .O(N__5498),
            .I(N__5495));
    Span4Mux_v I__827 (
            .O(N__5495),
            .I(N__5492));
    Sp12to4 I__826 (
            .O(N__5492),
            .I(N__5489));
    Span12Mux_h I__825 (
            .O(N__5489),
            .I(N__5486));
    Odrv12 I__824 (
            .O(N__5486),
            .I(D_LM_AMIGA_in_6));
    IoInMux I__823 (
            .O(N__5483),
            .I(N__5480));
    LocalMux I__822 (
            .O(N__5480),
            .I(N__5477));
    IoSpan4Mux I__821 (
            .O(N__5477),
            .I(N__5474));
    Sp12to4 I__820 (
            .O(N__5474),
            .I(N__5471));
    Span12Mux_s9_h I__819 (
            .O(N__5471),
            .I(N__5468));
    Odrv12 I__818 (
            .O(N__5468),
            .I(un2_D_LM_AMIGA_6));
    IoInMux I__817 (
            .O(N__5465),
            .I(N__5462));
    LocalMux I__816 (
            .O(N__5462),
            .I(N__5459));
    Span4Mux_s3_h I__815 (
            .O(N__5459),
            .I(N__5456));
    Span4Mux_h I__814 (
            .O(N__5456),
            .I(N__5452));
    InMux I__813 (
            .O(N__5455),
            .I(N__5449));
    Span4Mux_h I__812 (
            .O(N__5452),
            .I(N__5446));
    LocalMux I__811 (
            .O(N__5449),
            .I(N__5443));
    Sp12to4 I__810 (
            .O(N__5446),
            .I(N__5438));
    Span12Mux_v I__809 (
            .O(N__5443),
            .I(N__5438));
    Span12Mux_v I__808 (
            .O(N__5438),
            .I(N__5435));
    Span12Mux_h I__807 (
            .O(N__5435),
            .I(N__5432));
    Odrv12 I__806 (
            .O(N__5432),
            .I(D_LM_040_in_1));
    InMux I__805 (
            .O(N__5429),
            .I(N__5426));
    LocalMux I__804 (
            .O(N__5426),
            .I(N__5423));
    Span12Mux_v I__803 (
            .O(N__5423),
            .I(N__5420));
    Span12Mux_h I__802 (
            .O(N__5420),
            .I(N__5417));
    Odrv12 I__801 (
            .O(N__5417),
            .I(D_UU_040_in_1));
    IoInMux I__800 (
            .O(N__5414),
            .I(N__5411));
    LocalMux I__799 (
            .O(N__5411),
            .I(N__5408));
    Span4Mux_s3_h I__798 (
            .O(N__5408),
            .I(N__5405));
    Span4Mux_h I__797 (
            .O(N__5405),
            .I(N__5402));
    Span4Mux_h I__796 (
            .O(N__5402),
            .I(N__5399));
    Odrv4 I__795 (
            .O(N__5399),
            .I(un1_D_UU_040_1));
    IoInMux I__794 (
            .O(N__5396),
            .I(N__5392));
    InMux I__793 (
            .O(N__5395),
            .I(N__5389));
    LocalMux I__792 (
            .O(N__5392),
            .I(N__5386));
    LocalMux I__791 (
            .O(N__5389),
            .I(N__5383));
    IoSpan4Mux I__790 (
            .O(N__5386),
            .I(N__5380));
    Span4Mux_v I__789 (
            .O(N__5383),
            .I(N__5377));
    Span4Mux_s2_h I__788 (
            .O(N__5380),
            .I(N__5374));
    Sp12to4 I__787 (
            .O(N__5377),
            .I(N__5371));
    Span4Mux_v I__786 (
            .O(N__5374),
            .I(N__5368));
    Span12Mux_h I__785 (
            .O(N__5371),
            .I(N__5365));
    Sp12to4 I__784 (
            .O(N__5368),
            .I(N__5362));
    Span12Mux_v I__783 (
            .O(N__5365),
            .I(N__5359));
    Span12Mux_h I__782 (
            .O(N__5362),
            .I(N__5356));
    Span12Mux_v I__781 (
            .O(N__5359),
            .I(N__5353));
    Span12Mux_h I__780 (
            .O(N__5356),
            .I(N__5350));
    Odrv12 I__779 (
            .O(N__5353),
            .I(D_LL_040_in_5));
    Odrv12 I__778 (
            .O(N__5350),
            .I(D_LL_040_in_5));
    InMux I__777 (
            .O(N__5345),
            .I(N__5342));
    LocalMux I__776 (
            .O(N__5342),
            .I(N__5339));
    Span4Mux_v I__775 (
            .O(N__5339),
            .I(N__5336));
    Span4Mux_h I__774 (
            .O(N__5336),
            .I(N__5333));
    Sp12to4 I__773 (
            .O(N__5333),
            .I(N__5330));
    Span12Mux_h I__772 (
            .O(N__5330),
            .I(N__5327));
    Odrv12 I__771 (
            .O(N__5327),
            .I(D_UM_040_in_5));
    IoInMux I__770 (
            .O(N__5324),
            .I(N__5321));
    LocalMux I__769 (
            .O(N__5321),
            .I(N__5318));
    IoSpan4Mux I__768 (
            .O(N__5318),
            .I(N__5315));
    Span4Mux_s2_v I__767 (
            .O(N__5315),
            .I(N__5312));
    Span4Mux_h I__766 (
            .O(N__5312),
            .I(N__5309));
    Span4Mux_v I__765 (
            .O(N__5309),
            .I(N__5306));
    Odrv4 I__764 (
            .O(N__5306),
            .I(un1_D_UM_040_5));
    InMux I__763 (
            .O(N__5303),
            .I(N__5300));
    LocalMux I__762 (
            .O(N__5300),
            .I(WRITE_CYCLE_ACTIVE_rep13_i_ess));
    InMux I__761 (
            .O(N__5297),
            .I(N__5294));
    LocalMux I__760 (
            .O(N__5294),
            .I(WRITE_CYCLE_ACTIVE_rep4_i_ess));
    IoInMux I__759 (
            .O(N__5291),
            .I(N__5288));
    LocalMux I__758 (
            .O(N__5288),
            .I(N__5285));
    IoSpan4Mux I__757 (
            .O(N__5285),
            .I(N__5282));
    Span4Mux_s3_v I__756 (
            .O(N__5282),
            .I(N__5279));
    Odrv4 I__755 (
            .O(N__5279),
            .I(N_217_i));
    InMux I__754 (
            .O(N__5276),
            .I(N__5273));
    LocalMux I__753 (
            .O(N__5273),
            .I(N__5270));
    Span4Mux_v I__752 (
            .O(N__5270),
            .I(N__5267));
    Sp12to4 I__751 (
            .O(N__5267),
            .I(N__5264));
    Odrv12 I__750 (
            .O(N__5264),
            .I(D_LL_AMIGA_in_4));
    IoInMux I__749 (
            .O(N__5261),
            .I(N__5258));
    LocalMux I__748 (
            .O(N__5258),
            .I(N__5255));
    Span4Mux_s2_h I__747 (
            .O(N__5255),
            .I(N__5252));
    Sp12to4 I__746 (
            .O(N__5252),
            .I(N__5249));
    Span12Mux_s8_v I__745 (
            .O(N__5249),
            .I(N__5246));
    Span12Mux_h I__744 (
            .O(N__5246),
            .I(N__5243));
    Odrv12 I__743 (
            .O(N__5243),
            .I(un2_D_LL_AMIGA_4));
    IoInMux I__742 (
            .O(N__5240),
            .I(N__5236));
    InMux I__741 (
            .O(N__5239),
            .I(N__5233));
    LocalMux I__740 (
            .O(N__5236),
            .I(N__5230));
    LocalMux I__739 (
            .O(N__5233),
            .I(N__5227));
    IoSpan4Mux I__738 (
            .O(N__5230),
            .I(N__5224));
    Span4Mux_v I__737 (
            .O(N__5227),
            .I(N__5221));
    Span4Mux_s2_h I__736 (
            .O(N__5224),
            .I(N__5218));
    Sp12to4 I__735 (
            .O(N__5221),
            .I(N__5215));
    Sp12to4 I__734 (
            .O(N__5218),
            .I(N__5212));
    Span12Mux_h I__733 (
            .O(N__5215),
            .I(N__5209));
    Span12Mux_h I__732 (
            .O(N__5212),
            .I(N__5206));
    Span12Mux_v I__731 (
            .O(N__5209),
            .I(N__5203));
    Span12Mux_h I__730 (
            .O(N__5206),
            .I(N__5200));
    Odrv12 I__729 (
            .O(N__5203),
            .I(D_LL_040_in_0));
    Odrv12 I__728 (
            .O(N__5200),
            .I(D_LL_040_in_0));
    InMux I__727 (
            .O(N__5195),
            .I(N__5192));
    LocalMux I__726 (
            .O(N__5192),
            .I(N__5189));
    Span12Mux_h I__725 (
            .O(N__5189),
            .I(N__5186));
    Span12Mux_h I__724 (
            .O(N__5186),
            .I(N__5183));
    Odrv12 I__723 (
            .O(N__5183),
            .I(D_UM_040_in_0));
    IoInMux I__722 (
            .O(N__5180),
            .I(N__5177));
    LocalMux I__721 (
            .O(N__5177),
            .I(N__5174));
    IoSpan4Mux I__720 (
            .O(N__5174),
            .I(N__5171));
    Span4Mux_s1_h I__719 (
            .O(N__5171),
            .I(N__5168));
    Span4Mux_h I__718 (
            .O(N__5168),
            .I(N__5165));
    Span4Mux_h I__717 (
            .O(N__5165),
            .I(N__5162));
    Odrv4 I__716 (
            .O(N__5162),
            .I(un1_D_UM_040_0));
    InMux I__715 (
            .O(N__5159),
            .I(N__5156));
    LocalMux I__714 (
            .O(N__5156),
            .I(N__5153));
    Span12Mux_h I__713 (
            .O(N__5153),
            .I(N__5150));
    Odrv12 I__712 (
            .O(N__5150),
            .I(D_LM_AMIGA_in_3));
    IoInMux I__711 (
            .O(N__5147),
            .I(N__5144));
    LocalMux I__710 (
            .O(N__5144),
            .I(N__5141));
    IoSpan4Mux I__709 (
            .O(N__5141),
            .I(N__5138));
    Span4Mux_s0_h I__708 (
            .O(N__5138),
            .I(N__5135));
    Sp12to4 I__707 (
            .O(N__5135),
            .I(N__5132));
    Span12Mux_s9_h I__706 (
            .O(N__5132),
            .I(N__5129));
    Span12Mux_h I__705 (
            .O(N__5129),
            .I(N__5126));
    Odrv12 I__704 (
            .O(N__5126),
            .I(un2_D_LM_AMIGA_3));
    IoInMux I__703 (
            .O(N__5123),
            .I(N__5120));
    LocalMux I__702 (
            .O(N__5120),
            .I(N__5117));
    IoSpan4Mux I__701 (
            .O(N__5117),
            .I(N__5114));
    Span4Mux_s2_v I__700 (
            .O(N__5114),
            .I(N__5111));
    Span4Mux_v I__699 (
            .O(N__5111),
            .I(N__5108));
    Odrv4 I__698 (
            .O(N__5108),
            .I(LBENn_c_i));
    InMux I__697 (
            .O(N__5105),
            .I(N__5102));
    LocalMux I__696 (
            .O(N__5102),
            .I(WRITE_CYCLE_ACTIVE_rep2_i_ess));
    IoInMux I__695 (
            .O(N__5099),
            .I(N__5096));
    LocalMux I__694 (
            .O(N__5096),
            .I(N__5093));
    Span4Mux_s2_v I__693 (
            .O(N__5093),
            .I(N__5090));
    Span4Mux_h I__692 (
            .O(N__5090),
            .I(N__5087));
    Span4Mux_v I__691 (
            .O(N__5087),
            .I(N__5084));
    Odrv4 I__690 (
            .O(N__5084),
            .I(N_215_i));
    InMux I__689 (
            .O(N__5081),
            .I(N__5078));
    LocalMux I__688 (
            .O(N__5078),
            .I(N__5075));
    Span4Mux_v I__687 (
            .O(N__5075),
            .I(N__5072));
    Sp12to4 I__686 (
            .O(N__5072),
            .I(N__5069));
    Span12Mux_h I__685 (
            .O(N__5069),
            .I(N__5066));
    Odrv12 I__684 (
            .O(N__5066),
            .I(D_UM_040_in_6));
    IoInMux I__683 (
            .O(N__5063),
            .I(N__5060));
    LocalMux I__682 (
            .O(N__5060),
            .I(N__5057));
    IoSpan4Mux I__681 (
            .O(N__5057),
            .I(N__5054));
    Span4Mux_s1_h I__680 (
            .O(N__5054),
            .I(N__5050));
    InMux I__679 (
            .O(N__5053),
            .I(N__5047));
    Span4Mux_h I__678 (
            .O(N__5050),
            .I(N__5044));
    LocalMux I__677 (
            .O(N__5047),
            .I(N__5041));
    Span4Mux_h I__676 (
            .O(N__5044),
            .I(N__5036));
    Span4Mux_v I__675 (
            .O(N__5041),
            .I(N__5036));
    Sp12to4 I__674 (
            .O(N__5036),
            .I(N__5033));
    Span12Mux_v I__673 (
            .O(N__5033),
            .I(N__5030));
    Span12Mux_h I__672 (
            .O(N__5030),
            .I(N__5027));
    Odrv12 I__671 (
            .O(N__5027),
            .I(D_LL_040_in_6));
    IoInMux I__670 (
            .O(N__5024),
            .I(N__5021));
    LocalMux I__669 (
            .O(N__5021),
            .I(N__5018));
    Span12Mux_s2_h I__668 (
            .O(N__5018),
            .I(N__5015));
    Span12Mux_v I__667 (
            .O(N__5015),
            .I(N__5012));
    Odrv12 I__666 (
            .O(N__5012),
            .I(un1_D_UM_040_6));
    InMux I__665 (
            .O(N__5009),
            .I(N__5006));
    LocalMux I__664 (
            .O(N__5006),
            .I(N__5003));
    Odrv12 I__663 (
            .O(N__5003),
            .I(D_LM_AMIGA_in_2));
    IoInMux I__662 (
            .O(N__5000),
            .I(N__4997));
    LocalMux I__661 (
            .O(N__4997),
            .I(N__4994));
    Sp12to4 I__660 (
            .O(N__4994),
            .I(N__4991));
    Span12Mux_h I__659 (
            .O(N__4991),
            .I(N__4988));
    Span12Mux_v I__658 (
            .O(N__4988),
            .I(N__4985));
    Odrv12 I__657 (
            .O(N__4985),
            .I(un2_D_LM_AMIGA_2));
    InMux I__656 (
            .O(N__4982),
            .I(N__4979));
    LocalMux I__655 (
            .O(N__4979),
            .I(WRITE_CYCLE_ACTIVE_rep0_i_ess));
    IoInMux I__654 (
            .O(N__4976),
            .I(N__4973));
    LocalMux I__653 (
            .O(N__4973),
            .I(N__4970));
    Span4Mux_s3_v I__652 (
            .O(N__4970),
            .I(N__4967));
    Span4Mux_v I__651 (
            .O(N__4967),
            .I(N__4964));
    Odrv4 I__650 (
            .O(N__4964),
            .I(N_213_i));
    IoInMux I__649 (
            .O(N__4961),
            .I(N__4958));
    LocalMux I__648 (
            .O(N__4958),
            .I(N__4955));
    Span4Mux_s3_v I__647 (
            .O(N__4955),
            .I(N__4952));
    Span4Mux_h I__646 (
            .O(N__4952),
            .I(N__4949));
    Span4Mux_v I__645 (
            .O(N__4949),
            .I(N__4946));
    Odrv4 I__644 (
            .O(N__4946),
            .I(N_226_i));
    InMux I__643 (
            .O(N__4943),
            .I(N__4940));
    LocalMux I__642 (
            .O(N__4940),
            .I(N__4937));
    Odrv4 I__641 (
            .O(N__4937),
            .I(WRITE_CYCLE_ACTIVE_rep6_i_ess));
    InMux I__640 (
            .O(N__4934),
            .I(N__4931));
    LocalMux I__639 (
            .O(N__4931),
            .I(N__4928));
    Span12Mux_v I__638 (
            .O(N__4928),
            .I(N__4925));
    Odrv12 I__637 (
            .O(N__4925),
            .I(D_LL_AMIGA_in_1));
    IoInMux I__636 (
            .O(N__4922),
            .I(N__4919));
    LocalMux I__635 (
            .O(N__4919),
            .I(N__4916));
    Span4Mux_s3_h I__634 (
            .O(N__4916),
            .I(N__4913));
    Sp12to4 I__633 (
            .O(N__4913),
            .I(N__4910));
    Span12Mux_s8_v I__632 (
            .O(N__4910),
            .I(N__4907));
    Span12Mux_h I__631 (
            .O(N__4907),
            .I(N__4904));
    Odrv12 I__630 (
            .O(N__4904),
            .I(un2_D_LL_AMIGA_1));
    InMux I__629 (
            .O(N__4901),
            .I(N__4898));
    LocalMux I__628 (
            .O(N__4898),
            .I(N__4895));
    Span4Mux_v I__627 (
            .O(N__4895),
            .I(N__4892));
    Span4Mux_v I__626 (
            .O(N__4892),
            .I(N__4888));
    InMux I__625 (
            .O(N__4891),
            .I(N__4885));
    Sp12to4 I__624 (
            .O(N__4888),
            .I(N__4880));
    LocalMux I__623 (
            .O(N__4885),
            .I(N__4880));
    Span12Mux_h I__622 (
            .O(N__4880),
            .I(N__4877));
    Odrv12 I__621 (
            .O(N__4877),
            .I(A_040_c_1));
    InMux I__620 (
            .O(N__4874),
            .I(N__4871));
    LocalMux I__619 (
            .O(N__4871),
            .I(N__4868));
    Odrv4 I__618 (
            .O(N__4868),
            .I(WRITE_CYCLE_ACTIVE_rep21_i_ess));
    InMux I__617 (
            .O(N__4865),
            .I(N__4862));
    LocalMux I__616 (
            .O(N__4862),
            .I(N__4859));
    Span4Mux_v I__615 (
            .O(N__4859),
            .I(N__4856));
    Odrv4 I__614 (
            .O(N__4856),
            .I(WRITE_CYCLE_ACTIVE_rep23_i_ess));
    InMux I__613 (
            .O(N__4853),
            .I(N__4850));
    LocalMux I__612 (
            .O(N__4850),
            .I(WRITE_CYCLE_ACTIVE_rep7_i_ess));
    IoInMux I__611 (
            .O(N__4847),
            .I(N__4844));
    LocalMux I__610 (
            .O(N__4844),
            .I(N__4841));
    IoSpan4Mux I__609 (
            .O(N__4841),
            .I(N__4838));
    Span4Mux_s2_v I__608 (
            .O(N__4838),
            .I(N__4835));
    Span4Mux_v I__607 (
            .O(N__4835),
            .I(N__4832));
    Odrv4 I__606 (
            .O(N__4832),
            .I(N_220_i));
    InMux I__605 (
            .O(N__4829),
            .I(N__4826));
    LocalMux I__604 (
            .O(N__4826),
            .I(WRITE_CYCLE_ACTIVE_rep3_i_ess));
    IoInMux I__603 (
            .O(N__4823),
            .I(N__4820));
    LocalMux I__602 (
            .O(N__4820),
            .I(N__4817));
    IoSpan4Mux I__601 (
            .O(N__4817),
            .I(N__4814));
    Span4Mux_s3_v I__600 (
            .O(N__4814),
            .I(N__4811));
    Odrv4 I__599 (
            .O(N__4811),
            .I(N_219_i));
    InMux I__598 (
            .O(N__4808),
            .I(N__4805));
    LocalMux I__597 (
            .O(N__4805),
            .I(N__4802));
    Span4Mux_v I__596 (
            .O(N__4802),
            .I(N__4799));
    Sp12to4 I__595 (
            .O(N__4799),
            .I(N__4796));
    Odrv12 I__594 (
            .O(N__4796),
            .I(D_LL_AMIGA_in_0));
    IoInMux I__593 (
            .O(N__4793),
            .I(N__4790));
    LocalMux I__592 (
            .O(N__4790),
            .I(N__4787));
    Span12Mux_s11_h I__591 (
            .O(N__4787),
            .I(N__4784));
    Span12Mux_h I__590 (
            .O(N__4784),
            .I(N__4781));
    Odrv12 I__589 (
            .O(N__4781),
            .I(un2_D_LL_AMIGA_0));
    InMux I__588 (
            .O(N__4778),
            .I(N__4775));
    LocalMux I__587 (
            .O(N__4775),
            .I(N__4772));
    Odrv12 I__586 (
            .O(N__4772),
            .I(D_LM_AMIGA_in_1));
    IoInMux I__585 (
            .O(N__4769),
            .I(N__4766));
    LocalMux I__584 (
            .O(N__4766),
            .I(N__4763));
    Span4Mux_s3_h I__583 (
            .O(N__4763),
            .I(N__4760));
    Span4Mux_h I__582 (
            .O(N__4760),
            .I(N__4757));
    Sp12to4 I__581 (
            .O(N__4757),
            .I(N__4754));
    Span12Mux_v I__580 (
            .O(N__4754),
            .I(N__4751));
    Span12Mux_h I__579 (
            .O(N__4751),
            .I(N__4748));
    Odrv12 I__578 (
            .O(N__4748),
            .I(un2_D_LM_AMIGA_1));
    InMux I__577 (
            .O(N__4745),
            .I(N__4742));
    LocalMux I__576 (
            .O(N__4742),
            .I(N__4739));
    Span12Mux_h I__575 (
            .O(N__4739),
            .I(N__4736));
    Span12Mux_h I__574 (
            .O(N__4736),
            .I(N__4733));
    Odrv12 I__573 (
            .O(N__4733),
            .I(D_UM_040_in_2));
    IoInMux I__572 (
            .O(N__4730),
            .I(N__4726));
    InMux I__571 (
            .O(N__4729),
            .I(N__4723));
    LocalMux I__570 (
            .O(N__4726),
            .I(N__4720));
    LocalMux I__569 (
            .O(N__4723),
            .I(N__4717));
    IoSpan4Mux I__568 (
            .O(N__4720),
            .I(N__4714));
    Span4Mux_v I__567 (
            .O(N__4717),
            .I(N__4711));
    Span4Mux_s2_h I__566 (
            .O(N__4714),
            .I(N__4708));
    Sp12to4 I__565 (
            .O(N__4711),
            .I(N__4705));
    Sp12to4 I__564 (
            .O(N__4708),
            .I(N__4702));
    Span12Mux_v I__563 (
            .O(N__4705),
            .I(N__4699));
    Span12Mux_h I__562 (
            .O(N__4702),
            .I(N__4696));
    Span12Mux_h I__561 (
            .O(N__4699),
            .I(N__4693));
    Span12Mux_h I__560 (
            .O(N__4696),
            .I(N__4690));
    Odrv12 I__559 (
            .O(N__4693),
            .I(D_LL_040_in_2));
    Odrv12 I__558 (
            .O(N__4690),
            .I(D_LL_040_in_2));
    IoInMux I__557 (
            .O(N__4685),
            .I(N__4682));
    LocalMux I__556 (
            .O(N__4682),
            .I(N__4679));
    Span4Mux_s3_h I__555 (
            .O(N__4679),
            .I(N__4676));
    Span4Mux_h I__554 (
            .O(N__4676),
            .I(N__4673));
    Span4Mux_v I__553 (
            .O(N__4673),
            .I(N__4670));
    Odrv4 I__552 (
            .O(N__4670),
            .I(un1_D_UM_040_2));
    IoInMux I__551 (
            .O(N__4667),
            .I(N__4664));
    LocalMux I__550 (
            .O(N__4664),
            .I(N__4661));
    Span4Mux_s3_v I__549 (
            .O(N__4661),
            .I(N__4658));
    Span4Mux_h I__548 (
            .O(N__4658),
            .I(N__4655));
    Odrv4 I__547 (
            .O(N__4655),
            .I(N_216_i));
    InMux I__546 (
            .O(N__4652),
            .I(N__4649));
    LocalMux I__545 (
            .O(N__4649),
            .I(N__4646));
    Odrv12 I__544 (
            .O(N__4646),
            .I(WRITE_CYCLE_ACTIVE_rep5_i_ess));
    IoInMux I__543 (
            .O(N__4643),
            .I(N__4640));
    LocalMux I__542 (
            .O(N__4640),
            .I(N__4637));
    Span4Mux_s3_h I__541 (
            .O(N__4637),
            .I(N__4634));
    Span4Mux_v I__540 (
            .O(N__4634),
            .I(N__4631));
    Odrv4 I__539 (
            .O(N__4631),
            .I(N_218_i));
    InMux I__538 (
            .O(N__4628),
            .I(N__4625));
    LocalMux I__537 (
            .O(N__4625),
            .I(N__4622));
    Span4Mux_h I__536 (
            .O(N__4622),
            .I(N__4619));
    Span4Mux_v I__535 (
            .O(N__4619),
            .I(N__4616));
    Odrv4 I__534 (
            .O(N__4616),
            .I(A_040_c_0));
    IoInMux I__533 (
            .O(N__4613),
            .I(N__4610));
    LocalMux I__532 (
            .O(N__4610),
            .I(N__4607));
    Span4Mux_s2_v I__531 (
            .O(N__4607),
            .I(N__4604));
    Span4Mux_v I__530 (
            .O(N__4604),
            .I(N__4601));
    Odrv4 I__529 (
            .O(N__4601),
            .I(A_AMIGA_c_0));
    IoInMux I__528 (
            .O(N__4598),
            .I(N__4595));
    LocalMux I__527 (
            .O(N__4595),
            .I(N__4592));
    Odrv12 I__526 (
            .O(N__4592),
            .I(U111_CYCLE_SM_A_AMIGA_0_i_1));
    InMux I__525 (
            .O(N__4589),
            .I(N__4586));
    LocalMux I__524 (
            .O(N__4586),
            .I(WRITE_CYCLE_ACTIVE_rep28_i_ess));
    InMux I__523 (
            .O(N__4583),
            .I(N__4580));
    LocalMux I__522 (
            .O(N__4580),
            .I(N__4577));
    Span4Mux_v I__521 (
            .O(N__4577),
            .I(N__4574));
    Odrv4 I__520 (
            .O(N__4574),
            .I(WRITE_CYCLE_ACTIVE_rep27_i_ess));
    InMux I__519 (
            .O(N__4571),
            .I(N__4568));
    LocalMux I__518 (
            .O(N__4568),
            .I(WRITE_CYCLE_ACTIVE_rep19_i_ess));
    IoInMux I__517 (
            .O(N__4565),
            .I(N__4562));
    LocalMux I__516 (
            .O(N__4562),
            .I(N__4559));
    Odrv12 I__515 (
            .O(N__4559),
            .I(N_231_i));
    InMux I__514 (
            .O(N__4556),
            .I(N__4553));
    LocalMux I__513 (
            .O(N__4553),
            .I(WRITE_CYCLE_ACTIVE_rep18_i_ess));
    IoInMux I__512 (
            .O(N__4550),
            .I(N__4547));
    LocalMux I__511 (
            .O(N__4547),
            .I(N__4544));
    Odrv12 I__510 (
            .O(N__4544),
            .I(N_232_i));
    InMux I__509 (
            .O(N__4541),
            .I(N__4538));
    LocalMux I__508 (
            .O(N__4538),
            .I(WRITE_CYCLE_ACTIVE_rep8_i_ess));
    InMux I__507 (
            .O(N__4535),
            .I(N__4532));
    LocalMux I__506 (
            .O(N__4532),
            .I(WRITE_CYCLE_ACTIVE_rep20_i_ess));
    InMux I__505 (
            .O(N__4529),
            .I(N__4526));
    LocalMux I__504 (
            .O(N__4526),
            .I(WRITE_CYCLE_ACTIVE_rep11_i_ess));
    InMux I__503 (
            .O(N__4523),
            .I(N__4520));
    LocalMux I__502 (
            .O(N__4520),
            .I(WRITE_CYCLE_ACTIVE_rep22_i_ess));
    InMux I__501 (
            .O(N__4517),
            .I(N__4514));
    LocalMux I__500 (
            .O(N__4514),
            .I(WRITE_CYCLE_ACTIVE_rep14_i_ess));
    InMux I__499 (
            .O(N__4511),
            .I(N__4508));
    LocalMux I__498 (
            .O(N__4508),
            .I(WRITE_CYCLE_ACTIVE_rep1_i_ess));
    InMux I__497 (
            .O(N__4505),
            .I(N__4502));
    LocalMux I__496 (
            .O(N__4502),
            .I(WRITE_CYCLE_ACTIVE_rep12_i_ess));
    IoInMux I__495 (
            .O(N__4499),
            .I(N__4496));
    LocalMux I__494 (
            .O(N__4496),
            .I(N__4493));
    IoSpan4Mux I__493 (
            .O(N__4493),
            .I(N__4490));
    Span4Mux_s2_h I__492 (
            .O(N__4490),
            .I(N__4487));
    Odrv4 I__491 (
            .O(N__4487),
            .I(N_214_i));
    IoInMux I__490 (
            .O(N__4484),
            .I(N__4481));
    LocalMux I__489 (
            .O(N__4481),
            .I(N__4478));
    IoSpan4Mux I__488 (
            .O(N__4478),
            .I(N__4475));
    Span4Mux_s3_h I__487 (
            .O(N__4475),
            .I(N__4472));
    Odrv4 I__486 (
            .O(N__4472),
            .I(N_228_i));
    IoInMux I__485 (
            .O(N__4469),
            .I(N__4466));
    LocalMux I__484 (
            .O(N__4466),
            .I(N__4463));
    IoSpan4Mux I__483 (
            .O(N__4463),
            .I(N__4460));
    Span4Mux_s2_h I__482 (
            .O(N__4460),
            .I(N__4457));
    Odrv4 I__481 (
            .O(N__4457),
            .I(N_225_i));
    InMux I__480 (
            .O(N__4454),
            .I(N__4451));
    LocalMux I__479 (
            .O(N__4451),
            .I(WRITE_CYCLE_ACTIVE_rep15_i_ess));
    IoInMux I__478 (
            .O(N__4448),
            .I(N__4445));
    LocalMux I__477 (
            .O(N__4445),
            .I(N__4442));
    IoSpan4Mux I__476 (
            .O(N__4442),
            .I(N__4439));
    Span4Mux_s1_h I__475 (
            .O(N__4439),
            .I(N__4436));
    Span4Mux_h I__474 (
            .O(N__4436),
            .I(N__4433));
    Odrv4 I__473 (
            .O(N__4433),
            .I(N_241_i));
    InMux I__472 (
            .O(N__4430),
            .I(N__4427));
    LocalMux I__471 (
            .O(N__4427),
            .I(WRITE_CYCLE_ACTIVE_rep25_i_ess));
    InMux I__470 (
            .O(N__4424),
            .I(N__4421));
    LocalMux I__469 (
            .O(N__4421),
            .I(WRITE_CYCLE_ACTIVE_rep30_i_ess));
    InMux I__468 (
            .O(N__4418),
            .I(N__4415));
    LocalMux I__467 (
            .O(N__4415),
            .I(WRITE_CYCLE_ACTIVE_i_ess));
    InMux I__466 (
            .O(N__4412),
            .I(N__4409));
    LocalMux I__465 (
            .O(N__4409),
            .I(WRITE_CYCLE_ACTIVE_rep16_i_ess));
    IoInMux I__464 (
            .O(N__4406),
            .I(N__4403));
    LocalMux I__463 (
            .O(N__4403),
            .I(N__4400));
    Span12Mux_s4_h I__462 (
            .O(N__4400),
            .I(N__4397));
    Odrv12 I__461 (
            .O(N__4397),
            .I(N_223_i));
    IoInMux I__460 (
            .O(N__4394),
            .I(N__4391));
    LocalMux I__459 (
            .O(N__4391),
            .I(N__4388));
    IoSpan4Mux I__458 (
            .O(N__4388),
            .I(N__4385));
    Span4Mux_s3_h I__457 (
            .O(N__4385),
            .I(N__4382));
    Odrv4 I__456 (
            .O(N__4382),
            .I(N_233_i));
    InMux I__455 (
            .O(N__4379),
            .I(N__4376));
    LocalMux I__454 (
            .O(N__4376),
            .I(WRITE_CYCLE_ACTIVE_rep10_i_ess));
    IoInMux I__453 (
            .O(N__4373),
            .I(N__4370));
    LocalMux I__452 (
            .O(N__4370),
            .I(N__4367));
    Span12Mux_s4_h I__451 (
            .O(N__4367),
            .I(N__4364));
    Odrv12 I__450 (
            .O(N__4364),
            .I(N_234_i));
    InMux I__449 (
            .O(N__4361),
            .I(N__4358));
    LocalMux I__448 (
            .O(N__4358),
            .I(WRITE_CYCLE_ACTIVE_rep9_i_ess));
    IoInMux I__447 (
            .O(N__4355),
            .I(N__4352));
    LocalMux I__446 (
            .O(N__4352),
            .I(N__4349));
    IoSpan4Mux I__445 (
            .O(N__4349),
            .I(N__4346));
    Span4Mux_s3_h I__444 (
            .O(N__4346),
            .I(N__4343));
    Odrv4 I__443 (
            .O(N__4343),
            .I(N_222_i));
    IoInMux I__442 (
            .O(N__4340),
            .I(N__4337));
    LocalMux I__441 (
            .O(N__4337),
            .I(N__4334));
    IoSpan4Mux I__440 (
            .O(N__4334),
            .I(N__4331));
    Span4Mux_s3_h I__439 (
            .O(N__4331),
            .I(N__4328));
    Odrv4 I__438 (
            .O(N__4328),
            .I(N_236_i));
    IoInMux I__437 (
            .O(N__4325),
            .I(N__4322));
    LocalMux I__436 (
            .O(N__4322),
            .I(N__4319));
    Span4Mux_s0_h I__435 (
            .O(N__4319),
            .I(N__4316));
    Span4Mux_h I__434 (
            .O(N__4316),
            .I(N__4313));
    Odrv4 I__433 (
            .O(N__4313),
            .I(N_235_i));
    IoInMux I__432 (
            .O(N__4310),
            .I(N__4307));
    LocalMux I__431 (
            .O(N__4307),
            .I(N__4304));
    Span4Mux_s3_h I__430 (
            .O(N__4304),
            .I(N__4301));
    Span4Mux_v I__429 (
            .O(N__4301),
            .I(N__4298));
    Odrv4 I__428 (
            .O(N__4298),
            .I(N_224_i));
    IoInMux I__427 (
            .O(N__4295),
            .I(N__4292));
    LocalMux I__426 (
            .O(N__4292),
            .I(N__4289));
    Span12Mux_s4_h I__425 (
            .O(N__4289),
            .I(N__4286));
    Odrv12 I__424 (
            .O(N__4286),
            .I(N_227_i));
    IoInMux I__423 (
            .O(N__4283),
            .I(N__4280));
    LocalMux I__422 (
            .O(N__4280),
            .I(N__4277));
    Span4Mux_s0_h I__421 (
            .O(N__4277),
            .I(N__4274));
    Span4Mux_h I__420 (
            .O(N__4274),
            .I(N__4271));
    Odrv4 I__419 (
            .O(N__4271),
            .I(N_243_i));
    IoInMux I__418 (
            .O(N__4268),
            .I(N__4265));
    LocalMux I__417 (
            .O(N__4265),
            .I(N__4262));
    Span12Mux_s4_h I__416 (
            .O(N__4262),
            .I(N__4259));
    Odrv12 I__415 (
            .O(N__4259),
            .I(N_229_i));
    IoInMux I__414 (
            .O(N__4256),
            .I(N__4253));
    LocalMux I__413 (
            .O(N__4253),
            .I(N__4250));
    Span4Mux_s0_h I__412 (
            .O(N__4250),
            .I(N__4247));
    Span4Mux_h I__411 (
            .O(N__4247),
            .I(N__4244));
    Odrv4 I__410 (
            .O(N__4244),
            .I(N_244_i));
    InMux I__409 (
            .O(N__4241),
            .I(N__4238));
    LocalMux I__408 (
            .O(N__4238),
            .I(N__4235));
    Odrv4 I__407 (
            .O(N__4235),
            .I(WRITE_CYCLE_ACTIVE_rep29_i_ess));
    InMux I__406 (
            .O(N__4232),
            .I(N__4229));
    LocalMux I__405 (
            .O(N__4229),
            .I(WRITE_CYCLE_ACTIVE_rep17_i_ess));
    IoInMux I__404 (
            .O(N__4226),
            .I(N__4223));
    LocalMux I__403 (
            .O(N__4223),
            .I(N__4220));
    IoSpan4Mux I__402 (
            .O(N__4220),
            .I(N__4217));
    Span4Mux_s3_h I__401 (
            .O(N__4217),
            .I(N__4214));
    Odrv4 I__400 (
            .O(N__4214),
            .I(N_230_i));
    IoInMux I__399 (
            .O(N__4211),
            .I(N__4208));
    LocalMux I__398 (
            .O(N__4208),
            .I(N__4205));
    Odrv12 I__397 (
            .O(N__4205),
            .I(RESETn_c_i));
    IoInMux I__396 (
            .O(N__4202),
            .I(N__4199));
    LocalMux I__395 (
            .O(N__4199),
            .I(N__4196));
    IoSpan4Mux I__394 (
            .O(N__4196),
            .I(N__4193));
    Span4Mux_s1_h I__393 (
            .O(N__4193),
            .I(N__4190));
    Odrv4 I__392 (
            .O(N__4190),
            .I(\U111_CYCLE_SM.CYCLE_STATE_0_0 ));
    IoInMux I__391 (
            .O(N__4187),
            .I(N__4184));
    LocalMux I__390 (
            .O(N__4184),
            .I(N__4181));
    Odrv12 I__389 (
            .O(N__4181),
            .I(N_221_i));
    IoInMux I__388 (
            .O(N__4178),
            .I(N__4175));
    LocalMux I__387 (
            .O(N__4175),
            .I(N__4172));
    Span4Mux_s0_v I__386 (
            .O(N__4172),
            .I(N__4169));
    Sp12to4 I__385 (
            .O(N__4169),
            .I(N__4166));
    Span12Mux_h I__384 (
            .O(N__4166),
            .I(N__4163));
    Span12Mux_v I__383 (
            .O(N__4163),
            .I(N__4160));
    Span12Mux_v I__382 (
            .O(N__4160),
            .I(N__4157));
    Odrv12 I__381 (
            .O(N__4157),
            .I(TAn_in));
    IoInMux I__380 (
            .O(N__4154),
            .I(N__4151));
    LocalMux I__379 (
            .O(N__4151),
            .I(N__4148));
    IoSpan4Mux I__378 (
            .O(N__4148),
            .I(N__4145));
    Span4Mux_s3_h I__377 (
            .O(N__4145),
            .I(N__4142));
    Odrv4 I__376 (
            .O(N__4142),
            .I(N_240_i));
    IoInMux I__375 (
            .O(N__4139),
            .I(N__4136));
    LocalMux I__374 (
            .O(N__4136),
            .I(N__4133));
    Span4Mux_s3_h I__373 (
            .O(N__4133),
            .I(N__4130));
    Span4Mux_v I__372 (
            .O(N__4130),
            .I(N__4127));
    Odrv4 I__371 (
            .O(N__4127),
            .I(N_237_i));
    IoInMux I__370 (
            .O(N__4124),
            .I(N__4121));
    LocalMux I__369 (
            .O(N__4121),
            .I(N__4118));
    IoSpan4Mux I__368 (
            .O(N__4118),
            .I(N__4115));
    Span4Mux_s2_h I__367 (
            .O(N__4115),
            .I(N__4112));
    Odrv4 I__366 (
            .O(N__4112),
            .I(N_239_i));
    InMux I__365 (
            .O(N__4109),
            .I(N__4106));
    LocalMux I__364 (
            .O(N__4106),
            .I(WRITE_CYCLE_ACTIVE_rep26_i_ess));
    IoInMux I__363 (
            .O(N__4103),
            .I(N__4100));
    LocalMux I__362 (
            .O(N__4100),
            .I(N__4097));
    Span4Mux_s3_h I__361 (
            .O(N__4097),
            .I(N__4094));
    Span4Mux_v I__360 (
            .O(N__4094),
            .I(N__4091));
    Odrv4 I__359 (
            .O(N__4091),
            .I(N_238_i));
    InMux I__358 (
            .O(N__4088),
            .I(N__4085));
    LocalMux I__357 (
            .O(N__4085),
            .I(N__4082));
    Odrv4 I__356 (
            .O(N__4082),
            .I(WRITE_CYCLE_ACTIVE_rep24_i_ess));
    IoInMux I__355 (
            .O(N__4079),
            .I(N__4076));
    LocalMux I__354 (
            .O(N__4076),
            .I(N__4073));
    Span4Mux_s0_h I__353 (
            .O(N__4073),
            .I(N__4070));
    Span4Mux_h I__352 (
            .O(N__4070),
            .I(N__4067));
    Odrv4 I__351 (
            .O(N__4067),
            .I(N_242_i));
    IoInMux I__350 (
            .O(N__4064),
            .I(N__4061));
    LocalMux I__349 (
            .O(N__4061),
            .I(N__4058));
    IoSpan4Mux I__348 (
            .O(N__4058),
            .I(N__4055));
    Span4Mux_s3_h I__347 (
            .O(N__4055),
            .I(N__4052));
    Sp12to4 I__346 (
            .O(N__4052),
            .I(N__4049));
    Span12Mux_s8_h I__345 (
            .O(N__4049),
            .I(N__4046));
    Span12Mux_v I__344 (
            .O(N__4046),
            .I(N__4043));
    Span12Mux_v I__343 (
            .O(N__4043),
            .I(N__4040));
    Span12Mux_h I__342 (
            .O(N__4040),
            .I(N__4037));
    Odrv12 I__341 (
            .O(N__4037),
            .I(TCIn_c));
    INV \INVU111_CYCLE_SM.TSnC  (
            .O(\INVU111_CYCLE_SM.TSnC_net ),
            .I(N__12817));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__4211),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    ICE_GB \U111_CYCLE_SM.CYCLE_STATE_RNIICIM_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__4202),
            .GLOBALBUFFEROUTPUT(\U111_CYCLE_SM.CYCLE_STATE_0_g_0 ));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam D_LL_AMIGA_iobuf_RNO_3_LC_1_2_3.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_3_LC_1_2_3.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_3_LC_1_2_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_3_LC_1_2_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4583),
            .lcout(N_240_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_AMIGA_iobuf_RNO_0_LC_1_2_6.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_0_LC_1_2_6.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_0_LC_1_2_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_0_LC_1_2_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4088),
            .lcout(N_237_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_AMIGA_iobuf_RNO_2_LC_1_2_7.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_2_LC_1_2_7.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_2_LC_1_2_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_2_LC_1_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4109),
            .lcout(N_239_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep26_i_ess_LC_1_3_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep26_i_ess_LC_1_3_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep26_i_ess_LC_1_3_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep26_i_ess_LC_1_3_5  (
            .in0(N__10382),
            .in1(N__11764),
            .in2(N__12216),
            .in3(N__10703),
            .lcout(WRITE_CYCLE_ACTIVE_rep26_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12843),
            .ce(N__12626),
            .sr(N__12473));
    defparam D_LL_AMIGA_iobuf_RNO_1_LC_1_4_1.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_1_LC_1_4_1.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_1_LC_1_4_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_1_LC_1_4_1 (
            .in0(N__4430),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_238_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep24_i_ess_LC_1_5_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep24_i_ess_LC_1_5_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep24_i_ess_LC_1_5_4 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep24_i_ess_LC_1_5_4  (
            .in0(N__11077),
            .in1(N__12167),
            .in2(N__11630),
            .in3(N__10586),
            .lcout(WRITE_CYCLE_ACTIVE_rep24_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12837),
            .ce(N__12620),
            .sr(N__12469));
    defparam D_LL_AMIGA_iobuf_RNO_5_LC_1_6_4.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_5_LC_1_6_4.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_5_LC_1_6_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_5_LC_1_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4241),
            .lcout(N_242_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_AMIGA_iobuf_RNO_6_LC_1_6_5.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_6_LC_1_6_5.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_6_LC_1_6_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_6_LC_1_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4424),
            .lcout(N_243_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_AMIGA_iobuf_RNO_0_LC_1_7_3.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_0_LC_1_7_3.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_0_LC_1_7_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_0_LC_1_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4412),
            .lcout(N_229_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_AMIGA_iobuf_RNO_7_LC_1_7_7.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_7_LC_1_7_7.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_7_LC_1_7_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_7_LC_1_7_7 (
            .in0(N__4418),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_244_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep17_i_ess_LC_1_8_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep17_i_ess_LC_1_8_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep17_i_ess_LC_1_8_6 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep17_i_ess_LC_1_8_6  (
            .in0(N__10573),
            .in1(N__12116),
            .in2(N__11759),
            .in3(N__11023),
            .lcout(WRITE_CYCLE_ACTIVE_rep17_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12831),
            .ce(N__12614),
            .sr(N__12462));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep29_i_ess_LC_1_8_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep29_i_ess_LC_1_8_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep29_i_ess_LC_1_8_7 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep29_i_ess_LC_1_8_7  (
            .in0(N__11024),
            .in1(N__12117),
            .in2(N__10585),
            .in3(N__11748),
            .lcout(WRITE_CYCLE_ACTIVE_rep29_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12831),
            .ce(N__12614),
            .sr(N__12462));
    defparam D_LM_AMIGA_iobuf_RNO_1_LC_1_9_6.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_1_LC_1_9_6.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_1_LC_1_9_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_1_LC_1_9_6 (
            .in0(N__4232),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_230_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_1_10_2.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_1_10_2.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_1_10_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_1_10_2 (
            .in0(N__7241),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIICIM_0_LC_1_10_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIICIM_0_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIICIM_0_LC_1_10_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIICIM_0_LC_1_10_4  (
            .in0(N__12515),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6770),
            .lcout(\U111_CYCLE_SM.CYCLE_STATE_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_0_LC_1_12_6.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_0_LC_1_12_6.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_0_LC_1_12_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_0_LC_1_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4541),
            .lcout(N_221_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_2_LC_1_13_1.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_2_LC_1_13_1.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_2_LC_1_13_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_2_LC_1_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4379),
            .lcout(N_223_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_AMIGA_iobuf_RNO_4_LC_1_13_3.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_4_LC_1_13_3.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_4_LC_1_13_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_4_LC_1_13_3 (
            .in0(N__4535),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_233_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep10_i_ess_LC_1_14_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep10_i_ess_LC_1_14_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep10_i_ess_LC_1_14_4 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep10_i_ess_LC_1_14_4  (
            .in0(N__11109),
            .in1(N__12022),
            .in2(N__11716),
            .in3(N__10535),
            .lcout(WRITE_CYCLE_ACTIVE_rep10_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12820),
            .ce(N__12615),
            .sr(N__12466));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep9_i_ess_LC_1_14_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep9_i_ess_LC_1_14_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep9_i_ess_LC_1_14_7 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep9_i_ess_LC_1_14_7  (
            .in0(N__12023),
            .in1(N__11688),
            .in2(N__10572),
            .in3(N__11113),
            .lcout(WRITE_CYCLE_ACTIVE_rep9_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12820),
            .ce(N__12615),
            .sr(N__12466));
    defparam D_LM_AMIGA_iobuf_RNO_5_LC_1_15_1.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_5_LC_1_15_1.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_5_LC_1_15_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_5_LC_1_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4874),
            .lcout(N_234_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_1_LC_1_15_3.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_1_LC_1_15_3.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_1_LC_1_15_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_1_LC_1_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4361),
            .lcout(N_222_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_AMIGA_iobuf_RNO_7_LC_1_17_3.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_7_LC_1_17_3.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_7_LC_1_17_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_7_LC_1_17_3 (
            .in0(N__4865),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_236_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_AMIGA_iobuf_RNO_6_LC_1_17_5.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_6_LC_1_17_5.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_6_LC_1_17_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_6_LC_1_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4523),
            .lcout(N_235_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_3_LC_1_17_7.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_3_LC_1_17_7.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_3_LC_1_17_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_3_LC_1_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4529),
            .lcout(N_224_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_6_LC_1_18_6.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_6_LC_1_18_6.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_6_LC_1_18_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_6_LC_1_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4517),
            .lcout(N_227_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_AMIGA_iobuf_RNO_1_LC_1_18_7.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_1_LC_1_18_7.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_1_LC_1_18_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_1_LC_1_18_7 (
            .in0(N__4511),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_214_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_7_LC_1_19_1.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_7_LC_1_19_1.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_7_LC_1_19_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_7_LC_1_19_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4454),
            .lcout(N_228_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_4_LC_1_19_4.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_4_LC_1_19_4.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_4_LC_1_19_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_4_LC_1_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4505),
            .lcout(N_225_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep15_i_ess_LC_1_20_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep15_i_ess_LC_1_20_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep15_i_ess_LC_1_20_4 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep15_i_ess_LC_1_20_4  (
            .in0(N__10571),
            .in1(N__12166),
            .in2(N__11703),
            .in3(N__11168),
            .lcout(WRITE_CYCLE_ACTIVE_rep15_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12798),
            .ce(N__12630),
            .sr(N__12487));
    defparam D_LL_AMIGA_iobuf_RNO_4_LC_2_3_5.C_ON=1'b0;
    defparam D_LL_AMIGA_iobuf_RNO_4_LC_2_3_5.SEQ_MODE=4'b0000;
    defparam D_LL_AMIGA_iobuf_RNO_4_LC_2_3_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_AMIGA_iobuf_RNO_4_LC_2_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4589),
            .lcout(N_241_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep25_i_ess_LC_2_4_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep25_i_ess_LC_2_4_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep25_i_ess_LC_2_4_1 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep25_i_ess_LC_2_4_1  (
            .in0(N__10883),
            .in1(N__12243),
            .in2(N__11765),
            .in3(N__10584),
            .lcout(WRITE_CYCLE_ACTIVE_rep25_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12838),
            .ce(N__12627),
            .sr(N__12474));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep30_i_ess_LC_2_6_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep30_i_ess_LC_2_6_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep30_i_ess_LC_2_6_5 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep30_i_ess_LC_2_6_5  (
            .in0(N__10884),
            .in1(N__12089),
            .in2(N__11760),
            .in3(N__10582),
            .lcout(WRITE_CYCLE_ACTIVE_rep30_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12834),
            .ce(N__12621),
            .sr(N__12470));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_i_ess_LC_2_7_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_i_ess_LC_2_7_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_i_ess_LC_2_7_1 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_i_ess_LC_2_7_1  (
            .in0(N__12206),
            .in1(N__11744),
            .in2(N__10992),
            .in3(N__10581),
            .lcout(WRITE_CYCLE_ACTIVE_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12832),
            .ce(N__12619),
            .sr(N__12467));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep16_i_ess_LC_2_8_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep16_i_ess_LC_2_8_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep16_i_ess_LC_2_8_5 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep16_i_ess_LC_2_8_5  (
            .in0(N__10993),
            .in1(N__12205),
            .in2(N__11758),
            .in3(N__10554),
            .lcout(WRITE_CYCLE_ACTIVE_rep16_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12827),
            .ce(N__12617),
            .sr(N__12463));
    defparam D_LM_AMIGA_iobuf_RNO_3_LC_2_11_7.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_3_LC_2_11_7.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_3_LC_2_11_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_3_LC_2_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4571),
            .lcout(N_232_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep8_i_ess_LC_2_12_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep8_i_ess_LC_2_12_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep8_i_ess_LC_2_12_5 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep8_i_ess_LC_2_12_5  (
            .in0(N__11079),
            .in1(N__12204),
            .in2(N__11740),
            .in3(N__10504),
            .lcout(WRITE_CYCLE_ACTIVE_rep8_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12822),
            .ce(N__12613),
            .sr(N__12464));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep20_i_ess_LC_2_13_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep20_i_ess_LC_2_13_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep20_i_ess_LC_2_13_4 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep20_i_ess_LC_2_13_4  (
            .in0(N__12202),
            .in1(N__10503),
            .in2(N__11137),
            .in3(N__11588),
            .lcout(WRITE_CYCLE_ACTIVE_rep20_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12821),
            .ce(N__12616),
            .sr(N__12468));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep11_i_ess_LC_2_16_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep11_i_ess_LC_2_16_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep11_i_ess_LC_2_16_6 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep11_i_ess_LC_2_16_6  (
            .in0(N__12227),
            .in1(N__10485),
            .in2(N__11167),
            .in3(N__11684),
            .lcout(WRITE_CYCLE_ACTIVE_rep11_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12815),
            .ce(N__12622),
            .sr(N__12475));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep5_i_ess_LC_2_17_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep5_i_ess_LC_2_17_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep5_i_ess_LC_2_17_1 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep5_i_ess_LC_2_17_1  (
            .in0(N__11632),
            .in1(N__12230),
            .in2(N__10549),
            .in3(N__11150),
            .lcout(WRITE_CYCLE_ACTIVE_rep5_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12810),
            .ce(N__12624),
            .sr(N__12477));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep22_i_ess_LC_2_17_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep22_i_ess_LC_2_17_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep22_i_ess_LC_2_17_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep22_i_ess_LC_2_17_5  (
            .in0(N__11631),
            .in1(N__12229),
            .in2(N__10548),
            .in3(N__11149),
            .lcout(WRITE_CYCLE_ACTIVE_rep22_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12810),
            .ce(N__12624),
            .sr(N__12477));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep14_i_ess_LC_2_18_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep14_i_ess_LC_2_18_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep14_i_ess_LC_2_18_1 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep14_i_ess_LC_2_18_1  (
            .in0(N__10493),
            .in1(N__12252),
            .in2(N__11166),
            .in3(N__11649),
            .lcout(WRITE_CYCLE_ACTIVE_rep14_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12805),
            .ce(N__12628),
            .sr(N__12482));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep1_i_ess_LC_2_18_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep1_i_ess_LC_2_18_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep1_i_ess_LC_2_18_4 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep1_i_ess_LC_2_18_4  (
            .in0(N__11650),
            .in1(N__10494),
            .in2(N__12260),
            .in3(N__11142),
            .lcout(WRITE_CYCLE_ACTIVE_rep1_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12805),
            .ce(N__12628),
            .sr(N__12482));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep12_i_ess_LC_2_19_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep12_i_ess_LC_2_19_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep12_i_ess_LC_2_19_1 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep12_i_ess_LC_2_19_1  (
            .in0(N__11144),
            .in1(N__12257),
            .in2(N__11705),
            .in3(N__10498),
            .lcout(WRITE_CYCLE_ACTIVE_rep12_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12799),
            .ce(N__12631),
            .sr(N__12488));
    defparam D_UU_AMIGA_iobuf_RNO_3_LC_2_20_3.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_3_LC_2_20_3.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_3_LC_2_20_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_3_LC_2_20_3 (
            .in0(N__4829),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_216_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_AMIGA_iobuf_RNO_5_LC_2_20_7.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_5_LC_2_20_7.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_5_LC_2_20_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_5_LC_2_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4652),
            .lcout(N_218_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_0  (
            .in0(N__4628),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6025),
            .lcout(A_AMIGA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_3  (
            .in0(N__6026),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4891),
            .lcout(U111_CYCLE_SM_A_AMIGA_0_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep28_i_ess_LC_3_3_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep28_i_ess_LC_3_3_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep28_i_ess_LC_3_3_7 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep28_i_ess_LC_3_3_7  (
            .in0(N__10381),
            .in1(N__12244),
            .in2(N__11654),
            .in3(N__10693),
            .lcout(WRITE_CYCLE_ACTIVE_rep28_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12839),
            .ce(N__12634),
            .sr(N__12484));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep27_i_ess_LC_3_4_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep27_i_ess_LC_3_4_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep27_i_ess_LC_3_4_5 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep27_i_ess_LC_3_4_5  (
            .in0(N__12242),
            .in1(N__11589),
            .in2(N__11076),
            .in3(N__10583),
            .lcout(WRITE_CYCLE_ACTIVE_rep27_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12836),
            .ce(N__12632),
            .sr(N__12478));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep19_i_ess_LC_3_11_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep19_i_ess_LC_3_11_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep19_i_ess_LC_3_11_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep19_i_ess_LC_3_11_5  (
            .in0(N__10569),
            .in1(N__12203),
            .in2(N__11584),
            .in3(N__10994),
            .lcout(WRITE_CYCLE_ACTIVE_rep19_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12823),
            .ce(N__12612),
            .sr(N__12465));
    defparam D_LM_AMIGA_iobuf_RNO_2_LC_3_12_3.C_ON=1'b0;
    defparam D_LM_AMIGA_iobuf_RNO_2_LC_3_12_3.SEQ_MODE=4'b0000;
    defparam D_LM_AMIGA_iobuf_RNO_2_LC_3_12_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LM_AMIGA_iobuf_RNO_2_LC_3_12_3 (
            .in0(N__4556),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_231_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep18_i_ess_LC_3_13_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep18_i_ess_LC_3_13_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep18_i_ess_LC_3_13_1 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep18_i_ess_LC_3_13_1  (
            .in0(N__10502),
            .in1(N__12171),
            .in2(N__11587),
            .in3(N__11078),
            .lcout(WRITE_CYCLE_ACTIVE_rep18_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12819),
            .ce(N__12618),
            .sr(N__12471));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep21_i_ess_LC_3_15_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep21_i_ess_LC_3_15_3 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep21_i_ess_LC_3_15_3 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep21_i_ess_LC_3_15_3  (
            .in0(N__11506),
            .in1(N__12217),
            .in2(N__10372),
            .in3(N__11083),
            .lcout(WRITE_CYCLE_ACTIVE_rep21_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12816),
            .ce(N__12623),
            .sr(N__12476));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep23_i_ess_LC_3_16_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep23_i_ess_LC_3_16_2 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep23_i_ess_LC_3_16_2 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep23_i_ess_LC_3_16_2  (
            .in0(N__12226),
            .in1(N__11505),
            .in2(N__10568),
            .in3(N__11138),
            .lcout(WRITE_CYCLE_ACTIVE_rep23_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12811),
            .ce(N__12625),
            .sr(N__12479));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep7_i_ess_LC_3_17_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep7_i_ess_LC_3_17_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep7_i_ess_LC_3_17_7 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep7_i_ess_LC_3_17_7  (
            .in0(N__10486),
            .in1(N__12228),
            .in2(N__11453),
            .in3(N__11148),
            .lcout(WRITE_CYCLE_ACTIVE_rep7_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12806),
            .ce(N__12629),
            .sr(N__12483));
    defparam D_UU_AMIGA_iobuf_RNO_7_LC_3_18_1.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_7_LC_3_18_1.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_7_LC_3_18_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_7_LC_3_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4853),
            .lcout(N_220_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep3_i_ess_LC_3_19_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep3_i_ess_LC_3_19_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep3_i_ess_LC_3_19_1 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep3_i_ess_LC_3_19_1  (
            .in0(N__11601),
            .in1(N__12256),
            .in2(N__10550),
            .in3(N__11143),
            .lcout(WRITE_CYCLE_ACTIVE_rep3_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12793),
            .ce(N__12633),
            .sr(N__12490));
    defparam D_UU_AMIGA_iobuf_RNO_6_LC_3_20_5.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_6_LC_3_20_5.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_6_LC_3_20_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_6_LC_3_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4943),
            .lcout(N_219_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_5_1_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_5_1_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_5_1_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_5_1_6  (
            .in0(N__8827),
            .in1(N__4808),
            .in2(_gnd_net_),
            .in3(N__8975),
            .lcout(un2_D_LL_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_5_10_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_5_10_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_5_10_4  (
            .in0(N__8735),
            .in1(N__6530),
            .in2(_gnd_net_),
            .in3(N__4778),
            .lcout(un2_D_LM_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_5_10_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_5_10_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_5_10_6  (
            .in0(N__4745),
            .in1(N__8741),
            .in2(_gnd_net_),
            .in3(N__4729),
            .lcout(un1_D_UM_040_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_5_12_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_5_12_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_5_12_2  (
            .in0(N__5081),
            .in1(N__5053),
            .in2(_gnd_net_),
            .in3(N__8792),
            .lcout(un1_D_UM_040_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_5_12_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_5_12_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_5_12_5  (
            .in0(N__8791),
            .in1(N__7698),
            .in2(_gnd_net_),
            .in3(N__5009),
            .lcout(un2_D_LM_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep0_i_ess_LC_5_18_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep0_i_ess_LC_5_18_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep0_i_ess_LC_5_18_7 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep0_i_ess_LC_5_18_7  (
            .in0(N__10461),
            .in1(N__12251),
            .in2(N__11182),
            .in3(N__11560),
            .lcout(WRITE_CYCLE_ACTIVE_rep0_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12790),
            .ce(N__12635),
            .sr(N__12491));
    defparam D_UU_AMIGA_iobuf_RNO_0_LC_5_19_3.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_0_LC_5_19_3.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_0_LC_5_19_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_0_LC_5_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4982),
            .lcout(N_213_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_AMIGA_iobuf_RNO_5_LC_5_19_4.C_ON=1'b0;
    defparam D_UM_AMIGA_iobuf_RNO_5_LC_5_19_4.SEQ_MODE=4'b0000;
    defparam D_UM_AMIGA_iobuf_RNO_5_LC_5_19_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_AMIGA_iobuf_RNO_5_LC_5_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5303),
            .lcout(N_226_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep4_i_ess_LC_5_20_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep4_i_ess_LC_5_20_3 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep4_i_ess_LC_5_20_3 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep4_i_ess_LC_5_20_3  (
            .in0(N__12073),
            .in1(N__11558),
            .in2(N__11183),
            .in3(N__10528),
            .lcout(WRITE_CYCLE_ACTIVE_rep4_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12784),
            .ce(N__12638),
            .sr(N__12493));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep6_i_ess_LC_5_20_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep6_i_ess_LC_5_20_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep6_i_ess_LC_5_20_6 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep6_i_ess_LC_5_20_6  (
            .in0(N__11559),
            .in1(N__12074),
            .in2(N__10570),
            .in3(N__11181),
            .lcout(WRITE_CYCLE_ACTIVE_rep6_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12784),
            .ce(N__12638),
            .sr(N__12493));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_6_3_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_6_3_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_6_3_1  (
            .in0(N__6963),
            .in1(N__4934),
            .in2(_gnd_net_),
            .in3(N__8828),
            .lcout(un2_D_LL_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_6_6_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_6_6_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_6_6_4  (
            .in0(N__6088),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4901),
            .lcout(\U111_CYCLE_SM.FLIP_WORD_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep13_i_ess_LC_6_19_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep13_i_ess_LC_6_19_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep13_i_ess_LC_6_19_6 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep13_i_ess_LC_6_19_6  (
            .in0(N__11161),
            .in1(N__12259),
            .in2(N__11655),
            .in3(N__10527),
            .lcout(WRITE_CYCLE_ACTIVE_rep13_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12783),
            .ce(N__12637),
            .sr(N__12492));
    defparam D_UU_AMIGA_iobuf_RNO_4_LC_6_20_2.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_4_LC_6_20_2.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_4_LC_6_20_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_4_LC_6_20_2 (
            .in0(N__5297),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_217_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_7_3_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_7_3_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_7_3_1  (
            .in0(N__5276),
            .in1(N__8465),
            .in2(_gnd_net_),
            .in3(N__8823),
            .lcout(un2_D_LL_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_7_9_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_7_9_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_7_9_1  (
            .in0(N__5239),
            .in1(N__5195),
            .in2(_gnd_net_),
            .in3(N__8710),
            .lcout(un1_D_UM_040_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_7_11_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_7_11_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_7_11_2  (
            .in0(N__8645),
            .in1(N__8006),
            .in2(_gnd_net_),
            .in3(N__5159),
            .lcout(un2_D_LM_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep2_i_ess_LC_7_19_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep2_i_ess_LC_7_19_3 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep2_i_ess_LC_7_19_3 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_rep2_i_ess_LC_7_19_3  (
            .in0(N__11522),
            .in1(N__12258),
            .in2(N__10454),
            .in3(N__11157),
            .lcout(WRITE_CYCLE_ACTIVE_rep2_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12782),
            .ce(N__12639),
            .sr(N__12494));
    defparam BUFENn_obuf_RNO_LC_7_20_0.C_ON=1'b0;
    defparam BUFENn_obuf_RNO_LC_7_20_0.SEQ_MODE=4'b0000;
    defparam BUFENn_obuf_RNO_LC_7_20_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 BUFENn_obuf_RNO_LC_7_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11174),
            .lcout(LBENn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_AMIGA_iobuf_RNO_2_LC_7_20_6.C_ON=1'b0;
    defparam D_UU_AMIGA_iobuf_RNO_2_LC_7_20_6.SEQ_MODE=4'b0000;
    defparam D_UU_AMIGA_iobuf_RNO_2_LC_7_20_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_AMIGA_iobuf_RNO_2_LC_7_20_6 (
            .in0(N__5105),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_215_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_7_20_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_7_20_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_7_20_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_7_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_8_3_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_8_3_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_8_3_2  (
            .in0(N__9392),
            .in1(N__5687),
            .in2(_gnd_net_),
            .in3(N__8768),
            .lcout(un2_D_LL_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_8_7_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_8_7_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_8_7_6  (
            .in0(N__8769),
            .in1(N__6887),
            .in2(_gnd_net_),
            .in3(N__5648),
            .lcout(un2_D_LM_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TSn_LC_8_9_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TSn_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TSn_LC_8_9_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U111_CYCLE_SM.TSn_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__7240),
            .in2(_gnd_net_),
            .in3(N__5593),
            .lcout(TSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.TSnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_LC_8_10_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_LC_8_10_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TS_EN_LC_8_10_6 .LUT_INIT=16'b1110010011111111;
    LogicCell40 \U111_CYCLE_SM.TS_EN_LC_8_10_6  (
            .in0(N__6722),
            .in1(N__5594),
            .in2(N__5717),
            .in3(N__5729),
            .lcout(\U111_CYCLE_SM.TS_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12812),
            .ce(),
            .sr(N__12472));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_8_15_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_8_15_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_8_15_0  (
            .in0(N__5582),
            .in1(N__5557),
            .in2(_gnd_net_),
            .in3(N__8745),
            .lcout(un1_D_UM_040_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_8_17_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_8_17_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_8_17_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_8_17_5  (
            .in0(N__8746),
            .in1(N__7920),
            .in2(_gnd_net_),
            .in3(N__5501),
            .lcout(un2_D_LM_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_8_18_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_8_18_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_8_18_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_8_18_7  (
            .in0(N__5455),
            .in1(N__5429),
            .in2(_gnd_net_),
            .in3(N__8747),
            .lcout(un1_D_UU_040_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_8_20_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_8_20_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_8_20_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_8_20_1  (
            .in0(N__8797),
            .in1(N__5395),
            .in2(_gnd_net_),
            .in3(N__5345),
            .lcout(un1_D_UM_040_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_8_20_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_8_20_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_8_20_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_8_20_5  (
            .in0(N__8798),
            .in1(N__5840),
            .in2(_gnd_net_),
            .in3(N__5815),
            .lcout(un1_D_UU_040_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_9_2_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_9_2_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_9_2_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_9_2_5  (
            .in0(N__8734),
            .in1(N__5762),
            .in2(_gnd_net_),
            .in3(N__7540),
            .lcout(un2_D_LL_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LATCH_EN_LC_9_9_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LATCH_EN_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.LATCH_EN_LC_9_9_4 .LUT_INIT=16'b1100000011100010;
    LogicCell40 \U111_CYCLE_SM.LATCH_EN_LC_9_9_4  (
            .in0(N__6689),
            .in1(N__5728),
            .in2(N__9025),
            .in3(N__6766),
            .lcout(\U111_CYCLE_SM.LATCH_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12813),
            .ce(),
            .sr(N__12480));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIDUAQ_0_LC_9_10_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIDUAQ_0_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIDUAQ_0_LC_9_10_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIDUAQ_0_LC_9_10_0  (
            .in0(N__12094),
            .in1(N__11704),
            .in2(N__11133),
            .in3(N__6760),
            .lcout(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ),
            .ltout(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIC4111_3_LC_9_10_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIC4111_3_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIC4111_3_LC_9_10_1 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIC4111_3_LC_9_10_1  (
            .in0(N__6181),
            .in1(_gnd_net_),
            .in2(N__5732),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.un1_CYCLE_STATE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_4_LC_9_10_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_4_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_4_LC_9_10_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_4_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(N__7242),
            .in2(_gnd_net_),
            .in3(N__6182),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12807),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_RNO_1_LC_9_10_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_RNO_1_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN_RNO_1_LC_9_10_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U111_CYCLE_SM.TS_EN_RNO_1_LC_9_10_5  (
            .in0(N__6180),
            .in1(N__6598),
            .in2(N__7186),
            .in3(N__6228),
            .lcout(\U111_CYCLE_SM.TS_EN_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.BURST_LC_9_11_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_LC_9_11_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.BURST_LC_9_11_0 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U111_CYCLE_SM.BURST_LC_9_11_0  (
            .in0(N__6639),
            .in1(N__6154),
            .in2(N__6133),
            .in3(N__6599),
            .lcout(\U111_CYCLE_SM.BURSTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12800),
            .ce(),
            .sr(N__12481));
    defparam \U111_CYCLE_SM.BURST_COUNT_1_LC_9_11_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_COUNT_1_LC_9_11_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.BURST_COUNT_1_LC_9_11_1 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \U111_CYCLE_SM.BURST_COUNT_1_LC_9_11_1  (
            .in0(N__6671),
            .in1(N__6638),
            .in2(N__6302),
            .in3(N__6617),
            .lcout(\U111_CYCLE_SM.BURST_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12800),
            .ce(),
            .sr(N__12481));
    defparam \U111_CYCLE_SM.LW_TRANS_LC_9_11_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_TRANS_LC_9_11_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.LW_TRANS_LC_9_11_2 .LUT_INIT=16'b1101011110000010;
    LogicCell40 \U111_CYCLE_SM.LW_TRANS_LC_9_11_2  (
            .in0(N__6640),
            .in1(N__6155),
            .in2(N__6134),
            .in3(N__6046),
            .lcout(\U111_CYCLE_SM.LW_TRANSZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12800),
            .ce(),
            .sr(N__12481));
    defparam \U111_CYCLE_SM.TA_DIS_LC_9_11_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_DIS_LC_9_11_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TA_DIS_LC_9_11_3 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \U111_CYCLE_SM.TA_DIS_LC_9_11_3  (
            .in0(N__6184),
            .in1(N__6237),
            .in2(N__7123),
            .in3(N__6032),
            .lcout(\U111_CYCLE_SM.TA_DISZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12800),
            .ce(),
            .sr(N__12481));
    defparam \U111_CYCLE_SM.FLIP_WORD_LC_9_11_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_LC_9_11_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.FLIP_WORD_LC_9_11_5 .LUT_INIT=16'b1111000011101110;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_LC_9_11_5  (
            .in0(N__8596),
            .in1(N__6183),
            .in2(N__6110),
            .in3(N__6238),
            .lcout(\U111_CYCLE_SM.FLIP_WORDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12800),
            .ce(),
            .sr(N__12481));
    defparam \U111_CYCLE_SM.PORT_MISMATCH_LC_9_11_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.PORT_MISMATCH_LC_9_11_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.PORT_MISMATCH_LC_9_11_7 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \U111_CYCLE_SM.PORT_MISMATCH_LC_9_11_7  (
            .in0(N__6047),
            .in1(N__6239),
            .in2(N__6212),
            .in3(N__6084),
            .lcout(\U111_CYCLE_SM.PORT_MISMATCHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12800),
            .ce(),
            .sr(N__12481));
    defparam \U111_CYCLE_SM.TA_DIS_RNO_0_LC_9_12_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_DIS_RNO_0_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_DIS_RNO_0_LC_9_12_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U111_CYCLE_SM.TA_DIS_RNO_0_LC_9_12_4  (
            .in0(N__6092),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6045),
            .lcout(\U111_CYCLE_SM.PORT_MISMATCH_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A2_EN_LC_9_12_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A2_EN_LC_9_12_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.A2_EN_LC_9_12_5 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \U111_CYCLE_SM.A2_EN_LC_9_12_5  (
            .in0(N__6188),
            .in1(N__6010),
            .in2(_gnd_net_),
            .in3(N__6553),
            .lcout(\U111_CYCLE_SM.A2_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12795),
            .ce(),
            .sr(N__12485));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_9_15_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_9_15_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_9_15_2  (
            .in0(N__7029),
            .in1(N__5999),
            .in2(_gnd_net_),
            .in3(N__8666),
            .lcout(un2_D_LM_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_9_20_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_9_20_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_9_20_3  (
            .in0(N__5959),
            .in1(N__5915),
            .in2(_gnd_net_),
            .in3(N__8796),
            .lcout(un1_D_UU_040_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_10_6_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_10_6_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_10_6_0  (
            .in0(N__8807),
            .in1(N__9332),
            .in2(_gnd_net_),
            .in3(N__5882),
            .lcout(un2_D_LL_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_1_LC_10_9_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_1_LC_10_9_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_1_LC_10_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_1_LC_10_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6522),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12808),
            .ce(N__7868),
            .sr(N__7796));
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_10_10_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_10_10_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_10_10_0 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_1_LC_10_10_0  (
            .in0(N__6641),
            .in1(N__6557),
            .in2(N__7254),
            .in3(N__6597),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12801),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_10_10_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_10_10_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(N__7166),
            .in2(_gnd_net_),
            .in3(N__6711),
            .lcout(\U111_CYCLE_SM.N_124_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_10_10_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_10_10_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_10_10_2  (
            .in0(N__6712),
            .in1(N__6206),
            .in2(N__7414),
            .in3(N__6251),
            .lcout(),
            .ltout(\U111_CYCLE_SM.N_132_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_10_10_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_10_10_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_10_10_3 .LUT_INIT=16'b1111000111111111;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_0_LC_10_10_3  (
            .in0(N__7329),
            .in1(N__6311),
            .in2(N__6305),
            .in3(N__6569),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12801),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_10_10_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_10_10_4 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_10_10_4  (
            .in0(N__6298),
            .in1(N__6615),
            .in2(N__6287),
            .in3(N__6596),
            .lcout(\U111_CYCLE_SM.un7_CYCLE_STATE_0 ),
            .ltout(\U111_CYCLE_SM.un7_CYCLE_STATE_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_10_10_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_10_10_5 .LUT_INIT=16'b0111011101010111;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_10_10_5  (
            .in0(N__7330),
            .in1(N__7405),
            .in2(N__6245),
            .in3(N__6207),
            .lcout(),
            .ltout(\U111_CYCLE_SM.CYCLE_STATE_srsts_i_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_2_LC_10_10_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_2_LC_10_10_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_2_LC_10_10_6 .LUT_INIT=16'b1100110000001000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_2_LC_10_10_6  (
            .in0(N__6713),
            .in1(N__7255),
            .in2(N__6242),
            .in3(N__6236),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12801),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_3_LC_10_10_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_3_LC_10_10_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_3_LC_10_10_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_3_LC_10_10_7  (
            .in0(N__6663),
            .in1(N__7246),
            .in2(_gnd_net_),
            .in3(N__6208),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12801),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.BURST_COUNT_0_LC_10_11_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_COUNT_0_LC_10_11_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.BURST_COUNT_0_LC_10_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U111_CYCLE_SM.BURST_COUNT_0_LC_10_11_2  (
            .in0(N__6637),
            .in1(N__6664),
            .in2(_gnd_net_),
            .in3(N__6616),
            .lcout(\U111_CYCLE_SM.BURST_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12796),
            .ce(),
            .sr(N__12486));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_3_0_LC_10_11_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_3_0_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_3_0_LC_10_11_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_3_0_LC_10_11_6  (
            .in0(N__7410),
            .in1(N__7150),
            .in2(_gnd_net_),
            .in3(N__6595),
            .lcout(),
            .ltout(\U111_CYCLE_SM.N_131_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_10_11_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_10_11_7 .LUT_INIT=16'b0000100000001100;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_10_11_7  (
            .in0(N__6563),
            .in1(N__7267),
            .in2(N__6572),
            .in3(N__6765),
            .lcout(\U111_CYCLE_SM.CYCLE_STATE_srsts_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_4_0_LC_10_12_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_4_0_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_4_0_LC_10_12_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_4_0_LC_10_12_2  (
            .in0(N__11037),
            .in1(N__12013),
            .in2(_gnd_net_),
            .in3(N__11605),
            .lcout(\U111_CYCLE_SM.TS_EN6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_10_12_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_10_12_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_10_12_4  (
            .in0(N__7409),
            .in1(N__7332),
            .in2(_gnd_net_),
            .in3(N__7154),
            .lcout(\U111_CYCLE_SM.N_144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIUR6Q_1_LC_10_18_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIUR6Q_1_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIUR6Q_1_LC_10_18_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNIUR6Q_1_LC_10_18_5  (
            .in0(N__6542),
            .in1(N__6523),
            .in2(_gnd_net_),
            .in3(N__9096),
            .lcout(un1_D_UU_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_10_18_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_10_18_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_10_18_7  (
            .in0(N__6461),
            .in1(N__6446),
            .in2(_gnd_net_),
            .in3(N__8781),
            .lcout(un1_D_UM_040_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_10_20_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_10_20_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_10_20_7  (
            .in0(N__6373),
            .in1(N__6344),
            .in2(_gnd_net_),
            .in3(N__8815),
            .lcout(un1_D_UU_040_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LBENn_c_sbtinv_LC_11_1_0.C_ON=1'b0;
    defparam LBENn_c_sbtinv_LC_11_1_0.SEQ_MODE=4'b0000;
    defparam LBENn_c_sbtinv_LC_11_1_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 LBENn_c_sbtinv_LC_11_1_0 (
            .in0(N__10686),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(LBENn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_11_7_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_11_7_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_11_7_3  (
            .in0(N__8808),
            .in1(N__8318),
            .in2(_gnd_net_),
            .in3(N__6809),
            .lcout(un2_D_LL_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_RNO_2_LC_11_8_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_RNO_2_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN_RNO_2_LC_11_8_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U111_CYCLE_SM.TS_EN_RNO_2_LC_11_8_0  (
            .in0(N__7368),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7311),
            .lcout(\U111_CYCLE_SM.N_119_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_LC_11_9_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_LC_11_9_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_LC_11_9_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_LC_11_9_0  (
            .in0(N__10567),
            .in1(N__12093),
            .in2(N__11585),
            .in3(N__10876),
            .lcout(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12802),
            .ce(N__12636),
            .sr(N__12489));
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_10_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_10_2 .LUT_INIT=16'b0001000000010001;
    LogicCell40 \U111_CYCLE_SM.TS_EN_RNO_0_LC_11_10_2  (
            .in0(N__6710),
            .in1(N__6764),
            .in2(N__6734),
            .in3(N__7161),
            .lcout(\U111_CYCLE_SM.N_117_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_11_10_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_11_10_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_11_10_3  (
            .in0(N__7386),
            .in1(N__7331),
            .in2(_gnd_net_),
            .in3(N__6709),
            .lcout(\U111_CYCLE_SM.BURST_COUNT_0_sqmuxa ),
            .ltout(\U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3B1_LC_11_10_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3B1_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3B1_LC_11_10_4 .LUT_INIT=16'b0101010111110101;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3B1_LC_11_10_4  (
            .in0(N__7253),
            .in1(_gnd_net_),
            .in2(N__6692),
            .in3(N__6685),
            .lcout(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1 ),
            .ltout(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_esr_RNIPC3BZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI9Q9V1_2_LC_11_10_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI9Q9V1_2_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI9Q9V1_2_LC_11_10_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNI9Q9V1_2_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6674),
            .in3(N__6662),
            .lcout(\U111_CYCLE_SM.BURST_COUNT_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_5_LC_11_11_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_5_LC_11_11_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_5_LC_11_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_5_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7031),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12792),
            .ce(N__7858),
            .sr(N__7794));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_11_11_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_11_11_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_11_11_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_1_LC_11_11_5  (
            .in0(N__6968),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12792),
            .ce(N__7858),
            .sr(N__7794));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_0_LC_11_11_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_0_LC_11_11_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_0_LC_11_11_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_0_LC_11_11_7  (
            .in0(N__6886),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12792),
            .ce(N__7858),
            .sr(N__7794));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_11_12_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_11_12_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_11_12_6  (
            .in0(N__7387),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7333),
            .lcout(),
            .ltout(\U111_CYCLE_SM.CYCLE_STATE_srsts_i_o2_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_5_LC_11_12_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_5_LC_11_12_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_5_LC_11_12_7 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_5_LC_11_12_7  (
            .in0(N__7268),
            .in1(N__7190),
            .in2(N__7169),
            .in3(N__7165),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12788),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_11_13_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_11_13_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__11038),
            .in2(_gnd_net_),
            .in3(N__7127),
            .lcout(TAn_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_11_13_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_11_13_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_11_13_2  (
            .in0(N__7085),
            .in1(N__7600),
            .in2(_gnd_net_),
            .in3(N__8721),
            .lcout(un2_D_LM_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI647Q_5_LC_11_15_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI647Q_5_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI647Q_5_LC_11_15_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNI647Q_5_LC_11_15_3  (
            .in0(N__9105),
            .in1(N__7043),
            .in2(_gnd_net_),
            .in3(N__7030),
            .lcout(un1_D_UU_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_11_15_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_11_15_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIEBFL_1_LC_11_15_6  (
            .in0(N__6964),
            .in1(N__6926),
            .in2(_gnd_net_),
            .in3(N__9104),
            .lcout(un1_D_UM_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNISP6Q_0_LC_11_17_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNISP6Q_0_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNISP6Q_0_LC_11_17_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNISP6Q_0_LC_11_17_2  (
            .in0(N__6896),
            .in1(N__6867),
            .in2(_gnd_net_),
            .in3(N__9107),
            .lcout(un1_D_UU_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_12_6_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_12_6_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_12_6_7  (
            .in0(N__7457),
            .in1(N__8261),
            .in2(_gnd_net_),
            .in3(N__8756),
            .lcout(un2_D_LL_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_12_9_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_12_9_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_12_9_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_0_LC_12_9_6  (
            .in0(N__8967),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12794),
            .ce(N__7865),
            .sr(N__7797));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_12_10_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_12_10_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_12_10_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_7_LC_12_10_3  (
            .in0(N__8311),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12791),
            .ce(N__7867),
            .sr(N__7795));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_6_LC_12_10_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_6_LC_12_10_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_6_LC_12_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_6_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7928),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12791),
            .ce(N__7867),
            .sr(N__7795));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_12_10_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_12_10_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_12_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_2_LC_12_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9384),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12791),
            .ce(N__7867),
            .sr(N__7795));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_3_LC_12_11_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_3_LC_12_11_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_3_LC_12_11_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_3_LC_12_11_0  (
            .in0(N__8005),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12787),
            .ce(N__7866),
            .sr(N__7798));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_12_11_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_12_11_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_12_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_4_LC_12_11_1  (
            .in0(N__8464),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12787),
            .ce(N__7866),
            .sr(N__7798));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_12_11_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_12_11_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_12_11_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_6_LC_12_11_2  (
            .in0(N__9321),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12787),
            .ce(N__7866),
            .sr(N__7798));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_7_LC_12_11_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_7_LC_12_11_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_7_LC_12_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_7_LC_12_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8375),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12787),
            .ce(N__7866),
            .sr(N__7798));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_12_11_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_12_11_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_12_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_3_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7541),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12787),
            .ce(N__7866),
            .sr(N__7798));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_4_LC_12_11_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_4_LC_12_11_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_4_LC_12_11_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_4_LC_12_11_6  (
            .in0(N__7599),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12787),
            .ce(N__7866),
            .sr(N__7798));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_12_11_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_12_11_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_12_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_5_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8256),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12787),
            .ce(N__7866),
            .sr(N__7798));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_2_LC_12_12_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_2_LC_12_12_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_2_LC_12_12_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_2_LC_12_12_1  (
            .in0(N__7700),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12785),
            .ce(N__7857),
            .sr(N__7805));
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_13_6.C_ON=1'b0;
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_13_6.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7763),
            .lcout(GB_BUFFER_CLK80_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI0U6Q_2_LC_12_14_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI0U6Q_2_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI0U6Q_2_LC_12_14_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNI0U6Q_2_LC_12_14_0  (
            .in0(N__9085),
            .in1(N__7709),
            .in2(_gnd_net_),
            .in3(N__7699),
            .lcout(un1_D_UU_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIA87Q_7_LC_12_14_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIA87Q_7_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNIA87Q_7_LC_12_14_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNIA87Q_7_LC_12_14_1  (
            .in0(N__8371),
            .in1(N__7640),
            .in2(_gnd_net_),
            .in3(N__9089),
            .lcout(un1_D_UU_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI427Q_4_LC_12_14_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI427Q_4_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI427Q_4_LC_12_14_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNI427Q_4_LC_12_14_2  (
            .in0(N__7610),
            .in1(_gnd_net_),
            .in2(N__9106),
            .in3(N__7601),
            .lcout(un1_D_UU_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_12_16_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_12_16_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIIFFL_3_LC_12_16_1  (
            .in0(N__7536),
            .in1(N__7490),
            .in2(_gnd_net_),
            .in3(N__9090),
            .lcout(un1_D_UM_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_12_16_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_12_16_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIKHFL_4_LC_12_16_4  (
            .in0(N__9091),
            .in1(N__8474),
            .in2(_gnd_net_),
            .in3(N__8457),
            .lcout(un1_D_UM_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_12_17_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_12_17_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_12_17_7  (
            .in0(N__8393),
            .in1(N__8370),
            .in2(_gnd_net_),
            .in3(N__8757),
            .lcout(un2_D_LM_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_12_19_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_12_19_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIQNFL_7_LC_12_19_5  (
            .in0(N__9095),
            .in1(N__8327),
            .in2(_gnd_net_),
            .in3(N__8310),
            .lcout(un1_D_UM_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_12_20_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_12_20_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIMJFL_5_LC_12_20_0  (
            .in0(N__8260),
            .in1(N__8213),
            .in2(_gnd_net_),
            .in3(N__9108),
            .lcout(un1_D_UM_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_12_20_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_12_20_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_12_20_2  (
            .in0(N__8177),
            .in1(N__8159),
            .in2(_gnd_net_),
            .in3(N__8799),
            .lcout(un1_D_UU_040_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_12_20_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_12_20_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_12_20_3  (
            .in0(N__8800),
            .in1(N__8096),
            .in2(_gnd_net_),
            .in3(N__8068),
            .lcout(un1_D_UU_040_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI207Q_3_LC_12_20_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI207Q_3_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI207Q_3_LC_12_20_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNI207Q_3_LC_12_20_4  (
            .in0(N__7992),
            .in1(N__7961),
            .in2(_gnd_net_),
            .in3(N__9109),
            .lcout(un1_D_UU_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI867Q_6_LC_12_20_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI867Q_6_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_esr_RNI867Q_6_LC_12_20_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_esr_RNI867Q_6_LC_12_20_6  (
            .in0(N__7927),
            .in1(N__7898),
            .in2(_gnd_net_),
            .in3(N__9110),
            .lcout(un1_D_UU_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_13_10_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_13_10_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIGDFL_2_LC_13_10_7  (
            .in0(N__9398),
            .in1(N__9391),
            .in2(_gnd_net_),
            .in3(N__9051),
            .lcout(un1_D_UM_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_13_11_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_13_11_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIOLFL_6_LC_13_11_4  (
            .in0(N__9338),
            .in1(N__9328),
            .in2(_gnd_net_),
            .in3(N__9052),
            .lcout(un1_D_UM_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_13_19_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_13_19_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_13_19_1  (
            .in0(N__9268),
            .in1(N__9224),
            .in2(_gnd_net_),
            .in3(N__8816),
            .lcout(un1_D_UM_040_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_13_20_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_13_20_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_13_20_3  (
            .in0(N__8821),
            .in1(N__9182),
            .in2(_gnd_net_),
            .in3(N__9154),
            .lcout(un1_D_UU_040_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_14_9_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_14_9_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_esr_RNIC9FL_0_LC_14_9_2  (
            .in0(N__9026),
            .in1(N__8984),
            .in2(_gnd_net_),
            .in3(N__8971),
            .lcout(un1_D_UM_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_14_19_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_14_19_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_14_19_3  (
            .in0(N__8915),
            .in1(N__8890),
            .in2(_gnd_net_),
            .in3(N__8817),
            .lcout(un1_D_UM_040_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_14_20_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_14_20_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_14_20_4  (
            .in0(N__8822),
            .in1(N__8555),
            .in2(_gnd_net_),
            .in3(N__8527),
            .lcout(un1_D_UU_040_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep4_i_ess_LC_19_19_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep4_i_ess_LC_19_19_0 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep4_i_ess_LC_19_19_0 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep4_i_ess_LC_19_19_0  (
            .in0(N__12090),
            .in1(N__11126),
            .in2(N__10446),
            .in3(N__11507),
            .lcout(READ_CYCLE_ACTIVE_rep4_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12786),
            .ce(N__12643),
            .sr(N__12500));
    defparam D_UU_040_iobuf_RNO_4_LC_19_20_3.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_4_LC_19_20_3.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_4_LC_19_20_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_040_iobuf_RNO_4_LC_19_20_3 (
            .in0(N__9509),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_185_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep2_i_ess_LC_20_19_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep2_i_ess_LC_20_19_0 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep2_i_ess_LC_20_19_0 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep2_i_ess_LC_20_19_0  (
            .in0(N__12049),
            .in1(N__11513),
            .in2(N__10445),
            .in3(N__11162),
            .lcout(READ_CYCLE_ACTIVE_rep2_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12789),
            .ce(N__12645),
            .sr(N__12501));
    defparam D_UU_040_iobuf_RNO_2_LC_20_20_0.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_2_LC_20_20_0.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_2_LC_20_20_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UU_040_iobuf_RNO_2_LC_20_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9488),
            .lcout(N_183_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep0_i_ess_LC_22_17_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep0_i_ess_LC_22_17_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep0_i_ess_LC_22_17_5 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep0_i_ess_LC_22_17_5  (
            .in0(N__11053),
            .in1(N__11937),
            .in2(N__10350),
            .in3(N__11342),
            .lcout(READ_CYCLE_ACTIVE_rep0_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12809),
            .ce(N__12646),
            .sr(N__12502));
    defparam D_UU_040_iobuf_RNO_0_LC_22_18_7.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_0_LC_22_18_7.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_0_LC_22_18_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UU_040_iobuf_RNO_0_LC_22_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9467),
            .lcout(N_181_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep7_i_ess_LC_22_19_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep7_i_ess_LC_22_19_0 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep7_i_ess_LC_22_19_0 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep7_i_ess_LC_22_19_0  (
            .in0(N__11514),
            .in1(N__11938),
            .in2(N__10351),
            .in3(N__11054),
            .lcout(READ_CYCLE_ACTIVE_rep7_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12797),
            .ce(N__12649),
            .sr(N__12507));
    defparam D_UU_040_iobuf_RNO_7_LC_22_20_7.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_7_LC_22_20_7.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_7_LC_22_20_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_040_iobuf_RNO_7_LC_22_20_7 (
            .in0(N__9443),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_188_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_040_iobuf_RNO_4_LC_23_2_1.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_4_LC_23_2_1.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_4_LC_23_2_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_040_iobuf_RNO_4_LC_23_2_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9404),
            .lcout(N_209_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep28_i_ess_LC_23_3_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep28_i_ess_LC_23_3_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep28_i_ess_LC_23_3_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep28_i_ess_LC_23_3_4  (
            .in0(N__12092),
            .in1(N__11710),
            .in2(N__10820),
            .in3(N__10444),
            .lcout(READ_CYCLE_ACTIVE_rep28_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12842),
            .ce(N__12653),
            .sr(N__12505));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep26_i_ess_LC_23_4_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep26_i_ess_LC_23_4_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep26_i_ess_LC_23_4_5 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep26_i_ess_LC_23_4_5  (
            .in0(N__12091),
            .in1(N__10450),
            .in2(N__11064),
            .in3(N__11709),
            .lcout(READ_CYCLE_ACTIVE_rep26_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12840),
            .ce(N__12650),
            .sr(N__12503));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep18_i_ess_LC_23_6_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep18_i_ess_LC_23_6_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep18_i_ess_LC_23_6_1 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep18_i_ess_LC_23_6_1  (
            .in0(N__10449),
            .in1(N__12043),
            .in2(N__11708),
            .in3(N__10961),
            .lcout(READ_CYCLE_ACTIVE_rep18_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12835),
            .ce(N__12647),
            .sr(N__12498));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep17_i_ess_LC_23_6_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep17_i_ess_LC_23_6_2 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep17_i_ess_LC_23_6_2 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep17_i_ess_LC_23_6_2  (
            .in0(N__12042),
            .in1(N__10448),
            .in2(N__11065),
            .in3(N__11667),
            .lcout(READ_CYCLE_ACTIVE_rep17_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12835),
            .ce(N__12647),
            .sr(N__12498));
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_23_8_4.C_ON=1'b0;
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_23_8_4.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_23_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_CLK40_THRU_LUT4_0_LC_23_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12848),
            .lcout(GB_BUFFER_CLK40_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep21_i_ess_LC_23_10_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep21_i_ess_LC_23_10_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep21_i_ess_LC_23_10_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep21_i_ess_LC_23_10_4  (
            .in0(N__11971),
            .in1(N__11608),
            .in2(N__10447),
            .in3(N__11066),
            .lcout(READ_CYCLE_ACTIVE_rep21_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12825),
            .ce(N__12641),
            .sr(N__12495));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep5_i_ess_LC_23_19_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep5_i_ess_LC_23_19_0 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep5_i_ess_LC_23_19_0 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep5_i_ess_LC_23_19_0  (
            .in0(N__10238),
            .in1(N__12051),
            .in2(N__11131),
            .in3(N__11596),
            .lcout(READ_CYCLE_ACTIVE_rep5_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12803),
            .ce(N__12652),
            .sr(N__12509));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep6_i_ess_LC_23_19_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep6_i_ess_LC_23_19_2 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep6_i_ess_LC_23_19_2 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep6_i_ess_LC_23_19_2  (
            .in0(N__10239),
            .in1(N__12052),
            .in2(N__11132),
            .in3(N__11597),
            .lcout(READ_CYCLE_ACTIVE_rep6_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12803),
            .ce(N__12652),
            .sr(N__12509));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep15_i_ess_LC_23_19_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep15_i_ess_LC_23_19_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep15_i_ess_LC_23_19_4 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep15_i_ess_LC_23_19_4  (
            .in0(N__10237),
            .in1(N__12050),
            .in2(N__11130),
            .in3(N__11595),
            .lcout(READ_CYCLE_ACTIVE_rep15_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12803),
            .ce(N__12652),
            .sr(N__12509));
    defparam D_UU_040_iobuf_RNO_5_LC_23_20_3.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_5_LC_23_20_3.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_5_LC_23_20_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_040_iobuf_RNO_5_LC_23_20_3 (
            .in0(N__9551),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_186_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_040_iobuf_RNO_6_LC_23_20_4.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_6_LC_23_20_4.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_6_LC_23_20_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_040_iobuf_RNO_6_LC_23_20_4 (
            .in0(N__9530),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_187_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_040_iobuf_RNO_4_LC_23_20_6.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_4_LC_23_20_6.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_4_LC_23_20_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_040_iobuf_RNO_4_LC_23_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10028),
            .lcout(N_193_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_040_iobuf_RNO_5_LC_23_20_7.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_5_LC_23_20_7.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_5_LC_23_20_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UM_040_iobuf_RNO_5_LC_23_20_7 (
            .in0(N__12266),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_194_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_040_iobuf_RNO_0_LC_24_2_0.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_0_LC_24_2_0.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_0_LC_24_2_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LL_040_iobuf_RNO_0_LC_24_2_0 (
            .in0(N__9644),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_205_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_040_iobuf_RNO_1_LC_24_2_1.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_1_LC_24_2_1.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_1_LC_24_2_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_040_iobuf_RNO_1_LC_24_2_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9650),
            .lcout(N_206_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_040_iobuf_RNO_3_LC_24_2_6.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_3_LC_24_2_6.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_3_LC_24_2_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LL_040_iobuf_RNO_3_LC_24_2_6 (
            .in0(N__9638),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_208_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep25_i_ess_LC_24_3_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep25_i_ess_LC_24_3_2 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep25_i_ess_LC_24_3_2 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep25_i_ess_LC_24_3_2  (
            .in0(N__10442),
            .in1(N__12047),
            .in2(N__11739),
            .in3(N__10824),
            .lcout(READ_CYCLE_ACTIVE_rep25_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12844),
            .ce(N__12655),
            .sr(N__12508));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep24_i_ess_LC_24_3_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep24_i_ess_LC_24_3_5 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep24_i_ess_LC_24_3_5 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep24_i_ess_LC_24_3_5  (
            .in0(N__12046),
            .in1(N__11711),
            .in2(N__10953),
            .in3(N__10441),
            .lcout(READ_CYCLE_ACTIVE_rep24_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12844),
            .ce(N__12655),
            .sr(N__12508));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep27_i_ess_LC_24_3_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep27_i_ess_LC_24_3_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep27_i_ess_LC_24_3_7 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep27_i_ess_LC_24_3_7  (
            .in0(N__12048),
            .in1(N__11715),
            .in2(N__10954),
            .in3(N__10443),
            .lcout(READ_CYCLE_ACTIVE_rep27_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12844),
            .ce(N__12655),
            .sr(N__12508));
    defparam D_LL_040_iobuf_RNO_6_LC_24_4_0.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_6_LC_24_4_0.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_6_LC_24_4_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_040_iobuf_RNO_6_LC_24_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9824),
            .lcout(N_211_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_040_iobuf_RNO_2_LC_24_4_6.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_2_LC_24_4_6.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_2_LC_24_4_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LL_040_iobuf_RNO_2_LC_24_4_6 (
            .in0(N__9845),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_207_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep30_i_ess_LC_24_5_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep30_i_ess_LC_24_5_0 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep30_i_ess_LC_24_5_0 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep30_i_ess_LC_24_5_0  (
            .in0(N__10338),
            .in1(N__12044),
            .in2(N__11554),
            .in3(N__10839),
            .lcout(READ_CYCLE_ACTIVE_rep30_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12841),
            .ce(N__12651),
            .sr(N__12504));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep31_i_ess_LC_24_5_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep31_i_ess_LC_24_5_3 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep31_i_ess_LC_24_5_3 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep31_i_ess_LC_24_5_3  (
            .in0(N__12045),
            .in1(N__11457),
            .in2(N__10965),
            .in3(N__10339),
            .lcout(READ_CYCLE_ACTIVE_rep31_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12841),
            .ce(N__12651),
            .sr(N__12504));
    defparam D_LM_040_iobuf_RNO_1_LC_24_6_5.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_1_LC_24_6_5.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_1_LC_24_6_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_040_iobuf_RNO_1_LC_24_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9818),
            .lcout(N_198_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_040_iobuf_RNO_2_LC_24_6_6.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_2_LC_24_6_6.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_2_LC_24_6_6.LUT_INIT=16'b0011001100110011;
    LogicCell40 D_LM_040_iobuf_RNO_2_LC_24_6_6 (
            .in0(_gnd_net_),
            .in1(N__9797),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_199_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_040_iobuf_RNO_7_LC_24_6_7.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_7_LC_24_6_7.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_7_LC_24_6_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_040_iobuf_RNO_7_LC_24_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9779),
            .lcout(N_212_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_040_iobuf_RNO_0_LC_24_7_3.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_0_LC_24_7_3.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_0_LC_24_7_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_040_iobuf_RNO_0_LC_24_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9935),
            .lcout(N_197_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_040_iobuf_RNO_3_LC_24_7_7.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_3_LC_24_7_7.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_3_LC_24_7_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LM_040_iobuf_RNO_3_LC_24_7_7 (
            .in0(N__9731),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_200_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep19_i_ess_LC_24_8_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep19_i_ess_LC_24_8_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep19_i_ess_LC_24_8_1 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep19_i_ess_LC_24_8_1  (
            .in0(N__11973),
            .in1(N__11662),
            .in2(N__10966),
            .in3(N__10249),
            .lcout(READ_CYCLE_ACTIVE_rep19_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12833),
            .ce(N__12644),
            .sr(N__12497));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep16_i_ess_LC_24_8_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep16_i_ess_LC_24_8_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep16_i_ess_LC_24_8_4 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep16_i_ess_LC_24_8_4  (
            .in0(N__10248),
            .in1(N__11972),
            .in2(N__11706),
            .in3(N__10843),
            .lcout(READ_CYCLE_ACTIVE_rep16_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12833),
            .ce(N__12644),
            .sr(N__12497));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep20_i_ess_LC_24_8_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep20_i_ess_LC_24_8_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep20_i_ess_LC_24_8_6 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep20_i_ess_LC_24_8_6  (
            .in0(N__10250),
            .in1(N__11974),
            .in2(N__11707),
            .in3(N__10847),
            .lcout(READ_CYCLE_ACTIVE_rep20_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12833),
            .ce(N__12644),
            .sr(N__12497));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep8_i_ess_LC_24_8_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep8_i_ess_LC_24_8_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep8_i_ess_LC_24_8_7 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep8_i_ess_LC_24_8_7  (
            .in0(N__11975),
            .in1(N__11666),
            .in2(N__10967),
            .in3(N__10251),
            .lcout(READ_CYCLE_ACTIVE_rep8_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12833),
            .ce(N__12644),
            .sr(N__12497));
    defparam D_LM_040_iobuf_RNO_4_LC_24_9_2.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_4_LC_24_9_2.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_4_LC_24_9_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LM_040_iobuf_RNO_4_LC_24_9_2 (
            .in0(N__9929),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_201_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_040_iobuf_RNO_0_LC_24_9_4.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_0_LC_24_9_4.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_0_LC_24_9_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UM_040_iobuf_RNO_0_LC_24_9_4 (
            .in0(N__9911),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_189_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_040_iobuf_RNO_5_LC_24_10_0.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_5_LC_24_10_0.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_5_LC_24_10_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_LM_040_iobuf_RNO_5_LC_24_10_0 (
            .in0(N__9896),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_202_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LL_040_iobuf_RNO_5_LC_24_10_3.C_ON=1'b0;
    defparam D_LL_040_iobuf_RNO_5_LC_24_10_3.SEQ_MODE=4'b0000;
    defparam D_LL_040_iobuf_RNO_5_LC_24_10_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LL_040_iobuf_RNO_5_LC_24_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10022),
            .lcout(N_210_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_040_iobuf_RNO_2_LC_24_10_6.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_2_LC_24_10_6.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_2_LC_24_10_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_040_iobuf_RNO_2_LC_24_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9851),
            .lcout(N_191_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep10_i_ess_LC_24_11_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep10_i_ess_LC_24_11_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep10_i_ess_LC_24_11_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep10_i_ess_LC_24_11_4  (
            .in0(N__11606),
            .in1(N__11903),
            .in2(N__10336),
            .in3(N__10851),
            .lcout(READ_CYCLE_ACTIVE_rep10_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12826),
            .ce(N__12640),
            .sr(N__12496));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep29_i_ess_LC_24_11_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep29_i_ess_LC_24_11_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep29_i_ess_LC_24_11_6 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep29_i_ess_LC_24_11_6  (
            .in0(N__11607),
            .in1(N__11904),
            .in2(N__10337),
            .in3(N__10852),
            .lcout(READ_CYCLE_ACTIVE_rep29_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12826),
            .ce(N__12640),
            .sr(N__12496));
    defparam D_UM_040_iobuf_RNO_6_LC_24_12_2.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_6_LC_24_12_2.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_6_LC_24_12_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UM_040_iobuf_RNO_6_LC_24_12_2 (
            .in0(N__10004),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_195_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep22_i_ess_LC_24_13_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep22_i_ess_LC_24_13_0 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep22_i_ess_LC_24_13_0 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep22_i_ess_LC_24_13_0  (
            .in0(N__10854),
            .in1(N__11901),
            .in2(N__10241),
            .in3(N__11489),
            .lcout(READ_CYCLE_ACTIVE_rep22_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12824),
            .ce(N__12642),
            .sr(N__12499));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep23_i_ess_LC_24_13_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep23_i_ess_LC_24_13_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep23_i_ess_LC_24_13_1 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep23_i_ess_LC_24_13_1  (
            .in0(N__11902),
            .in1(N__10170),
            .in2(N__11586),
            .in3(N__10855),
            .lcout(READ_CYCLE_ACTIVE_rep23_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12824),
            .ce(N__12642),
            .sr(N__12499));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep14_i_ess_LC_24_13_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep14_i_ess_LC_24_13_6 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep14_i_ess_LC_24_13_6 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep14_i_ess_LC_24_13_6  (
            .in0(N__10853),
            .in1(N__11900),
            .in2(N__10240),
            .in3(N__11488),
            .lcout(READ_CYCLE_ACTIVE_rep14_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12824),
            .ce(N__12642),
            .sr(N__12499));
    defparam D_LM_040_iobuf_RNO_6_LC_24_14_6.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_6_LC_24_14_6.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_6_LC_24_14_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_040_iobuf_RNO_6_LC_24_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9998),
            .lcout(N_203_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_LM_040_iobuf_RNO_7_LC_24_15_3.C_ON=1'b0;
    defparam D_LM_040_iobuf_RNO_7_LC_24_15_3.SEQ_MODE=4'b0000;
    defparam D_LM_040_iobuf_RNO_7_LC_24_15_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_LM_040_iobuf_RNO_7_LC_24_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9980),
            .lcout(N_204_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep9_i_ess_LC_24_16_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep9_i_ess_LC_24_16_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep9_i_ess_LC_24_16_1 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep9_i_ess_LC_24_16_1  (
            .in0(N__11925),
            .in1(N__11538),
            .in2(N__10232),
            .in3(N__10968),
            .lcout(READ_CYCLE_ACTIVE_rep9_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12818),
            .ce(N__12648),
            .sr(N__12506));
    defparam D_UM_040_iobuf_RNO_1_LC_24_17_1.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_1_LC_24_17_1.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_1_LC_24_17_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UM_040_iobuf_RNO_1_LC_24_17_1 (
            .in0(N__9956),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_190_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep11_i_ess_LC_24_18_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep11_i_ess_LC_24_18_1 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep11_i_ess_LC_24_18_1 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep11_i_ess_LC_24_18_1  (
            .in0(N__11926),
            .in1(N__11535),
            .in2(N__10233),
            .in3(N__10969),
            .lcout(READ_CYCLE_ACTIVE_rep11_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12814),
            .ce(N__12654),
            .sr(N__12510));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep1_i_ess_LC_24_18_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep1_i_ess_LC_24_18_2 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep1_i_ess_LC_24_18_2 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep1_i_ess_LC_24_18_2  (
            .in0(N__11536),
            .in1(N__11927),
            .in2(N__11067),
            .in3(N__10148),
            .lcout(READ_CYCLE_ACTIVE_rep1_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12814),
            .ce(N__12654),
            .sr(N__12510));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep3_i_ess_LC_24_18_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep3_i_ess_LC_24_18_7 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep3_i_ess_LC_24_18_7 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep3_i_ess_LC_24_18_7  (
            .in0(N__11928),
            .in1(N__11537),
            .in2(N__10234),
            .in3(N__10973),
            .lcout(READ_CYCLE_ACTIVE_rep3_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12814),
            .ce(N__12654),
            .sr(N__12510));
    defparam D_UM_040_iobuf_RNO_3_LC_24_19_1.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_3_LC_24_19_1.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_3_LC_24_19_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UM_040_iobuf_RNO_3_LC_24_19_1 (
            .in0(N__12350),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_192_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_040_iobuf_RNO_3_LC_24_19_4.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_3_LC_24_19_4.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_3_LC_24_19_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_040_iobuf_RNO_3_LC_24_19_4 (
            .in0(N__12329),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_184_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UM_040_iobuf_RNO_7_LC_24_19_5.C_ON=1'b0;
    defparam D_UM_040_iobuf_RNO_7_LC_24_19_5.SEQ_MODE=4'b0000;
    defparam D_UM_040_iobuf_RNO_7_LC_24_19_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 D_UM_040_iobuf_RNO_7_LC_24_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12305),
            .lcout(N_196_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam D_UU_040_iobuf_RNO_1_LC_24_19_6.C_ON=1'b0;
    defparam D_UU_040_iobuf_RNO_1_LC_24_19_6.SEQ_MODE=4'b0000;
    defparam D_UU_040_iobuf_RNO_1_LC_24_19_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 D_UU_040_iobuf_RNO_1_LC_24_19_6 (
            .in0(N__12284),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_182_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep13_i_ess_LC_24_20_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep13_i_ess_LC_24_20_0 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep13_i_ess_LC_24_20_0 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep13_i_ess_LC_24_20_0  (
            .in0(N__11994),
            .in1(N__11594),
            .in2(N__11069),
            .in3(N__10236),
            .lcout(READ_CYCLE_ACTIVE_rep13_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12804),
            .ce(N__12656),
            .sr(N__12511));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep12_i_ess_LC_24_20_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep12_i_ess_LC_24_20_4 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep12_i_ess_LC_24_20_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_rep12_i_ess_LC_24_20_4  (
            .in0(N__11993),
            .in1(N__11593),
            .in2(N__11068),
            .in3(N__10235),
            .lcout(READ_CYCLE_ACTIVE_rep12_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12804),
            .ce(N__12656),
            .sr(N__12511));
endmodule // U111_TOP
